// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 15:05:47 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FKTTsukS/C69SFhV4NRC4OvoXtM6nDjk/bpKYtELB20fo5/ua01sPQ5iceCA1bBp
zswKgyLxEqV0drkF3G6EF4m43QHMO6+yekDl3VmeEyYxj0QNsWLiRR20VoFrXChU
YKFzEu4ZxLhaDeadMjF2uhVyxo/dPrSSJznEpNb6KZ8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14080)
KFmZWB4SEfY/iPbcKfTbYtWxic0nCgVgrnpENSZh7PWR3GZadd3X13kNs6cHLZtj
V2BWRkXhGkMyIJBbs0QyIzhhSzcj86d+9QR5lRL4Xb582NC6wh4WoQVAn0zYy2qH
vJJC2Klw2yXw5WdNQHYenlAIyBBkfdbMomZeANnECjCtS9lWLZKMWynrVZzBqUy5
yCPePP8XiJteSp14OVLORX66Zw9ljNU98Miw0FyPEQ3ZX3V3WjfooWvBSM3AA6/2
I1oeKMkvMGYfzjRMGx3RMXeT8Jkd9na682LbRaEc7VN5cJE/1vnDeUetp76+N1JO
yD3stepy4ZhT9ZAuTJe76g8F7RBe3o/nGudeRCjYi/PualSWoTtWyz/JwrUa1oaY
GJNnvTVVXyjMq/BnSc8Lx/7j7Zelr/Fz/puC2abJRnRlm0zQpVrmOnSBYhulqlRk
9UF/AxnvFhMV0cbimiuoml97CLDnibFlwBirRbaOLGjBkur8UnK2FD/PNjpQrSmZ
KNkdVDMGofwzj60O9krZVXSHTnVoge7K0MJzwPIZX92ieMuNTLBPX/aQv9g6t0yH
+ridjfnT1mSQ5DI8vgLbzEaSGBhsD7HgYvnEctfWgosegQ6kDKsfwrsSNENP8fZB
hdsnkCQhnwjbiiZwuFxM6VpTTwsEeQ2kUQ2DyEqaglvv7oF/bw+VXwFwjlseUIWN
y95tWMLEPQUFI4oy4YrFD+RlbCJop9PPK/MDnTdBC/QjmJMfOXhs3gHkzcfJXGQk
pJTLfkzlkAL5zw/d5qjfBuuWrN6PgCgqJu1rij4J3maePuhB/vPbBwfPxes/55Be
4fL32OM+DbFD4yYF5RqOped2tgT7Hw8vYdPIc/1BRKeQlQGT7bTE76vvDfckXiQk
aDvfY7sbYuht49BzCBQPaXLebHIjdtfc5ehtToQSAEjpA59qKKS84qIyeBBuo0Qt
IFJaLhVfMnpz77kmCGmb/tsi68EoN5TJ7zmxq/JUyorSdKXbM0NTyD5WDPeTVhNZ
B/Sdy2AAOzKz1uwTfptKvJWTNTAbqrZrfbXnmLUIfELGtfzh6zTsYatx7pRwmgD3
cIU/0gS96ftvAVPO6RaXXWss4VwKf8RwdJTf5jq7Sjiu2zHRE6EEVXjfMoOmLDfD
iKzhC/heFmJk07XDLKrQzo17F6a9qscVQ4a+60fWjCOGMaRGncuvPNGOfsHNMdDp
9jRcItnfgDRfXNjXC3PJLSSX+ooSnwCxGojbfaqi+kBjHKFkerNk4h0H7LsHhmr9
4QY5Ga06/srimHMh/y5CS9KJLR3ryFGy0hLmKK0q/V0eC1uB37OkOhAx+hz5t51i
xAoBZ+858R4Rjak3P0p05DLlET45QZcS/JgbY++q31N33rWv0fFZPc/OR7fUeBlf
teolihHcuhR42nNkZ6k8mBvp5AvzDNN4d0xXwv6H2ThOH/nN/Lx3ZXd2e+ONcnAR
g5vB7BxHg729syyzK6QZqarYs9ozvJH7ZkoAaJOku8FIPqD/Htn+lAa296wg+C+x
+6XG1qZCrFIWTBfkkdexhvkBMpdQqs6LAQqKKQ7WpVO0oBd0KlcqhN3ilMlx59XX
BnS35PyvkSTEjiPFRq5ONXFe/rLBgz/2WxTMo6ypDSx6QexuLmIKFOQaS6E6bP75
v9h/jUME1pCAWh/jRtNKjNatz3j4msLxHcsnmsIVKR9jyIG0ItrZcHJSuiLVuqf8
9qa0v8+1qFIBuHbq/HfETkm7NpXKNv/WycMIO9WMgICgOdqP7m8Ln4GnSzwTzE+N
ixm9FQjoIWQD9rO0eGaNSLrYWcIB1rVJ9dyesWjXwnNh17cwQOgkmqI4d33QClGx
kTR0fH09dwZb4DU7lGlZB+CTBEQqM1XVm4icaFzaiZxSr7tsTDezqnBIdPmahFuP
a8c7f8wTZVmrJyFMnqusiCC+LnMW4W/nIZDssfQAUXB5tv7OT8nwDe4rQjCo2kzB
dBjXjz+kz0zGPoKMy/xr30JF5q26gz8uP91UAm35QcnlcOLJqczsxebI5mpeZv74
43wLDjnh+0tER37RLMZRJMltRzPaSxdrpv+R6M0O84qdE3yXS4Er1hGeLSSndnOX
DfGzewlcoSryMBomP5tJjgXMuG8KOQ3AROTeF0QND8Nr6aCY1F54nolCUYlj6kU3
BuFamz9DMXto8YKh9sJ2dTMnJ9jqsh6zw2kumWMN0WznP2jrl/Ul5P0TVQxpvaJi
8GLS5Eq5BW3Zw+Sye6+2DS3r6OfypbpekfwDYtozjTcsAC7Is7EM9v2MVxEtXPqP
BckJm38JzhCj8x94VK2WLEN4q2RdI7S2sleLp1/gYpmWsX0uvbNf25FNFwTlsJR+
F3nc94ubcM7IVlp9wbHiE5+3buIQy0kJNWzK0dWfqD/JB6Z62aeHzrh0Y2/b4dp9
HXV7pRddQiN4QMxm3RbHjxjG7qeRrHBelPA29t3V8E3+FQWMxJFUirjZiKLplvPt
itxBDdd6B+L7B4hvWAECWpjAOsLrw9wXl+fTTjNjc5EMuQmtQs8To7bCHOUOYRwy
iOaUg+dV738sIU+0Xzc6I4j6bHm4jJTo2Dr0YpGSK7yxUEC5zM9oKIDQb872gosV
VwqlKKAbDzHa0Rfeurq+Gl1Jb0Ie+FlGZX0a/vZf9LvJ7hgc6J70JFoOdsY3dLeM
QV6FF3Qf0yr0fixl5dDclixjuyzwXpxmOjZERcG6f/47X2jkXK3f/TOfTSuPESQK
TBMyL8QjqMunlb/UVmg/xCmEdrxQHsrqT309C5f/Nu3Xvg6DSCXZkgKUTnxxi6K8
jWT8kcX1R/s90GV8xOqU8sVAmcvgMNhqLrZCpmJlEAjMKdsvtWRrwDqs1+kUeyKP
w9bAOdyJ9oWMyK7ntpylfvYtHH4YhoLjFNwgZECDP4i7QgclSar6W6uemttOz1Su
zPhK44nPNEL32KB8WuLLFEfes4Jzk9PgrbQfJio3VlMHD00HGvm9l0TflKZxsKjC
t/v2hb6j6fYBfNXXimk+WnsGmGgdnrL9AT4cOcn0NR2C0WWlHLkgDNcbDWDfZL34
gnV96xzHdx6OtCMbNmMt0Vg2dYnZp2SIB5VmP896J/tgMofae9ONT9SMnqNf6UVT
dZ6K04XOiIATeO1CKWTKnrBjxMU3t3aYz+dKLOVfly4aUEpCDb2DE+V+QWugsfeP
qShX8PEcBWCbr53Cgv0ICU4TqS6SQHSaJV3hCrLhWt9DpiDVV+ZqDDPpWieajH1B
Ux29RjTawbAp/imLR8SJ1yGMVzXbrzJw1nqlEPn66Dbqw5vNrzGqoxnZoFBoVDxu
7CP4y3/WRCm05wqoAbHQ3Tjpf5TNPu5VXXn37jqgjh3SBuJtU9Ea9yC7ypxOVJ0c
1COUPQ4TfhNOeDlZ+AfW1047nbsUsq+07iq5IITqzssyIAUJwzdJ7ZaGJx3ehUjM
vfpHdcrZG0k8UfvXfEGfx3Qs7x2tZXWy/Q17Oag4ITq0VfbU4uTJVskr4d+WppHc
1Yn8sdqSoP2g+fBm62rgJVXVrmCtU3Nca/fz7Dhc2VFwX9JyKhWI1wUytw7gBOsO
aOmnyr5pbxbuIPTWNbNr8ZJJP/6AT2PJ2wIue/CpLtDQMC7zZqYz+XPJWsXzuxXZ
0xJQTD/LbzjLbpPVAKQzkKa2B7fseeltBTbvnyC9t8ri6IpU/jFi1SoRg5bHb9Tq
Y3+IH/jIEQJN16Ce3lBnknUwUni94RuI9y6VSQrjSc0YHdi1Gi35KANm7tz1GaQr
xxzyQ0TWF+KTwXdjpZLVTojzk/DzuCw7FlzdN0qNXon5XDWI8aWVtbKsC3Woax2S
GrwcygR8w9lQ6Nrwsl4j4ExYiMoXxtSQjPBAVHrUIhipN+WBsOlaBu9SjQ2b9/Zn
W/gBcGMD9a0McEWa15q1K8/sMNP1s8qdFhdy7COADf4D6JNGjtPoIk1P15sDXWvx
riMvAnfsFVDKZCXl0AMjfndhi0YfsJrd7FOxjg1rFO5nZNrVT6k2Wz09Tlgv8nKI
ZI/9BFZIAtqsd4RMs4vVNhfFf2uuYQPUTmHVHQs4OGai6ZAjqikXZZMBqsjjI45M
2ScZm4W0KkM+ukiHZEIOT4Fe6BHajNQujf0jE3bo42lFrKiLemRNElIBsrZ4MKMf
JOJnESMq9/65f7Nv4QZ843Geqwp8XFMj0OpqlxmRmtY+w4yX64iQ9KzIZnFQN1CF
l42IuBAt+knwaN4PvxfRXsANiowaLd6HlIMvjplS191s6UtOEm5yqLOngxGWIpWg
RLJoG81N1mVqi7UL/d+ptpyiWaMVKpi4VeyayKnwQQQI5JEX1xV4spcSqauPclYY
2uRSopewj1L/lnCBkJPi8zradlybHjwLlhG6dAh+mcyE8/ErQJEN0Uk6y8sDKYA4
Vj0MuwzMmuxphVUEDgIrFxA9P+CtTASgCgGXyUao1JE12WwnnCWAOto9km5Qdh3X
CQNPhL3AWMFnSl7NzE6sgvR0iMgGTEi/A6XErgx1WV5nIgH2XDz94vIsliG4qOpK
bnQ82ysh1SDaX1WLfBk1ld1d9PMlSi1gc2o+o2wdQv0qhZEjDRqAPI+b/KUJh6e6
ygMsJi3W4NFR83qoUa3dkFKuQKjtrc+G0aMrTMysIu9y0XTr6f2VjV671JPrlkUb
hYqfU8OTgADUy8iZ1aC/vpCKWroK/wNoWKPx7FMqqw15ywYTzHh1U9vYZv7So4sI
f1SM8BLLIMevygR/IJhtSIJdYqHiPHTqO7aEVu61dvV7V0sOIaz76bDZvKq93msf
njgAocVTzIQd/oFbZsLBCtnCxVnzm32TpF8x4756nrRGs2FSWsclxm1jzS/WokJJ
18+PrgprT+JsGd0jD9tjeBzjZyFiDdBR+Qp9z2z/1BzuhA6SH9tWLey6Mdgwl91b
DFZg/tIpACmOxhuKkg6B2skcJSnvDrISeZJMOTx1VnAI8omJc/Wqex+ob5ena4J+
J8KUb4+WHYEXArK5cDY76Dm9TB7upRIRevlahm9mkuxIoUtZcQ9NZkUR8vccweV8
u87pSxQmR3w4Vf4lcf0hjEiJXOk5vwJXULYb/eoEdcB7SGjfsinuJdBAqeZM638w
cai1sXipJkAGGLKWQtHjZdYtTP4iGH2DIt9kyji3RKRapNdKvk8MWaHwtNXkcYgd
UOPI7PX2kvo2DKHjfQ8dBWcqyZ+jOO7Nt5WyOhuagNZiEasArHUcezzhLyRvNfLk
n1px2PMl1ON7ENjheW2Buu65y3mqJV8mmHLUqWXKmhiE62dV6RCkgrfZ6v3IWhBC
xGDdEfspFz41JNk5c/l5qK/9NX9Yzsj2AVa231R2U55bRHDgZgX+zDO6ry4MSZyr
4w5BBA4Np7ferpNg8SucuFnAbb7LSUjAOQ389RuXWBha9t72AqU4ba/+cFBqEzdA
vDmOp9q2UGXs0KHB7mITcay8j0vIQGN4+p82Vf6smtpPRa2pwet+esSk1Q0yBTs7
Kp59v6oKokZaHef3zkAzNPkbrZVkBisgiKM7VtgcAu4l+mzCNc+7rWUQqB3sa2EW
wRhkDBumbpVlntq6ybKN3b5xgLZF1cQUBzG8EuXiD++E8A/rq8oMOpC5nw8ce+ML
oFFld0P7skHjb9x0ItfC37wL+SC+SIHEJr0XwSOXw4yAO6eW76QR9ipUxPhsJtd6
f8FvVyDW6H1cVgIDf0u/r/u6+DxFy3jTJjXGekoHC+ptd4rhF55Y8bh87mYUFgYS
EJUPKPYJcif7ZAmRONLt7tJSaFoba6BtR6A6nR98mPXqqqhhnOzeqm8d1QGxZdbE
Xtob+hVl+Swvx0j9ZirlwtmBxPE7d50vXZto2uQ2W3UD8n8e2NNpzFpTcf7cUGHM
xu2rExSxxF4pyKLbR1R8v/l0xD3WRtN+S0W0yzipiGxd889kFcP/+Mhn7GoBgo9v
EbrP2HwJQ6U5FH5nbb1Hd9GwYFywhWThxxe0RxeVzwyT5LPHmh+FswN5dLqU+w4f
nT2UFt4ltH4ocL29E+i4DLjqYio0XAM2+m4c1gim5TsCabfto0gdmfOn5SZTLyRy
ijf6MfxJoMr7LRAY1tvlRjbNbk71yHLAPMjbun5JC9EaJd2lFluNDcH98tFB2FYK
7hOAlnHbojNjhbf7PSEi05V67n8jUMxk3ABmlgspQnIsm+GNwd2l0VZlyQ4V1dZW
+7s2aIFIAuqyYd3aul/Lgi11fwg2tPNzZ9h2YrHQIHJN1xpxNKjjHVoBj73OOAM1
tulQwGhdrLSpvjtAIryFQW4ih6JNNedEhldQjS8GscHWDj0g2wQI0gydw48xjk7z
ZgUsjselj3gNeTxQFu810BjokXnnK4gRe9R0cbNpNfyVBHpYNlkebE3JZrueNqTX
npp4cEdk2WqLre/eXn5l28VET7Coz4Wn57dBXkUKPrQ9lQVnFwBJv0NBinMFUvrB
AbQFwHEAfsHduJa4ZY2Bwc9hV8Dp71CLjuxh85kP+H2VqNRfCMOwrhapHGX71WOE
+RcwSf+bOxt1C/jpZICWo5SbIcSrbx4itw0Dn77ly6+oMwPuD/6wYokD/7Y+M+je
BKaYj29dC2THEiNyNYHHd+p5s6vssVw+dCEnuJ0kEt67NekAA8veVldBTWdfOqXr
X8YfX9a6FghdmnWE4Az9fcymT753EjsySRLxaVWkjap2v6uTZd08k9HCe1YcXAiU
LGgH9Xin4HM+EtXRF4ihl/4d+1+JkPMnclaJSF3jUX40ldK525uMe919THqSyxWn
paCUTjbTzqR83KN7K2FlpXNFL1jhkhzBzPRPHNVpIGsWMUyCqoJnOEWZp+FFBkhT
Y218A3/NPNYlLkhgmldOwStKlBeBcG6aXS/xVHojP35e0H2XEOG3uifnrYwzzRhv
iFt9T9RYFW5PnvJ5U91ENl3LOfkOSj2JeyxcAgFfMgvw87y/J7F6Gwy4xpr3V9yp
Ex15v6RYODM3kQKkLfEMQM8iFF5ceSWxmvMp/Meg/bTTpNcnP9EzosM+1aIuSKpt
VGw3w3xQ/P++Q5s2oOyqoBEsmHVUW9Gh5CAGOnvzR4b7Welx4rW1Id19UvpIrmj4
Jv68QFcCt4VINJ1sv+JBVzAB7sPpzMwba+XH7zwoDEwWsMFVdwsR9PMy/i3mAtNM
9rz3AUrJ33ngo9HpS+S45GCd/mqqCbWYHBJ0PQxu1Omfo+/kmFxyTWy8M6oGgv8+
zqBuUV9dPUgJ8xSbbckpKq1Zot+/eXyErihuAQ4oOn9nHbC9yPCmQIJyPLJvSe9x
8nQiNrtDczNeajKTqR9PyvnL/ORm+s0RRfuGpTY1Wf3uNQqvmseXSh8IVtpP+dbJ
AIrF4mUs+pQiaT7V+qP5isePWizcZ4kA60SLlVBOKyUermFxXzVwgmcRdSLpWAur
N1UNfpGg55piI3m52y+p54SbKQ0xZtabSFDjBekEa6WqbC81zPWNrUQoCOMpihu2
R3menDcPQuI9PkQ2RAZRDB/Pq8RcF8ZmkSzlY9YBJYjhjRC3QY1uRuvF9INzZtO3
AlYUR99aoKb1W/9ATxSCpFAn/P9fHrn4WVrAlgQUhVb79WaFViA80J/Vkbs6pyC5
uac9kR6dkFn/txPVHB/4TAhsGYbYo7Xh6RdExjfuFI7Y+IM8Vt338Oh91rcTKVBY
amefwnuQER4BobhWqOofJWOrmsHt0Yi26HCWiOZVrNj4gDazY5Gkhjdr7VyrvxJ/
x+FpVZu/H/uYeVKovHYblxXlzrlcmtIwNPUGNLFV81j9BJM+VecpURShAbh5aBeh
zVyozz4xFRys/5FAsJXnSWhijFwWQaAc676jAFKg5wG4x5nGz3jOgX+LAGQ3Jd2Q
i/QaIMdpxd8csqfgUMQfmJ0pyp2O2wnOD6hAJhdEQof4XoRjoW/TARslQkSEWHbO
uTBf+n5EQvqJPcdslOevq70tIPsquJOs1IHCw+tODbpysgl0FLf9bxvnIXdoccIh
QH0pPbeVGDa/6M/EIvvJJHaKNmjYUKjhfJez3ffFFjIpbbhQomPHKPtpV+Iqeg7x
jEyD3/FLQYqAcSlnkv2KShVePHFPtAoC/zJUpUO25HFJTpn38xBxNff4FYsBV6kc
EpFoGLYYRiXnT8CGC/WX7VnTgm40wUzVNFybhw6MGELLrwIt8oaXzfnSKdKzB3Lz
Pou4l9/H9Tjoc+q5UNbxu8hN7LaFHCwSB+vC8DECxaiVoucjvuwObSkA86QG6F01
kdhGlOgqrgQTkxxWaHS5mCVBX9fjQlTy2G8m+qEIZPvyIQ8uBAEZvQ+5OScJaLXR
RQ8l2UBjBy4zzXK27A+Qu2TgT2WZvCH7/WOvKzua43+baFaKI7e6PzdAbPlz7SPp
rxDpfUyPsq0cPX1AsYcistNl4iVw5Pb48tE+nDps37QZvVh3PEHd8S838Nw8O9G9
6ebPEuwt55+MktWzPqxNWkPgCTN+WKUjSbRU43g2xREVF/z4pYGwUPuAH64oLbIg
3EdKzNUhViLieShzt8/LIGsl9bmqU41Whu5FgdaX/5GrfXR7sdt3KWeOVTajoMX8
GksSik3vZI709vytH9VEr+rOP+JYIlDj10EuQ9vbtX7fgdVzl49+zpe41pCFhz6P
TnGqn7TGd3x9tcS2dJCQIgfOlOB2Hhfvz2Mcu16ikvoRVITgBErHDhz2yeKXAtyk
QdDuXOV8QkPYmKjWQ6yTAuP0kAPTxRMOzDfB4AihMCulT7D7y2qlIrxHzKZ14QJD
ucLgcaKyclI0Yb+lMV6yfrFZZgAARL5QhgdOB3g6Z3PsI/L2dXqnlBOpBVTBdmSJ
ymHCkwyRN+qHSjDl9V2ToUxTdc7XZzthZZ63vnQjfBoLhmUu/YNiB2V6dUW4YawO
D4op+kk7PdqdcZqk561T47zT96fzMPLl9hDYgJT0TDsM72d62YJUQvSySukAbr3W
vFoyflfLliYUK8tnqkJ2yhmUc92OZKfsDPiKPDefMP6JWzjHLTv/8V4YLyS7sU6j
4FE6oQ3mnt+OFHHSLgOaIeOBA5B2GJikkPZ8rFJSEK5IuxmfgEY6sDXYvM+tH9cR
c616dMU9oo/DZ4t28DvG5Rkn+XSsIVS4HmlNqNKRY0wwAxDxEN2Y48IrUi8bgnE5
xL3AQMIz9pgYIQO/AYJZ4487uZJ4ijn3NmDClOfhpycKGvK3L4waaxIrAZPNbISx
tUMvGqaeRdnH4Xs3/OzlINQarzBrH+AlCS9C2FUHW0x0MPSquw5qou3ZqNc2vWbO
YTPDxCvnq6s30pKQRI326VkAvxv2ajqApWEBv23lCfABI1z4brFzrOvifeESKPI6
pp2XFGQW8h8ORScfBuKppuSebEMvnrSRjMIxyyfZCluLfzhRCohzv3TzbGqAfofk
AYo8kChrxSigEJp6oE6i23QE3EzcrfVIGoaBchxj8Oa0a1dwB9zLqu60qCy/vmEq
9ehZ7vMoQD9mDMRCv6YtLIItexH/Txqly/fdVPztS7QrPl2kop4XNvRz4nC+ODq4
vyIqTqBd23Q4gkGovkWhQex6R6DkCi+VXzzMKfy1PrGEw8Ds9yalOkJfgSiPmBTK
qHJF4ZsiqLYd8ERHKryhaMT4Yv1TqdJ8hnEXAF9noYhTmW7yLZlW0lIAo9T6kviU
bMxPsQdGtv1jhmDrcbT4J9ZkDF+aj5kqJ+oInQUQ9bWFDKsQu2KxS1dXz0BwwM7O
L8iMLVgTYV3p57xU0WgFAuGpPdASehgGrkcc0FEcH7VidvnYv9XfGRUpr8o981G9
g8RG6/zLVoOjoYVXA1enj71ZCOJ0/FYrNJ+o9mIQ0s/QZoY8T9MXMXyi0nGjPBTC
03kNx99vOw9z4thr1Rtbj/EUSl0z7KaaRxw9Wd7FzBduCC4nx3M52+Pjs62dAsI4
ulNvkJ9Y7lQdBEYaSsMZFn7niJ4e6ZPvfVzyteAmIPVXZKrn5wXD/TPQA+kagFBS
VGZFmwRMO/ktokT853NwS8r8H6xlhft76PlASRKstktYtfsXI7hY+Xei2yAeZfYU
fnkVanxRvvbKp6t8mfXcA+MxkLV8AS5ufk/c7WSYJ0rN/agyPpuXCcExhHjO4zbL
ZkYAnRjNU8FPiFh2VI7oL62tmDkseRZnJR3k6+6rIea5FUeKfyDAqw28OfG9UpiV
dKU1JYC7NzkuTp7kUc/i07NKeXSitcbh7xqOBc3amh2OEh0+WYLDnU0uR1QfEU0N
L+SnSX2OiXKSbqS05mn5e/m5lThQmt8cCc9uIdvhiTwOUZHFirlhs5k++tfrMgue
GY1XqqjfQZ0BgnF+m8yAdYtAO9I1eXLZE3q60u6Jw+GvZ67TQUzHi80tgrF3sAy3
VadbBuORAcTCYluwpPRaL8G9jBBbzuwMC4aya7d1lVEUR1ANQbmimeBnqvGTp8RV
G8hPntDwF5XwAuNbovOF9ueI7J4cGbSuYlBY5onWpGYMizyoq1fPLljMUIOsCjfL
4WhvSmqNb30speXvAWm1r+soi0uTKQwgDXt27xVhjIob5PdwgFJsqOEvbBnUODbx
9Xdkh+0xsV/4ehB92L6bY1BsL34MHSR+w/G8qc9hhIPB2ImFfHdBFCIEN3dPVHCv
8Cx3diaDrTxvBy5GkSXrPMritOmtiPgiAXJwTX2ww42WhgJ7IRAXEJQKHhc9ykSd
kg9gd4quss4wbRane6sY0/pGWoRs+dli+CxcD1F75wSV0AjQlEqtVl3tfYX7OJJI
/MSh3BU/rykcR+7rN3igwyMjKiWRR16iMwsWg3ocADY1qxsCf2mCFpW9k0WiGbXv
0BP/p/yCWVWf+QF9/onR2GW+OH+JYC//ZdPFXkZFzeRZO6Uv8/hv8uIzTisiTn5e
h7ZE7YAwdzSMLENz0qf7AlPNku7NZcyfbE/PnON/K0XaX0A2aVWIEAH1Caj7ZJyB
Zs3/QVicqBpQE5UkEVe0DskBN7I538kXKnql7Q7ZZl963iJOk1apAf+tfFkcp1qy
u4FsiHuAWyxy3iuzn9uu7cUrUF8VjiZmMqSwviPrPXnIOgsXruf075/t0Q4xaBcW
t2ezSuC9Ze1FpDUcSMx0Z/K7BLu7lZXSak4TgoRW4MCeFz7YPucqCxqCXq6/L7Q4
hfsDoIVhSLOOpRYZaIRP25vjrjfxZT2lSaI9J6/FBs/hKzPYLKlnAHPTHwhOw34P
zngI6AaGJYk7Kg8jSakf2SpeFwTfY1I4HoQJGl5OYBokcmo0eUfJTCJvGAfNNwwP
I8FZvX8RuVUu2jVd0J8gvxLoMhLpt4TQhR5w34YgYBpk08rf8Ewv95vikFUji9DS
aZ3gbnbj0GmQAMxvBJdQ6C+eyu3Tm0bnPr+Lr+pLRAlRZ4yn/njZk/5CQm1RbaOI
G2UF05GTI/c0TQeG/TyvYKHpX/iasOhitb2BeLdT9jixAsu0F5T1B2ivDt67VI6h
sVzY/9QDq2SsGP+fGDsI+1KemzelU8NU/4bXgf7O4wLK4cR5e+319qMAV918Vqnf
uUeMzx4jwAcL99nkP9iK+z9s/UTzL27GB1yvhIaptdhqPbOKtxJKcx+RKdKIEB8e
xObwcfHyksOzoiOavFRA+gczSdynRDe9fMXNL/G0qYS7Xc0a8GfkkTf4Uo1ZlTmv
a+ULMhD7TcibXVXqhQ2gY7JnXlRniDZgRl3F129aupLgRXzszt0D4xwfC+1ATUrt
tNA8Cgv1Kkz1b05Z/lavibPPlXVfwCAXvy9ZpZVjU3jqZZlZEOSiBtJolFVS2WCd
3UoyMA+u6Z39B9iFJ7h6fNpCOTpTGHSvuSuncER4qlo5TKZ47wbZhG2894tkTlWH
lD4Tkm68aO7k/dlLsV1TjNJCKbt0QdgTCS5JmQuRivdLePbxUdQFnY8BiOTMlgVP
elmNv9hBpNJHbSu/5NvyDBZW6YTU0+vcep7nbpnFwkzmwIq85ZK+NZn6oETNPreu
DpZrHz3jfPVkD0RyVQ5W3I1U5KtgFEGp9t9b87isgXES8CEyt32uBDa8J9oiVoFq
veZVwGMqOsMmVXSNQJVHrPcg8jwQ72j5tz8wDn1l7Sbt2qhswBA28fjCsGzwqJFj
U+9fU8m368kDU+2vQ9xcqdLOju6vHKy5aqkxGn7VaMKQuYLk8J5A0YovqGMMUmXO
rJ0x1xgRkxT8NJIvDIZCAzocGYytf9mDRBBcSTjXSKT77X/ZKy5E2r+gEzigD5Q5
gwwKjRfYycgTtHO4O17lLIxLbSXai/JJmG9PE3gZXyjSDP9pcsNvrXcBbu2TBV+h
eCmFwH0wNekqeraXaeHkvqV8myMMY6RkP6/pXm379zrhmp19eLcwvCmSVtCSZAmU
qQkcbkf3Y0zCQ0HezE361he/IVEe+HD7uSyJ/NyTeAy+o2KxETIEm9AKrztoV6y8
FfM5ZOEbSVuWiOrOa3JJEKTghN/QZux4ViFj9cKfIqti/yLWKAO+8xb3ABLMbHXE
mkyCo1wFQxx8wRcaO7K7zBr0DkKFcE4yRiJ0h42r+tM4L4nKR5fgADcZ/PNKQoFI
gujkEivXSj/p5bM2X5VTgAwCeQMiNDrmNfOVlXOPMWrMcMFZ10Rg219DFYenQrfc
NBvYYQxveZejHZrf0MVXEro39SOI7W+2SKX4LgmNio4Y6x6kcyFqHUgub+IJmrSl
RawOfni9KPwF5vcZxijWgQR2lXJbNR7Whj2W7H/n5ZipwtdPAj8s8x5ubgVlTyyh
gqpjWCc7USJih5Ey6+7e2XVmmKf8GRdRuZ1bW0P2aKpomPnYms5V6JRZ7/gz7gr/
7o+51nTPxlHV2sd3qS/iSLAAeoCOQ/9HCNgkz9Vu/xw8LAsWks3/d0+/eIh4+Ed0
yxndYHpwwYlnC2OSZgBmAWAuAj/Y8Hvs4GWwCKLRs9qozr+bunqUVecrV2jC+S6W
gzY7vglMxDOCMdOaXf9tHNBjANMo5Dt6svNsngbc/KHPxCu+rOQ5lddi0A4ZxOzp
cwCKbK0WP4WoMquz2wl6/KcK/mRAABZ0Uw975r/YmsK5DInZHoWfB5/CpKN9Cpfh
WMnjWNJcTHwjcUZpdXRIX00NuGml5UDvGRvwixKFBDvBHxwe0ae9YiBYQPo1qnAB
HftOJNEufQzDlHTppI2mj8adLXlArIMAJxKqxfsqIpkl0t/TDQ+10/aH3WkXFw8v
vvVrL1sdrQTuzLKfqprYNU+JPnrq24WnyDD1mgMK5v7PfEY39x77yRjU6pokaJKD
uXqVIm1+8cKxgWh3dAPO5sfwwf0cG1E4EfOUZN4JXSdpl2tvLsXn68GTCfle2z65
7/di5Y39ubP5yIUD/Iwj/f9n4Uq/+V3Sp/3WzWezWdHu+d/Kjiu7zeJjct0PpUgn
F3Kk5uYQDU9QT2QgT0NLmcFyqbL4BVbaekIjZTGYDxycDFPHc8zU8KjLi4j6uBlX
ZjZznwHWaO4ZFUR9u7aPtSLG+ngMBRbx5G3wnStscUttPWOQy0J5vsas1TLpD/ny
0R64QHne7Rsf16pQpbWqq7+po63YeX4TF8SWjsd6S2n+fiSlzqPT1CmCX7zmdipP
MF0VvQUx/Is4SNsd2BRVLjFdt8+I/QruoJPcaMcK7ooEttg8pA2hR0z/1UgiS5zD
7AhBg82MElbKyYrpPENF2Diq4jeDEz18FDTa0WLpVssS5obPPSfiQdLFFYGhpXmy
3O9KOldjhWRz952VLdKBQyCmTS/X3iPHW4kCbqzkjz7MX+8XV8emlclPOOn+2dSo
gtogII7x5E5N6uZzF0052Mg7HTMZ4bbUTMZ/+gxkKthUbIXDYgyCap8PUTLsp8jc
BT006NqucQmxVYYvNzBxcPbu8r2i8sgKKxDCKOBj4OA+QD5VuwJIa43LKUj6KB0F
ebyFO1URhzLUoayqEd4N6gHLSiXZVWWtN/NgjXonhcQ1P/YRjUarXs+eIjr6OfU+
by1N0WV2+fhkW9rI+g2LEdyA+xuNJiALOYrUjfO3W9XIWAZps+SwwNmWV+lC0x1q
DQqx9qHkC719Ri4rC+r5GAdxAte19bMgatl7XeDeZFMrMOOkFkMNogvxZZmRRI6M
17EBh/Lx33RonmiV40ILKuDwHVjV3w6TprIa53yUDAiCmjnPgTzcFEIybVzneqxu
2Ks92bXSUuJuOtga+3wEotJt8W4po7D50SzMgDI+3cYn9gQE/EWbenKuJKVZaMdE
i2RHfCL0J3b+LoT/NF5R4M4nShCD5wVTbnCWaM87t8v9JLkcPnoBtrVZhI5eG42i
XnCGGzUEd9VsMtu5nU/d4os7YvuJ97VtT7tB2ubA58O1GEU4+6yEssvdLo4Uloe2
+zaeltVWtkxAJ9QrA9FiaqmZLw/C5ofs2UaOpBtpOr07SrJfxXgsdNOZKmE0np25
HmvXfXfbxoYrb80Z0BBg83T90lZib9s31gv6Aya9SJY5AG/blpS66DNbmoQQDPkh
ozx1kWfAtDbcU7r4jEE2iVA6s1rj7UTq8pXVbgfDxxpcriMEmrn6FDOlCljMqLUa
D9Ci/tEUl7gsRHmez/FIf0M8DWseApF2f+UVWn/BlKSzA/2a/irgJ/8bi3GoV4re
jG93qfzZ5UH1W1MBS6vGW5UlnpG4X4eRbNIE2M6NUYkEd3nElGcKmoN5nin3VL8w
cbIRtQ0L+z/+dXmUev/Z6JTYsw6AXkJTQFUM2F62zDk52YJukY0J1f94F/7Batxn
ge6meZMcKU2KbgGWWI3YNeKfeVtpP1+wuoeMLl34p3PH0Mh4GvYwPthyvI7oP255
GOzRtXTERGz14WWnY3iUvp7UARDKqNmHoA8z12jzHRZYUhpSB+jWXX1j4byPPF4Q
KxT6jQp/KZO65OZCC1IZpT4C6FbEIgXrAAv7GHanIFiV8uG/q/mVW0TwRYY1AVhr
sY9St34ICZsjfLcBtf3YLPl7UIIFN/VAUmlj5rzdRzFL5g7eNoM4EAg2roRssfnD
nIhd2D8iik8PYxheDNy02lMT5m6BzDRpyumjWt1A2+7Mv+vWOvjpgryq5IWQeN0h
ZfGKlQ8LkQNOF151kV0m4z34tb1r51E0nF+DCHUaY3nu5gcCK2JJQC7YwnDH7FwC
km24MSeW5rjclViMmLfIFMABPYI1ngPuktZl1w1tjoRSFqbFkkORA8D418Z6Vcqr
lt8PE3mnEwVZ1hOFBBgLhhXXHphRtbuc23cMdSfuqXzrqD/BQPBKBQicGnSw5XvZ
rhZqc9x+stzNVYNHfhfqifaZvbmnvRGnqtonuH/fEDQWq9hOm8YK3a4Sh5tkX6YX
atZT6Si+74taoH9RE7pD5mXjDAevCQozRHWH+L15wSUEVla4PJuZldDdhjErYI+Y
oYsC6m9ClreomX5v1iCuHQdhSM19LRsyPj6zmTMpCmeeR1WuPCTbDkLmDiyyeJRI
tanWD+FFrzgeBp+6ULlEP1d/oZVpu7wWhSwZgtZbd246KopcIYgQTBdIgmKzJeZg
QrGoUOHt9ofOTZW3y6zagUWTTCZzoKl8XgjYmHwIn1Fr2V9XIqpt6QQaXwVHWFNo
38C24dxyFt5YfNvjqFZGRN+lvO6RWjfjjivPyPHhthZS0GmN2qOvUajc9xWkaizj
hPtDlggCF35dpIm9FBBqBx8CqStdKLfwIIe2XfxyzPSwUyyf7bbbuJfM4gILN8em
tnXu+nNC2It4RScxJoolobg4CcIswtUVQ0kAD+9k9ubwEiwH+j2QjVsZxUB+Ljbd
UvxPoi6p8JrvK+ZBC26biRfnF9NpAjWfyerFgYFRDWkWhMXNa/HJTi1wucG9/pV1
VJu0IL7X8Q986OIc9aXAZjsl3kI4KtdzNQuH9f5p2Ofdyx4ZSBz8iT6SxbEioxSj
zt63RjKTOd4eLNy3sZwPGSe651E3O1+ooJcLDdd2fbUlj7CERJDgLPC4hoZqNdTV
B/P+qif813AhrR5hrmrz1eIxqi7+Kpdj9MrPQjPRCQXwvy/YzXafSpce5eQ/MIyl
HyQT9i7xLr6jcBzlansLINXeMRio4cElZq5bIoaCTvTdnQNQtuSFj1rVF1lr3azG
IAc52FVCzjXGK+Vp7W2FGJmjzmzu8+pn/f21UJSx0btsygY0XYjPqyi0A4iFioYu
9NwhcNwf5BlvMMKO4M5r5mc293VA8XHFXIg1VsMr3I7NG5/PBtKNsNV3D6Cc0C4q
Pxd4LKIb2ykVykequm3N9GpMseLchUVhJFq8MRc5aGtOQiRYwlfo3HG1t40oA56l
w+vnBdwnm7AmUAZmZQ1WuYZ+XsxzQpA0p8aR34ZGUz1SIdKfHPJlOxTE1rWQBUkg
+edvy7GFoEeEWvae+qZoJfxOoK72Z64YBv82CfPE+3GLBy/p2kXDZQaNa1S9fXff
GJ6qCR50vb6iPXSkwVBRxtzZS7P+WltmKge55GZU7l6I4Doq1IX4jz+mtnK3R7bF
JwsYVFFQk8LMBYy7b+qs6C+Ft3OTVnKQnv7u6e9+J4aAGTMfGhjkRPn1zSN+P7Ht
RmVeEhka76ojA064++gU+eHRpUmIHSzmryvES7SF2aiupHUiWR2R+YM27mQ9ZUYu
DrlB3/+ikBTZtjWaLfzX4oJpM2mOvFSJQCjVrzxvYgQP6k2x1VYjc+MMR8N17p5u
1ZbikLmc4/TpnKFPtU76otL0UspTMjA2VMMosstYW/tv9v5Ipea0TjOHyvl4dIOq
7GaQYLDcXlF1QHiRCKNhcquPrbqjewL+uoGAPv4meGjNkGxD/tQQAhbcfbn3q96g
dR2kgfULJXLvUu7l21pLeILu9LqCNgoe8Yk1sdjNMRBw+lVW5ped4ZWvW8gKDhfG
WBFjkVMx/wmlqTc4ZL9V/sgP1A7hKeoIO5KiXcSWgB2A9Rh6W2VBjkDoHE+6QtmQ
POTIE+lj1tqYYEnd2DAZn4WTn5KQkb+fUBtpeLB3BLnn3Ihe7vPxinu9d5ReTPDd
muwgcngETlx+QKWAd0lzdkmh3KYXMueCZ0M95rKvajwj0qFgcbSXrM9GK/U2qM1L
mvx7rF+QL4WUB9k/whX93+vKPYYUrHsg65v1ac4nRYv3JI7fGMNlP4LHxiMh6/nK
CBYznYE2Jdtyh3MDM3KDRanmJzxSWmw1gq0+dGD9t686MJZZR7vtGNz90zW4puVk
qyZY4BIHea0WTPvP9IYzwnmH9LlqHwFCl70XkwiLgAlE3cD6CFR1ug5SzcuV4X4r
3F0MYyF8nN+eQZXWFk2jlBKk/UnHTrvsnyKmZrOT5aEDDcPP5v3+Xdy2nlbKryFU
82+SwWOGbSW4s8FFhzYlPeRlUnp0tBcrhuYNJSKdCS1O7k7+Q8cz2gJZWvuoLJ5o
3MblcvMSiAXqcvQ/77CoUtP3YzP4UG4uejzVrUc8+m99ZKH6jOsewrKwSvEWgcxJ
ZP05yb7DNfnv0eoHfNvm2ru+0QHDgT8fdtBDjxNmu/YK0slUjVTWEHoV2g3Be8xv
uFzjZJu3SfkSkjlHNatWCO2tT7qX+PgQ6MveRfrYYPaSMrPvot0G3rpWAswZ+r5b
3ltSEaMzSEe2OU2MgyoHfhu1VJqkRAiSMeKGIOyFNEKnkjJMLIEjhGoPUGE9jsJ6
5zOAi8iH+o37XsKl1YxOHL3ZPpXBqC8cEkCdO6rdrsQdJjsEqt1EjmWe917Wrp5z
fEqVkTrBt+e2Sxur8oRDy4NCxPVrzuC3yYPwkV4FHbstRo+4+BkVWrPkDex1z5jK
N1hf8Um2TuqQ120w2KNWG3Ge9TBzz+OpWESUxovE3iXTDO8HVMtoFD6XP1Yjlm9w
WUUwPqJMTYJl4U08VW19xSd1owyxYv4wf16FAD/Vqb0TGWVVrcfJFsPGwcR+TrDN
FB4onET3n66Wp/3ZEbwJZc2n+pHM+W+3RzKScBenzBLcBo8pcAkQ89ZcZc+jb6KY
Vrk6+BFmIsg33o0st9Hnrjsmw+MXVQZm26c6+hlBgu4JRe8NGBYdAzWtGmhgKzJG
UST/1JAWM+mGAZKpK3G8yyyM4IHMK8H3rsAply8xfHuxrbOt40TwFzD9/opKzb9C
PEhsbwrR/GD3afjuZR/C4Y/a63QYQ+19k0m2jldiJqrXoHguUdmDQkmfJlEOD5QS
4nAe0birloN7mHFfgthiBjnmHp0J9MiAiIVHKnZ+H8U9nu0qFHV0uP9MIAugGjna
EQkQnnJGEytiIT5fH430674ChCNWrfmdu2hc1jmdFp5ni9t1saTQBeyv/YQqjyOb
Csb8+GwN0TItfodfu8MNUCrILSk4CkodA4fzboe7aJZL9Iz4oi8ACAnK8ZLoAcwd
3F/Yhs/xj08ln3Uw5UB99LKauZx3WDQZYJkzkPLKFkQnHarzaMcswYhyX4qwqOy7
nY98dJaw2fnpb1Rwf7kSNNhZlUWinlZhj0pzz9gH8AJ79IF+u0wyg5H9kohskZ1/
6oMaKebPRY6BIneAv4LPMKd3ufoH4Rmo25oj9cDfl3YhY+1HjyIxJQbP3lOgD1DE
wZJoqpSbWjkQytG1t/kINBDr2UD2rQaVL5NSdKCprNavbYy/5Ui4PwI9dL8OoC/L
8c/nqwc2Onrn7H1BZrIAs7ol5cGNWPWyF9qVUZH72tNlguMTApzk/PVBPFT9nVOC
qIxWN4ldBFlSXEh6lkhrvWk5mEl5PxSKOkIwy5GUmDjRBZidfqR08x6Mp+bzFMnM
eTcUZSN0ORBdtLlbxRfgsg3JVwblsf6OXfV+HAYVGPvClUNIPsVwOz0yq84CHuIZ
b0zHvDgDejMB840AZhzEnw==
`pragma protect end_protected
