// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 15:05:48 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EqOEzQbz+m68eH9tjb/BR5RGnT8wN7TEshjv3dCuBZkoF6Ct6D4YYLazk45lihUT
CMxjwdv0i7lrBg5vHXyZVP+0UnN2TFEwyEtoNaESd/1a0ZXY9S4vwNXeTPPu3mzz
v7EPWT2EPTJvK7GM2nVrC89RXMLVe7kWjwfe/825GTs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
/6wlMIZ/49jjnkqhXPbgxmMLMLcmEJ3fSouic0x9XQQ2fAyr0tcl8J/M5xrynk16
atEgdQs44CvFN6lHtNn+cVGl6Vem4ZZjtrYrD1x9+E3YDwtR1Er35uBrZSy/IPvB
3hpC2UcApHOLMLof3EBTIiwe97oc3PhDWQzlSbcvh1DjwSHUCiwE84pzJl+BZI5N
Dhm0qmCiPx5/CWgyRdkRqvqWFzTgMYrL6iatgNPmR4PfV//H7VICw5FhfC+hq8Ls
nCfG8lDTu4/Rq6IjrFf5Aq31MEqATaZWRqe8fmSQpFIEtPoh11usfVN8Vtpl0xNU
HHvfsHOSmNZ7RE8sI/cdOTUcUwK318dBGYBUWkC5I7hS0qqz9XOYAxqb73OnrLAq
WA0Wm1zBpc/QgnZyh1UZBf2oaJbzgHUUSOP3A2LVUYwHfH5nyB+4WUG2ijYBS3TG
k7K+b9wQJsIhfME7KvjimmTdEcbxCZ/56KW+61fyAPTZA8827JbtbgdrOsANl6EH
A13u7QwV4ZWyIiYQO0p2aPIHMZwxjyzOMLEk3wtvj6Eyp6taid1VOVgS8B4Ayo0J
rHOn+qoqMdxV4KJwiXViKn9uVlH0XdPYVC8ggXI6BP4uQHHgxsGsEdBRgvaizlHN
orxkkINaDrCYy3uf6uMqhGfcjCHsfJU6SefWAKnrUqAoGkSBSInzR5cL71v14+TS
lF4+sklh6J7FuxoBtfG/x3R9c1dNfiFSzaEkflK/pW9UToLZjph6wZgpElBoNxfw
Zmo7APRPpiZv6s6B0Ok4G0FwD5285AsLt9EU5HK3B1v8GiTK32j40NqZAxln1UHl
ZFX0q0JKquzLxNNWH2uDy7m3fF/JhUJEj2r2Z/xn8TWOaTc4GGUXUIXrFQcj/njc
JZeR+2DBxswJ9mIAPATpf7JU9fRBSoD0QJlRDzcKSA1uQQM4v4A9hd6dbuGeRiHy
el95oj3OBGzhV6ZekfLUYIJICbqJZKkBtC4Vd2jXT7H5ihG5oQKT5uQkYWrKDZRU
UQkUgElL55eUQOHsdLWjPGtH1EjtWOFMBjbY1ld7782mGfyJqw+FxBdijMRc7biE
ghcivqleYbjypj9J0oKeZxy3ADbwijJ4xa+pLVeXUzC1XCXXEZm/LIBqplB+lTR0
eV4MmFfxBIfwUM8ZgAU/s050372xaqY5gwmWD2Ad3c01NDhLI4myNA+6jSPORyA/
+xk6RRWmIYWPj+0jFuO0IkUbB/QN3hbDh4NsogQQTWkOCrtcqw4PTwNF9lNRqrmt
QGZAaRGOor4Q+Dpzf2BdmODRjHlAse895zr3cKf61iXUvVO+SmmtXPcfqhuv65zq
eXSvUUp49AYxRHFMEEq3iwA3qbA1mvOsVvq/EKhEPRluiWypRU+hpOu0jZZv/8Kv
/WoD7IGZdoZVrPVPjXOP5P/8ZeTMIeZJuOJ2Q456QOAE3ycL/ckzl0sFT0pP3G+V
lAGjhBQyN1tDcMK8b6aoVg35953qKJPJWPSd/eyD7Z6ofmq0O1XrmNes6PthMLty
OpCmToD3mn2o7egdhudP30Vkydcuf7PYE3VbIf8ZBo2dx1vxaPeQ6oMltjvYl/px
X3o8EP0FfDpCTXe7XHTyy1eaiwaZPTAoPkBRGhJ0snhAXnzkJ1wu2P/Exh75Z1C/
F0dyC1lcqY/BuxPcK9EDOKVFAgvlUEseJK9KC8NAQvCiyXx5VooS8XTlrvmXU2j6
v6kSsWU4KLqmINyRYjjWBVdIgDyltpIgQwGHx1rWQUQJ86VRhJDvI13PSrlf2aL/
1nM9texmKZ9fHtv5axYGSCl5rvzusL1X2d9p1U5DuwoKWP0oQOgnknFmNR/J1Wq8
VG+4tWy8NFY11yOBYFdldzGRi06tVTihRascR80VMYy9IZxFqc0/lJmtHFK/EnGV
uUELzySH6SUgy10P5Xa5CalCRR058UwZssW3AROyz1scLtWmW4++fYI6Kn5wsJQ7
3zUkm6VmWOeTXmfsXjaALYvtaUwNnTB5iKXvBNvbZdXMGBVmmTnW9OaNOlBSqeUr
O0shvE8YFH9L/Kmh+iVLV6duTHLLuWKlcS1LYZyAzk+kRKc/XKjF2SBOzerxcBoh
2GuzOlgrN4NBCziFxFxp7nBk+CVPlCBuGGFsIfgQ06Gp0VS2/W1Ca0/dyiZF/qmt
sBk72UwaD5ubtQ4Q/QZ/8gb9iZqoVIcjbBtTGKKN249A9az2wqx1wFR0GWElWH0K
yqTS6wxhSFhMajDzDo1v6+v3bPp41n3x956kXaNxXy8naBZYbZmVjXw13+lu0WyP
xiHB/cnTd14266fep1uOEiYyCRBL999a3xoxp47pH3+KcxeN2QHtJbMoAwPboVh9
59Gj5f8YUOKSbTTImBOuJZ3bQbbKV1DVkwjzyuneMBd8z0kcEWGYoSBnt/io65ag
UXR710W10gtmMShHCSp8ZV8eJQxsko6S8b5Crdcxj+EgSjPcQ7Z/l7MUQTCygNlA
mL8ypDR8fgjV53ubmeGjyL/xi2AzJbwTTtwSwQYm9KrUn8RJnL5iFhPvbBSBHIis
QLf7R4nyP/4cUKSqsVEvjFwEcITQoYIPeEm3Vu/0D+L3NHI7nM7TmjC6Y3xT3peT
xx3maARRIvT4JRI/fD+VC5aW8ajNHtBAH8I9wACN0o2vSmWvGpHrEIWTdfxiuo/l
XUovNDySNCb9ktMR4z4KCYrFGGdmMl7W7LTpzcnkIA+yG+GPGq4N1xt7QvzTPyc4
TQ0uasRmhsOefznPKDBYBY4ehxVSVVnKPGIi9VWeumbSlxg59NQjcPWLdLWLyUz2
jP2nUR0dK0MyPdi+b/n7Sj81xFebH+lni78DS5zOvg8gHUrkQBiltq/1Wan52KRU
ybizQqBYnagPi/MTIEEYA6g2yRZ+boF0Csv804QEa3v4RJHVocMJjacpKDtaWTsb
B0wQHso6568xcOgyYgqoQ8J+Kwyw+o99dE/kZKP0sj1g7QNW33B3MTHC9rMksdEM
dtCSbRHOjOh9KrCUJb9xUlYfJZv4P5RchvPI5ShTGEP/gOAv19yLThDSk8HP0hv5
YWZTQ+RtRkMSSM+0u38eGRUsa4vER0jZl5/d6oY9Xhgfe4wYwHC73TCOLbiQTrGK
hWuhxzxfoAEAo+mg3cFJQqQCdv6Mj2Gadwn5n+QDpBYJpVQ7VytaUD+yH8nnPpzf
DA6m4IbSBMOUKZIvpRGDpVXHSd30WP/YrKMIZEwzfnI5dcGQCo3xsLZ6TPnbdqpY
muI0OQbWOgeq2puXBRVksjgbvvvkjTvGZU3PrPS1z02MpEIEkqp2+ICEh4lt8oSG
HJYIEr/oP1nhabEa8zbZXHHA+ORj1qMCV4KLyNI0gEpjTPA764VfJqQsIAFGDA3s
Bt+nhpkWo2X8vyh25DjxFIx31WgbjLZYPZv5ffNyQ9Uj4cxeTYdg1N4SRf6AkZM0
3Vkp9liyllqdAO1fqZ7saFsyD8805HDV/Wz467+2e4UVp8/9I3wqY8L06JTWH4rt
fMJv+nY1UH1EWhsZtxiJ8RgY7yPSGmiJLP79kpwnAT+b5REnOkFc5Rrf8/94hq88
COasLJb7GRRO9q1YzOGJFwbwx/VfZMnERV505FuhqGn0AhM61h6eHPrmS4KSRAum
cBbzguqJ4zbXLIKAIIbr/6zQmq3+37OGKA/+wkMuM1n/LuRT2mw5mJ4ZMgfNi2Cf
VXXLI6Z67F/Ibb3cTm7P2gi1HrKsEW9ZdXwuqh42u7yhTNfGKVPVmeWAI80fa+88
ALesgrPatKoAJ69/JyGmMiJ2dMvuIpw9xVSS6Iql1FZFPcx92Yl2+Kw81iyqdTaK
aO7Ww+9a0h9lue9V4PImU98mjdRCETnIOk7O79piSGlZtyylTMlYcfsiXBjze/o2
2P8vaIbGD3XqAvlo2ogFkd+8zFmWKjsMhnE541efNF/NSGX5dQ0YAoRKLHHqCqHu
eBXVOF1J3oGA/Vz25jH1S4EUbogUBmOC5p0/qbiHJp1LpMFL32SEwX75F2waGsCw
mxYlft/UC4G348jh59cpXA==
`pragma protect end_protected
