//------------------------------------------------------------
// Project: HYBRID_CONTROL
// Author: Nicola Zaupa
// Date: (2021/01/19) (23:11:22)
// File: tb_hybrid_control.v
//------------------------------------------------------------
// Description:
// testbench code to test the control behavior
//------------------------------------------------------------



`timescale 1 ns / 1 ps
//`default_nettype none


module tb_hybrid_control;

//=======================================================
//  REG/WIRE declarations
//=======================================================

reg     clk_main;
reg     clk_10;
reg     clk_100;
wire    w_sigma;
wire    w_sigma_delay;
wire    w_sigma_delay_2;
reg [13:0] jump;
reg [13:0] SIGNAL_A;
reg [13:0] SIGNAL_B;

//=======================================================
//  Structural coding
//=======================================================
hybrid_control HC_inst(
   .o_sigma( w_sigma ),  //
   .o_debug(  ),       //
   .i_clock(clk_100),   //
   .i_RESET( reset ),    //
   .i_vC( SIGNAL_A ),       //
   .i_iC( SIGNAL_B ),       //
   .i_theta( 32'sd236 ) // 3/4 pi
);

hybrid_control_half HC_half_inst(
   .o_sigma(  ),  //
   .o_debug(  ),       //
   .i_clock(clk_100),   //
   .i_RESET( reset ),    //
   .i_vC( SIGNAL_A ),       //
   .i_iC( SIGNAL_B ),       //
   .i_theta( 32'sd236 ) // 3/4 pi
);

dead_time dead_time_inst(
   .o_signal( w_sigma_delay ),     // output switching variable
   .i_clock( clk_10 ),     // for sequential behavior
   .i_signal( w_sigma ),
   .deadtime( 10'd10 )
);

dead_time dead_time_2_inst(
   .o_signal( w_sigma_delay_2 ),     // output switching variable
   .i_clock( clk_10 ),     // for sequential behavior
   .i_signal( ~w_sigma ),
   .deadtime( 10'd10 )
);

always
   begin //300MHz
      clk_main = 1'b1;
      #1.666
      clk_main = 1'b0;
      #1.666;
end

always
   begin //10MHz
      clk_10 = 1'b1;
      #50
      clk_10 = 1'b0;
      #50;
end

always
   begin //100MHz
      clk_100 = 1'b1;
      #5
      clk_100 = 1'b0;
      #5;
end


initial
begin
// Data from SRC simulation in Simulink
// frequency ADC: 1.000000e+01 MSPS

SIGNAL_A = 14'b00000000000000;
SIGNAL_B = 14'b00000000000000;
#100;
SIGNAL_A = 14'b00000000000000;
SIGNAL_B = 14'b00000000110000;
#100;
SIGNAL_A = 14'b00000000000010;
SIGNAL_B = 14'b00000001110000;
#100;
SIGNAL_A = 14'b00000000000111;
SIGNAL_B = 14'b00000010101111;
#100;
SIGNAL_A = 14'b00000000001101;
SIGNAL_B = 14'b00000011101110;
#100;
SIGNAL_A = 14'b00000000010101;
SIGNAL_B = 14'b00000100101011;
#100;
SIGNAL_A = 14'b00000000011111;
SIGNAL_B = 14'b00000101101000;
#100;
SIGNAL_A = 14'b00000000101011;
SIGNAL_B = 14'b00000110100100;
#100;
SIGNAL_A = 14'b00000000111000;
SIGNAL_B = 14'b00000111011111;
#100;
SIGNAL_A = 14'b00000001000111;
SIGNAL_B = 14'b00001000011000;
#100;
SIGNAL_A = 14'b00000001011000;
SIGNAL_B = 14'b00001001010001;
#100;
SIGNAL_A = 14'b00000001101011;
SIGNAL_B = 14'b00001010001001;
#100;
SIGNAL_A = 14'b00000001111111;
SIGNAL_B = 14'b00001010111111;
#100;
SIGNAL_A = 14'b00000010010101;
SIGNAL_B = 14'b00001011110100;
#100;
SIGNAL_A = 14'b00000010101101;
SIGNAL_B = 14'b00001100101000;
#100;
SIGNAL_A = 14'b00000011000110;
SIGNAL_B = 14'b00001101011010;
#100;
SIGNAL_A = 14'b00000011100000;
SIGNAL_B = 14'b00001110001011;
#100;
SIGNAL_A = 14'b00000011111100;
SIGNAL_B = 14'b00001110111011;
#100;
SIGNAL_A = 14'b00000100011010;
SIGNAL_B = 14'b00001111101010;
#100;
SIGNAL_A = 14'b00000100111000;
SIGNAL_B = 14'b00010000010110;
#100;
SIGNAL_A = 14'b00000101011000;
SIGNAL_B = 14'b00010001000010;
#100;
SIGNAL_A = 14'b00000101111010;
SIGNAL_B = 14'b00010001101100;
#100;
SIGNAL_A = 14'b00000110011100;
SIGNAL_B = 14'b00010010010100;
#100;
SIGNAL_A = 14'b00000111000000;
SIGNAL_B = 14'b00010010111011;
#100;
SIGNAL_A = 14'b00000111100101;
SIGNAL_B = 14'b00010011100000;
#100;
SIGNAL_A = 14'b00001000001011;
SIGNAL_B = 14'b00010100000100;
#100;
SIGNAL_A = 14'b00001000110010;
SIGNAL_B = 14'b00010100100110;
#100;
SIGNAL_A = 14'b00001001011010;
SIGNAL_B = 14'b00010101000111;
#100;
SIGNAL_A = 14'b00001010000011;
SIGNAL_B = 14'b00010101100101;
#100;
SIGNAL_A = 14'b00001010101101;
SIGNAL_B = 14'b00010110000011;
#100;
SIGNAL_A = 14'b00001011011000;
SIGNAL_B = 14'b00010110011110;
#100;
SIGNAL_A = 14'b00001100000011;
SIGNAL_B = 14'b00010110111000;
#100;
SIGNAL_A = 14'b00001100110000;
SIGNAL_B = 14'b00010111010000;
#100;
SIGNAL_A = 14'b00001101011101;
SIGNAL_B = 14'b00010111100110;
#100;
SIGNAL_A = 14'b00001110001010;
SIGNAL_B = 14'b00010111111011;
#100;
SIGNAL_A = 14'b00001110111000;
SIGNAL_B = 14'b00011000001110;
#100;
SIGNAL_A = 14'b00001111100111;
SIGNAL_B = 14'b00011000011111;
#100;
SIGNAL_A = 14'b00010000010110;
SIGNAL_B = 14'b00011000101110;
#100;
SIGNAL_A = 14'b00010001000110;
SIGNAL_B = 14'b00011000111100;
#100;
SIGNAL_A = 14'b00010001110110;
SIGNAL_B = 14'b00011001001000;
#100;
SIGNAL_A = 14'b00010010100111;
SIGNAL_B = 14'b00011001010011;
#100;
SIGNAL_A = 14'b00010011010111;
SIGNAL_B = 14'b00011001011011;
#100;
SIGNAL_A = 14'b00010100001000;
SIGNAL_B = 14'b00011001100010;
#100;
SIGNAL_A = 14'b00010100111001;
SIGNAL_B = 14'b00011001101000;
#100;
SIGNAL_A = 14'b00010101101011;
SIGNAL_B = 14'b00011001101011;
#100;
SIGNAL_A = 14'b00010110011100;
SIGNAL_B = 14'b00011001101101;
#100;
SIGNAL_A = 14'b00010111001101;
SIGNAL_B = 14'b00011001101110;
#100;
SIGNAL_A = 14'b00010111111111;
SIGNAL_B = 14'b00011001101100;
#100;
SIGNAL_A = 14'b00011000110000;
SIGNAL_B = 14'b00011001101010;
#100;
SIGNAL_A = 14'b00011001100001;
SIGNAL_B = 14'b00011001100101;
#100;
SIGNAL_A = 14'b00011010010010;
SIGNAL_B = 14'b00011001011111;
#100;
SIGNAL_A = 14'b00011011000011;
SIGNAL_B = 14'b00011001011000;
#100;
SIGNAL_A = 14'b00011011110100;
SIGNAL_B = 14'b00011001001110;
#100;
SIGNAL_A = 14'b00011100100100;
SIGNAL_B = 14'b00011001000100;
#100;
SIGNAL_A = 14'b00011101010100;
SIGNAL_B = 14'b00011000111000;
#100;
SIGNAL_A = 14'b00011110000100;
SIGNAL_B = 14'b00011000101010;
#100;
SIGNAL_A = 14'b00011110110011;
SIGNAL_B = 14'b00011000011011;
#100;
SIGNAL_A = 14'b00011111100001;
SIGNAL_B = 14'b00011000001011;
#100;
SIGNAL_A = 14'b00100000010000;
SIGNAL_B = 14'b00010111111001;
#100;
SIGNAL_A = 14'b00100000111101;
SIGNAL_B = 14'b00010111100110;
#100;
SIGNAL_A = 14'b00100001101010;
SIGNAL_B = 14'b00010111010010;
#100;
SIGNAL_A = 14'b00100010010111;
SIGNAL_B = 14'b00010110111100;
#100;
SIGNAL_A = 14'b00100011000010;
SIGNAL_B = 14'b00010110100101;
#100;
SIGNAL_A = 14'b00100011101101;
SIGNAL_B = 14'b00010110001101;
#100;
SIGNAL_A = 14'b00100100011000;
SIGNAL_B = 14'b00010101110100;
#100;
SIGNAL_A = 14'b00100101000001;
SIGNAL_B = 14'b00010101011010;
#100;
SIGNAL_A = 14'b00100101101010;
SIGNAL_B = 14'b00010100111110;
#100;
SIGNAL_A = 14'b00100110010010;
SIGNAL_B = 14'b00010100100010;
#100;
SIGNAL_A = 14'b00100110111001;
SIGNAL_B = 14'b00010100000100;
#100;
SIGNAL_A = 14'b00100111011111;
SIGNAL_B = 14'b00010011100110;
#100;
SIGNAL_A = 14'b00101000000100;
SIGNAL_B = 14'b00010011000110;
#100;
SIGNAL_A = 14'b00101000101000;
SIGNAL_B = 14'b00010010100110;
#100;
SIGNAL_A = 14'b00101001001011;
SIGNAL_B = 14'b00010010000101;
#100;
SIGNAL_A = 14'b00101001101110;
SIGNAL_B = 14'b00010001100011;
#100;
SIGNAL_A = 14'b00101010001111;
SIGNAL_B = 14'b00010001000000;
#100;
SIGNAL_A = 14'b00101010101111;
SIGNAL_B = 14'b00010000011101;
#100;
SIGNAL_A = 14'b00101011001110;
SIGNAL_B = 14'b00001111111001;
#100;
SIGNAL_A = 14'b00101011101100;
SIGNAL_B = 14'b00001111010100;
#100;
SIGNAL_A = 14'b00101100001001;
SIGNAL_B = 14'b00001110101110;
#100;
SIGNAL_A = 14'b00101100011100;
SIGNAL_B = 14'b00001110001100;
#100;
SIGNAL_A = 14'b00101100110101;
SIGNAL_B = 14'b00001011100100;
#100;
SIGNAL_A = 14'b00101101001000;
SIGNAL_B = 14'b00001000111110;
#100;
SIGNAL_A = 14'b00101101010111;
SIGNAL_B = 14'b00000110011001;
#100;
SIGNAL_A = 14'b00101101100001;
SIGNAL_B = 14'b00000011110101;
#100;
SIGNAL_A = 14'b00101101100110;
SIGNAL_B = 14'b00000001010010;
#100;
SIGNAL_A = 14'b00101101100110;
SIGNAL_B = 14'b11111110110010;
#100;
SIGNAL_A = 14'b00101101100001;
SIGNAL_B = 14'b11111100010010;
#100;
SIGNAL_A = 14'b00101101011000;
SIGNAL_B = 14'b11111001110100;
#100;
SIGNAL_A = 14'b00101101001001;
SIGNAL_B = 14'b11110111011000;
#100;
SIGNAL_A = 14'b00101100110110;
SIGNAL_B = 14'b11110100111111;
#100;
SIGNAL_A = 14'b00101100011111;
SIGNAL_B = 14'b11110010100111;
#100;
SIGNAL_A = 14'b00101100000011;
SIGNAL_B = 14'b11110000010010;
#100;
SIGNAL_A = 14'b00101011100011;
SIGNAL_B = 14'b11101101111111;
#100;
SIGNAL_A = 14'b00101010111110;
SIGNAL_B = 14'b11101011101111;
#100;
SIGNAL_A = 14'b00101010010101;
SIGNAL_B = 14'b11101001100010;
#100;
SIGNAL_A = 14'b00101001101000;
SIGNAL_B = 14'b11100111010111;
#100;
SIGNAL_A = 14'b00101000110110;
SIGNAL_B = 14'b11100101001111;
#100;
SIGNAL_A = 14'b00101000000001;
SIGNAL_B = 14'b11100011001011;
#100;
SIGNAL_A = 14'b00100111001000;
SIGNAL_B = 14'b11100001001001;
#100;
SIGNAL_A = 14'b00100110001010;
SIGNAL_B = 14'b11011111001011;
#100;
SIGNAL_A = 14'b00100101001001;
SIGNAL_B = 14'b11011101010000;
#100;
SIGNAL_A = 14'b00100100000101;
SIGNAL_B = 14'b11011011011000;
#100;
SIGNAL_A = 14'b00100010111101;
SIGNAL_B = 14'b11011001100100;
#100;
SIGNAL_A = 14'b00100001110001;
SIGNAL_B = 14'b11010111110100;
#100;
SIGNAL_A = 14'b00100000100010;
SIGNAL_B = 14'b11010110000111;
#100;
SIGNAL_A = 14'b00011111010000;
SIGNAL_B = 14'b11010100011101;
#100;
SIGNAL_A = 14'b00011101111011;
SIGNAL_B = 14'b11010010111000;
#100;
SIGNAL_A = 14'b00011100100011;
SIGNAL_B = 14'b11010001010110;
#100;
SIGNAL_A = 14'b00011011001000;
SIGNAL_B = 14'b11001111111001;
#100;
SIGNAL_A = 14'b00011001101010;
SIGNAL_B = 14'b11001110011111;
#100;
SIGNAL_A = 14'b00011000001010;
SIGNAL_B = 14'b11001101001001;
#100;
SIGNAL_A = 14'b00010110100111;
SIGNAL_B = 14'b11001011111000;
#100;
SIGNAL_A = 14'b00010101000010;
SIGNAL_B = 14'b11001010101010;
#100;
SIGNAL_A = 14'b00010011011010;
SIGNAL_B = 14'b11001001100001;
#100;
SIGNAL_A = 14'b00010001110001;
SIGNAL_B = 14'b11001000011011;
#100;
SIGNAL_A = 14'b00010000000101;
SIGNAL_B = 14'b11000111011010;
#100;
SIGNAL_A = 14'b00001110010111;
SIGNAL_B = 14'b11000110011101;
#100;
SIGNAL_A = 14'b00001100101000;
SIGNAL_B = 14'b11000101100101;
#100;
SIGNAL_A = 14'b00001010110111;
SIGNAL_B = 14'b11000100110000;
#100;
SIGNAL_A = 14'b00001001000101;
SIGNAL_B = 14'b11000100000000;
#100;
SIGNAL_A = 14'b00000111010001;
SIGNAL_B = 14'b11000011010100;
#100;
SIGNAL_A = 14'b00000101011100;
SIGNAL_B = 14'b11000010101101;
#100;
SIGNAL_A = 14'b00000011100101;
SIGNAL_B = 14'b11000010001001;
#100;
SIGNAL_A = 14'b00000001101110;
SIGNAL_B = 14'b11000001101010;
#100;
SIGNAL_A = 14'b11111111110111;
SIGNAL_B = 14'b11000001001111;
#100;
SIGNAL_A = 14'b11111101111110;
SIGNAL_B = 14'b11000000111001;
#100;
SIGNAL_A = 14'b11111100000101;
SIGNAL_B = 14'b11000000100110;
#100;
SIGNAL_A = 14'b11111010001011;
SIGNAL_B = 14'b11000000011000;
#100;
SIGNAL_A = 14'b11111000010000;
SIGNAL_B = 14'b11000000001110;
#100;
SIGNAL_A = 14'b11110110010110;
SIGNAL_B = 14'b11000000001000;
#100;
SIGNAL_A = 14'b11110100011011;
SIGNAL_B = 14'b11000000000110;
#100;
SIGNAL_A = 14'b11110010100000;
SIGNAL_B = 14'b11000000001000;
#100;
SIGNAL_A = 14'b11110000100110;
SIGNAL_B = 14'b11000000001110;
#100;
SIGNAL_A = 14'b11101110101011;
SIGNAL_B = 14'b11000000011000;
#100;
SIGNAL_A = 14'b11101100110001;
SIGNAL_B = 14'b11000000100110;
#100;
SIGNAL_A = 14'b11101010111000;
SIGNAL_B = 14'b11000000111000;
#100;
SIGNAL_A = 14'b11101000111111;
SIGNAL_B = 14'b11000001001110;
#100;
SIGNAL_A = 14'b11100111000111;
SIGNAL_B = 14'b11000001100111;
#100;
SIGNAL_A = 14'b11100101001111;
SIGNAL_B = 14'b11000010000100;
#100;
SIGNAL_A = 14'b11100011011001;
SIGNAL_B = 14'b11000010100101;
#100;
SIGNAL_A = 14'b11100001100011;
SIGNAL_B = 14'b11000011001001;
#100;
SIGNAL_A = 14'b11011111101111;
SIGNAL_B = 14'b11000011110001;
#100;
SIGNAL_A = 14'b11011101111100;
SIGNAL_B = 14'b11000100011100;
#100;
SIGNAL_A = 14'b11011100001010;
SIGNAL_B = 14'b11000101001010;
#100;
SIGNAL_A = 14'b11011010011010;
SIGNAL_B = 14'b11000101111100;
#100;
SIGNAL_A = 14'b11011000101100;
SIGNAL_B = 14'b11000110110001;
#100;
SIGNAL_A = 14'b11010110111110;
SIGNAL_B = 14'b11000111101001;
#100;
SIGNAL_A = 14'b11010101010011;
SIGNAL_B = 14'b11001000100100;
#100;
SIGNAL_A = 14'b11010011101010;
SIGNAL_B = 14'b11001001100010;
#100;
SIGNAL_A = 14'b11010010000010;
SIGNAL_B = 14'b11001010100011;
#100;
SIGNAL_A = 14'b11010000011100;
SIGNAL_B = 14'b11001011100110;
#100;
SIGNAL_A = 14'b11001110111001;
SIGNAL_B = 14'b11001100101100;
#100;
SIGNAL_A = 14'b11001101010111;
SIGNAL_B = 14'b11001101110101;
#100;
SIGNAL_A = 14'b11001011111000;
SIGNAL_B = 14'b11001111000000;
#100;
SIGNAL_A = 14'b11001010011011;
SIGNAL_B = 14'b11010000001101;
#100;
SIGNAL_A = 14'b11001001000000;
SIGNAL_B = 14'b11010001011101;
#100;
SIGNAL_A = 14'b11000111101000;
SIGNAL_B = 14'b11010010101111;
#100;
SIGNAL_A = 14'b11000110010011;
SIGNAL_B = 14'b11010100000011;
#100;
SIGNAL_A = 14'b11000101000000;
SIGNAL_B = 14'b11010101011001;
#100;
SIGNAL_A = 14'b11000011101111;
SIGNAL_B = 14'b11010110110000;
#100;
SIGNAL_A = 14'b11000010100001;
SIGNAL_B = 14'b11011000001010;
#100;
SIGNAL_A = 14'b11000001010110;
SIGNAL_B = 14'b11011001100101;
#100;
SIGNAL_A = 14'b11000000001110;
SIGNAL_B = 14'b11011011000001;
#100;
SIGNAL_A = 14'b10111111010001;
SIGNAL_B = 14'b11011100010011;
#100;
SIGNAL_A = 14'b10111110110010;
SIGNAL_B = 14'b11011101111010;
#100;
SIGNAL_A = 14'b10111101110100;
SIGNAL_B = 14'b11100001011011;
#100;
SIGNAL_A = 14'b10111100111100;
SIGNAL_B = 14'b11100100111010;
#100;
SIGNAL_A = 14'b10111100001100;
SIGNAL_B = 14'b11101000011010;
#100;
SIGNAL_A = 14'b10111011100010;
SIGNAL_B = 14'b11101011111001;
#100;
SIGNAL_A = 14'b10111010111110;
SIGNAL_B = 14'b11101111010110;
#100;
SIGNAL_A = 14'b10111010100010;
SIGNAL_B = 14'b11110010110011;
#100;
SIGNAL_A = 14'b10111010001100;
SIGNAL_B = 14'b11110110001110;
#100;
SIGNAL_A = 14'b10111001111100;
SIGNAL_B = 14'b11111001101000;
#100;
SIGNAL_A = 14'b10111001110011;
SIGNAL_B = 14'b11111101000000;
#100;
SIGNAL_A = 14'b10111001110000;
SIGNAL_B = 14'b00000000010101;
#100;
SIGNAL_A = 14'b10111001110100;
SIGNAL_B = 14'b00000011101001;
#100;
SIGNAL_A = 14'b10111001111110;
SIGNAL_B = 14'b00000110111011;
#100;
SIGNAL_A = 14'b10111010001111;
SIGNAL_B = 14'b00001010001010;
#100;
SIGNAL_A = 14'b10111010100101;
SIGNAL_B = 14'b00001101010110;
#100;
SIGNAL_A = 14'b10111011000010;
SIGNAL_B = 14'b00010000100000;
#100;
SIGNAL_A = 14'b10111011100101;
SIGNAL_B = 14'b00010011100111;
#100;
SIGNAL_A = 14'b10111100001101;
SIGNAL_B = 14'b00010110101010;
#100;
SIGNAL_A = 14'b10111100111100;
SIGNAL_B = 14'b00011001101010;
#100;
SIGNAL_A = 14'b10111101110000;
SIGNAL_B = 14'b00011100100110;
#100;
SIGNAL_A = 14'b10111110101010;
SIGNAL_B = 14'b00011111011111;
#100;
SIGNAL_A = 14'b10111111101001;
SIGNAL_B = 14'b00100010010100;
#100;
SIGNAL_A = 14'b11000000101101;
SIGNAL_B = 14'b00100101000101;
#100;
SIGNAL_A = 14'b11000001110111;
SIGNAL_B = 14'b00100111110010;
#100;
SIGNAL_A = 14'b11000011000110;
SIGNAL_B = 14'b00101010011011;
#100;
SIGNAL_A = 14'b11000100011010;
SIGNAL_B = 14'b00101101000000;
#100;
SIGNAL_A = 14'b11000101110011;
SIGNAL_B = 14'b00101111100000;
#100;
SIGNAL_A = 14'b11000111010000;
SIGNAL_B = 14'b00110001111011;
#100;
SIGNAL_A = 14'b11001000110011;
SIGNAL_B = 14'b00110100010010;
#100;
SIGNAL_A = 14'b11001010011001;
SIGNAL_B = 14'b00110110100100;
#100;
SIGNAL_A = 14'b11001100000100;
SIGNAL_B = 14'b00111000110001;
#100;
SIGNAL_A = 14'b11001101110011;
SIGNAL_B = 14'b00111010111001;
#100;
SIGNAL_A = 14'b11001111100110;
SIGNAL_B = 14'b00111100111100;
#100;
SIGNAL_A = 14'b11010001011101;
SIGNAL_B = 14'b00111110111010;
#100;
SIGNAL_A = 14'b11010011011000;
SIGNAL_B = 14'b01000000110011;
#100;
SIGNAL_A = 14'b11010101010110;
SIGNAL_B = 14'b01000010100110;
#100;
SIGNAL_A = 14'b11010111010111;
SIGNAL_B = 14'b01000100010100;
#100;
SIGNAL_A = 14'b11011001011100;
SIGNAL_B = 14'b01000101111101;
#100;
SIGNAL_A = 14'b11011011100100;
SIGNAL_B = 14'b01000111100000;
#100;
SIGNAL_A = 14'b11011101101111;
SIGNAL_B = 14'b01001000111110;
#100;
SIGNAL_A = 14'b11011111111100;
SIGNAL_B = 14'b01001010010110;
#100;
SIGNAL_A = 14'b11100010001100;
SIGNAL_B = 14'b01001011101001;
#100;
SIGNAL_A = 14'b11100100011111;
SIGNAL_B = 14'b01001100110110;
#100;
SIGNAL_A = 14'b11100110110011;
SIGNAL_B = 14'b01001101111110;
#100;
SIGNAL_A = 14'b11101001001010;
SIGNAL_B = 14'b01001111000000;
#100;
SIGNAL_A = 14'b11101011100011;
SIGNAL_B = 14'b01001111111100;
#100;
SIGNAL_A = 14'b11101101111101;
SIGNAL_B = 14'b01010000110011;
#100;
SIGNAL_A = 14'b11110000011001;
SIGNAL_B = 14'b01010001100100;
#100;
SIGNAL_A = 14'b11110010110110;
SIGNAL_B = 14'b01010010001111;
#100;
SIGNAL_A = 14'b11110101010101;
SIGNAL_B = 14'b01010010110101;
#100;
SIGNAL_A = 14'b11110111110100;
SIGNAL_B = 14'b01010011010101;
#100;
SIGNAL_A = 14'b11111010010101;
SIGNAL_B = 14'b01010011101111;
#100;
SIGNAL_A = 14'b11111100110110;
SIGNAL_B = 14'b01010100000100;
#100;
SIGNAL_A = 14'b11111111010111;
SIGNAL_B = 14'b01010100010100;
#100;
SIGNAL_A = 14'b00000001111000;
SIGNAL_B = 14'b01010100011110;
#100;
SIGNAL_A = 14'b00000100011011;
SIGNAL_B = 14'b01010100100011;
#100;
SIGNAL_A = 14'b00000110111101;
SIGNAL_B = 14'b01010100100010;
#100;
SIGNAL_A = 14'b00001001011111;
SIGNAL_B = 14'b01010100011100;
#100;
SIGNAL_A = 14'b00001100000001;
SIGNAL_B = 14'b01010100010001;
#100;
SIGNAL_A = 14'b00001110100011;
SIGNAL_B = 14'b01010100000000;
#100;
SIGNAL_A = 14'b00010001000100;
SIGNAL_B = 14'b01010011101011;
#100;
SIGNAL_A = 14'b00010011100100;
SIGNAL_B = 14'b01010011010000;
#100;
SIGNAL_A = 14'b00010110000011;
SIGNAL_B = 14'b01010010110000;
#100;
SIGNAL_A = 14'b00011000100010;
SIGNAL_B = 14'b01010010001100;
#100;
SIGNAL_A = 14'b00011010111111;
SIGNAL_B = 14'b01010001100010;
#100;
SIGNAL_A = 14'b00011101011011;
SIGNAL_B = 14'b01010000110100;
#100;
SIGNAL_A = 14'b00011111110101;
SIGNAL_B = 14'b01010000000001;
#100;
SIGNAL_A = 14'b00100010001110;
SIGNAL_B = 14'b01001111001010;
#100;
SIGNAL_A = 14'b00100100100101;
SIGNAL_B = 14'b01001110001110;
#100;
SIGNAL_A = 14'b00100110111010;
SIGNAL_B = 14'b01001101001110;
#100;
SIGNAL_A = 14'b00101001001110;
SIGNAL_B = 14'b01001100001010;
#100;
SIGNAL_A = 14'b00101011011111;
SIGNAL_B = 14'b01001011000001;
#100;
SIGNAL_A = 14'b00101101101110;
SIGNAL_B = 14'b01001001110101;
#100;
SIGNAL_A = 14'b00101111111010;
SIGNAL_B = 14'b01001000100100;
#100;
SIGNAL_A = 14'b00110010000100;
SIGNAL_B = 14'b01000111010000;
#100;
SIGNAL_A = 14'b00110100001100;
SIGNAL_B = 14'b01000101111000;
#100;
SIGNAL_A = 14'b00110110010001;
SIGNAL_B = 14'b01000100011101;
#100;
SIGNAL_A = 14'b00111000010011;
SIGNAL_B = 14'b01000010111110;
#100;
SIGNAL_A = 14'b00111010010010;
SIGNAL_B = 14'b01000001011100;
#100;
SIGNAL_A = 14'b00111100001110;
SIGNAL_B = 14'b00111111110110;
#100;
SIGNAL_A = 14'b00111110000111;
SIGNAL_B = 14'b00111110001110;
#100;
SIGNAL_A = 14'b00111111111101;
SIGNAL_B = 14'b00111100100011;
#100;
SIGNAL_A = 14'b01000001110000;
SIGNAL_B = 14'b00111010110101;
#100;
SIGNAL_A = 14'b01000011011111;
SIGNAL_B = 14'b00111001000100;
#100;
SIGNAL_A = 14'b01000101001011;
SIGNAL_B = 14'b00110111010001;
#100;
SIGNAL_A = 14'b01000110110011;
SIGNAL_B = 14'b00110101011100;
#100;
SIGNAL_A = 14'b01001000011000;
SIGNAL_B = 14'b00110011100100;
#100;
SIGNAL_A = 14'b01001001111001;
SIGNAL_B = 14'b00110001101011;
#100;
SIGNAL_A = 14'b01001011010111;
SIGNAL_B = 14'b00101111101111;
#100;
SIGNAL_A = 14'b01001011111000;
SIGNAL_B = 14'b00101110110100;
#100;
SIGNAL_A = 14'b01001101001110;
SIGNAL_B = 14'b00101010110101;
#100;
SIGNAL_A = 14'b01001110011101;
SIGNAL_B = 14'b00100110110110;
#100;
SIGNAL_A = 14'b01001111100011;
SIGNAL_B = 14'b00100010110110;
#100;
SIGNAL_A = 14'b01010000100011;
SIGNAL_B = 14'b00011110111000;
#100;
SIGNAL_A = 14'b01010001011010;
SIGNAL_B = 14'b00011010111001;
#100;
SIGNAL_A = 14'b01010010001010;
SIGNAL_B = 14'b00010110111100;
#100;
SIGNAL_A = 14'b01010010110010;
SIGNAL_B = 14'b00010010111111;
#100;
SIGNAL_A = 14'b01010011010011;
SIGNAL_B = 14'b00001111000100;
#100;
SIGNAL_A = 14'b01010011101100;
SIGNAL_B = 14'b00001011001011;
#100;
SIGNAL_A = 14'b01010011111110;
SIGNAL_B = 14'b00000111010011;
#100;
SIGNAL_A = 14'b01010100001000;
SIGNAL_B = 14'b00000011011101;
#100;
SIGNAL_A = 14'b01010100001011;
SIGNAL_B = 14'b11111111101010;
#100;
SIGNAL_A = 14'b01010100000111;
SIGNAL_B = 14'b11111011111001;
#100;
SIGNAL_A = 14'b01010011111011;
SIGNAL_B = 14'b11111000001011;
#100;
SIGNAL_A = 14'b01010011101001;
SIGNAL_B = 14'b11110100011111;
#100;
SIGNAL_A = 14'b01010011001111;
SIGNAL_B = 14'b11110000110110;
#100;
SIGNAL_A = 14'b01010010101111;
SIGNAL_B = 14'b11101101010001;
#100;
SIGNAL_A = 14'b01010010000111;
SIGNAL_B = 14'b11101001101111;
#100;
SIGNAL_A = 14'b01010001011001;
SIGNAL_B = 14'b11100110010000;
#100;
SIGNAL_A = 14'b01010000100100;
SIGNAL_B = 14'b11100010110110;
#100;
SIGNAL_A = 14'b01001111101001;
SIGNAL_B = 14'b11011111011111;
#100;
SIGNAL_A = 14'b01001110100111;
SIGNAL_B = 14'b11011100001101;
#100;
SIGNAL_A = 14'b01001101100000;
SIGNAL_B = 14'b11011000111111;
#100;
SIGNAL_A = 14'b01001100010010;
SIGNAL_B = 14'b11010101110101;
#100;
SIGNAL_A = 14'b01001010111110;
SIGNAL_B = 14'b11010010110000;
#100;
SIGNAL_A = 14'b01001001100100;
SIGNAL_B = 14'b11001111110000;
#100;
SIGNAL_A = 14'b01001000000100;
SIGNAL_B = 14'b11001100110101;
#100;
SIGNAL_A = 14'b01000110011111;
SIGNAL_B = 14'b11001001111111;
#100;
SIGNAL_A = 14'b01000100110101;
SIGNAL_B = 14'b11000111001110;
#100;
SIGNAL_A = 14'b01000011000101;
SIGNAL_B = 14'b11000100100010;
#100;
SIGNAL_A = 14'b01000001010001;
SIGNAL_B = 14'b11000001111100;
#100;
SIGNAL_A = 14'b00111111010111;
SIGNAL_B = 14'b10111111011100;
#100;
SIGNAL_A = 14'b00111101011001;
SIGNAL_B = 14'b10111101000001;
#100;
SIGNAL_A = 14'b00111011010110;
SIGNAL_B = 14'b10111010101011;
#100;
SIGNAL_A = 14'b00111001001111;
SIGNAL_B = 14'b10111000011100;
#100;
SIGNAL_A = 14'b00110111000011;
SIGNAL_B = 14'b10110110010011;
#100;
SIGNAL_A = 14'b00110100110100;
SIGNAL_B = 14'b10110100001111;
#100;
SIGNAL_A = 14'b00110010100000;
SIGNAL_B = 14'b10110010010010;
#100;
SIGNAL_A = 14'b00110000001001;
SIGNAL_B = 14'b10110000011010;
#100;
SIGNAL_A = 14'b00101101101111;
SIGNAL_B = 14'b10101110101001;
#100;
SIGNAL_A = 14'b00101011010001;
SIGNAL_B = 14'b10101100111111;
#100;
SIGNAL_A = 14'b00101000110000;
SIGNAL_B = 14'b10101011011010;
#100;
SIGNAL_A = 14'b00100110001100;
SIGNAL_B = 14'b10101001111100;
#100;
SIGNAL_A = 14'b00100011100101;
SIGNAL_B = 14'b10101000100100;
#100;
SIGNAL_A = 14'b00100000111100;
SIGNAL_B = 14'b10100111010011;
#100;
SIGNAL_A = 14'b00011110010001;
SIGNAL_B = 14'b10100110001000;
#100;
SIGNAL_A = 14'b00011011100011;
SIGNAL_B = 14'b10100101000011;
#100;
SIGNAL_A = 14'b00011000110100;
SIGNAL_B = 14'b10100100000101;
#100;
SIGNAL_A = 14'b00010110000010;
SIGNAL_B = 14'b10100011001101;
#100;
SIGNAL_A = 14'b00010011001111;
SIGNAL_B = 14'b10100010011011;
#100;
SIGNAL_A = 14'b00010000011011;
SIGNAL_B = 14'b10100001110000;
#100;
SIGNAL_A = 14'b00001101100101;
SIGNAL_B = 14'b10100001001100;
#100;
SIGNAL_A = 14'b00001010101111;
SIGNAL_B = 14'b10100000101101;
#100;
SIGNAL_A = 14'b00000111111000;
SIGNAL_B = 14'b10100000010101;
#100;
SIGNAL_A = 14'b00000101000000;
SIGNAL_B = 14'b10100000000100;
#100;
SIGNAL_A = 14'b00000010000111;
SIGNAL_B = 14'b10011111111000;
#100;
SIGNAL_A = 14'b11111111001111;
SIGNAL_B = 14'b10011111110011;
#100;
SIGNAL_A = 14'b11111100010111;
SIGNAL_B = 14'b10011111110011;
#100;
SIGNAL_A = 14'b11111001011110;
SIGNAL_B = 14'b10011111111010;
#100;
SIGNAL_A = 14'b11110110100110;
SIGNAL_B = 14'b10100000000111;
#100;
SIGNAL_A = 14'b11110011101110;
SIGNAL_B = 14'b10100000011010;
#100;
SIGNAL_A = 14'b11110000110111;
SIGNAL_B = 14'b10100000110010;
#100;
SIGNAL_A = 14'b11101110000000;
SIGNAL_B = 14'b10100001010001;
#100;
SIGNAL_A = 14'b11101011001011;
SIGNAL_B = 14'b10100001110101;
#100;
SIGNAL_A = 14'b11101000010111;
SIGNAL_B = 14'b10100010011110;
#100;
SIGNAL_A = 14'b11100101100100;
SIGNAL_B = 14'b10100011001101;
#100;
SIGNAL_A = 14'b11100010110010;
SIGNAL_B = 14'b10100100000010;
#100;
SIGNAL_A = 14'b11100000000011;
SIGNAL_B = 14'b10100100111100;
#100;
SIGNAL_A = 14'b11011101010101;
SIGNAL_B = 14'b10100101111010;
#100;
SIGNAL_A = 14'b11011010101001;
SIGNAL_B = 14'b10100110111110;
#100;
SIGNAL_A = 14'b11010111111111;
SIGNAL_B = 14'b10101000000111;
#100;
SIGNAL_A = 14'b11010101010111;
SIGNAL_B = 14'b10101001010101;
#100;
SIGNAL_A = 14'b11010010110010;
SIGNAL_B = 14'b10101010101000;
#100;
SIGNAL_A = 14'b11010000001111;
SIGNAL_B = 14'b10101011111111;
#100;
SIGNAL_A = 14'b11001101101111;
SIGNAL_B = 14'b10101101011010;
#100;
SIGNAL_A = 14'b11001011010010;
SIGNAL_B = 14'b10101110111010;
#100;
SIGNAL_A = 14'b11001000111000;
SIGNAL_B = 14'b10110000011110;
#100;
SIGNAL_A = 14'b11000110100001;
SIGNAL_B = 14'b10110010000110;
#100;
SIGNAL_A = 14'b11000100001101;
SIGNAL_B = 14'b10110011110010;
#100;
SIGNAL_A = 14'b11000001111100;
SIGNAL_B = 14'b10110101100001;
#100;
SIGNAL_A = 14'b10111111101111;
SIGNAL_B = 14'b10110111010100;
#100;
SIGNAL_A = 14'b10111101100101;
SIGNAL_B = 14'b10111001001011;
#100;
SIGNAL_A = 14'b10111011011111;
SIGNAL_B = 14'b10111011000101;
#100;
SIGNAL_A = 14'b10111001011100;
SIGNAL_B = 14'b10111101000010;
#100;
SIGNAL_A = 14'b10110111011110;
SIGNAL_B = 14'b10111111000010;
#100;
SIGNAL_A = 14'b10110101100011;
SIGNAL_B = 14'b11000001000101;
#100;
SIGNAL_A = 14'b10110011101100;
SIGNAL_B = 14'b11000011001011;
#100;
SIGNAL_A = 14'b10110001111001;
SIGNAL_B = 14'b11000101010011;
#100;
SIGNAL_A = 14'b10110000001011;
SIGNAL_B = 14'b11000111011101;
#100;
SIGNAL_A = 14'b10101110100000;
SIGNAL_B = 14'b11001001101010;
#100;
SIGNAL_A = 14'b10101101111010;
SIGNAL_B = 14'b11001010101011;
#100;
SIGNAL_A = 14'b10101100011000;
SIGNAL_B = 14'b11001110111011;
#100;
SIGNAL_A = 14'b10101010111101;
SIGNAL_B = 14'b11010011001100;
#100;
SIGNAL_A = 14'b10101001101011;
SIGNAL_B = 14'b11010111011101;
#100;
SIGNAL_A = 14'b10101000100010;
SIGNAL_B = 14'b11011011101110;
#100;
SIGNAL_A = 14'b10100111100000;
SIGNAL_B = 14'b11011111111110;
#100;
SIGNAL_A = 14'b10100110100111;
SIGNAL_B = 14'b11100100001110;
#100;
SIGNAL_A = 14'b10100101110101;
SIGNAL_B = 14'b11101000011101;
#100;
SIGNAL_A = 14'b10100101001100;
SIGNAL_B = 14'b11101100101010;
#100;
SIGNAL_A = 14'b10100100101011;
SIGNAL_B = 14'b11110000110110;
#100;
SIGNAL_A = 14'b10100100010010;
SIGNAL_B = 14'b11110101000001;
#100;
SIGNAL_A = 14'b10100100000001;
SIGNAL_B = 14'b11111001001001;
#100;
SIGNAL_A = 14'b10100011111000;
SIGNAL_B = 14'b11111101010000;
#100;
SIGNAL_A = 14'b10100011110110;
SIGNAL_B = 14'b00000001010011;
#100;
SIGNAL_A = 14'b10100011111100;
SIGNAL_B = 14'b00000101010100;
#100;
SIGNAL_A = 14'b10100100001011;
SIGNAL_B = 14'b00001001010011;
#100;
SIGNAL_A = 14'b10100100100000;
SIGNAL_B = 14'b00001101001110;
#100;
SIGNAL_A = 14'b10100100111101;
SIGNAL_B = 14'b00010001000110;
#100;
SIGNAL_A = 14'b10100101100010;
SIGNAL_B = 14'b00010100111011;
#100;
SIGNAL_A = 14'b10100110001110;
SIGNAL_B = 14'b00011000101100;
#100;
SIGNAL_A = 14'b10100111000001;
SIGNAL_B = 14'b00011100011001;
#100;
SIGNAL_A = 14'b10100111111011;
SIGNAL_B = 14'b00100000000001;
#100;
SIGNAL_A = 14'b10101000111100;
SIGNAL_B = 14'b00100011100110;
#100;
SIGNAL_A = 14'b10101010000011;
SIGNAL_B = 14'b00100111000110;
#100;
SIGNAL_A = 14'b10101011010010;
SIGNAL_B = 14'b00101010100001;
#100;
SIGNAL_A = 14'b10101100100110;
SIGNAL_B = 14'b00101101110111;
#100;
SIGNAL_A = 14'b10101110000010;
SIGNAL_B = 14'b00110001001001;
#100;
SIGNAL_A = 14'b10101111100011;
SIGNAL_B = 14'b00110100010101;
#100;
SIGNAL_A = 14'b10110001001011;
SIGNAL_B = 14'b00110111011100;
#100;
SIGNAL_A = 14'b10110010111000;
SIGNAL_B = 14'b00111010011110;
#100;
SIGNAL_A = 14'b10110100101011;
SIGNAL_B = 14'b00111101011010;
#100;
SIGNAL_A = 14'b10110110100100;
SIGNAL_B = 14'b01000000010000;
#100;
SIGNAL_A = 14'b10111000100010;
SIGNAL_B = 14'b01000011000000;
#100;
SIGNAL_A = 14'b10111010100101;
SIGNAL_B = 14'b01000101101011;
#100;
SIGNAL_A = 14'b10111100101101;
SIGNAL_B = 14'b01001000001111;
#100;
SIGNAL_A = 14'b10111110111010;
SIGNAL_B = 14'b01001010101101;
#100;
SIGNAL_A = 14'b11000001001100;
SIGNAL_B = 14'b01001101000101;
#100;
SIGNAL_A = 14'b11000011100010;
SIGNAL_B = 14'b01001111010110;
#100;
SIGNAL_A = 14'b11000101111101;
SIGNAL_B = 14'b01010001100010;
#100;
SIGNAL_A = 14'b11001000011011;
SIGNAL_B = 14'b01010011100110;
#100;
SIGNAL_A = 14'b11001010111110;
SIGNAL_B = 14'b01010101100100;
#100;
SIGNAL_A = 14'b11001101100100;
SIGNAL_B = 14'b01010111011100;
#100;
SIGNAL_A = 14'b11010000001101;
SIGNAL_B = 14'b01011001001100;
#100;
SIGNAL_A = 14'b11010010111010;
SIGNAL_B = 14'b01011010110110;
#100;
SIGNAL_A = 14'b11010101101010;
SIGNAL_B = 14'b01011100011001;
#100;
SIGNAL_A = 14'b11011000011101;
SIGNAL_B = 14'b01011101110110;
#100;
SIGNAL_A = 14'b11011011010011;
SIGNAL_B = 14'b01011111001011;
#100;
SIGNAL_A = 14'b11011110001011;
SIGNAL_B = 14'b01100000011010;
#100;
SIGNAL_A = 14'b11100001000101;
SIGNAL_B = 14'b01100001100010;
#100;
SIGNAL_A = 14'b11100100000001;
SIGNAL_B = 14'b01100010100011;
#100;
SIGNAL_A = 14'b11100110111111;
SIGNAL_B = 14'b01100011011101;
#100;
SIGNAL_A = 14'b11101001111111;
SIGNAL_B = 14'b01100100010000;
#100;
SIGNAL_A = 14'b11101101000000;
SIGNAL_B = 14'b01100100111101;
#100;
SIGNAL_A = 14'b11110000000010;
SIGNAL_B = 14'b01100101100010;
#100;
SIGNAL_A = 14'b11110011000110;
SIGNAL_B = 14'b01100110000001;
#100;
SIGNAL_A = 14'b11110110001010;
SIGNAL_B = 14'b01100110011001;
#100;
SIGNAL_A = 14'b11111001001111;
SIGNAL_B = 14'b01100110101011;
#100;
SIGNAL_A = 14'b11111100010100;
SIGNAL_B = 14'b01100110110110;
#100;
SIGNAL_A = 14'b11111111011010;
SIGNAL_B = 14'b01100110111010;
#100;
SIGNAL_A = 14'b00000010011110;
SIGNAL_B = 14'b01100110110111;
#100;
SIGNAL_A = 14'b00000101100100;
SIGNAL_B = 14'b01100110101111;
#100;
SIGNAL_A = 14'b00001000101001;
SIGNAL_B = 14'b01100110100000;
#100;
SIGNAL_A = 14'b00001011101101;
SIGNAL_B = 14'b01100110001010;
#100;
SIGNAL_A = 14'b00001110110001;
SIGNAL_B = 14'b01100101101110;
#100;
SIGNAL_A = 14'b00010001110100;
SIGNAL_B = 14'b01100101001100;
#100;
SIGNAL_A = 14'b00010100110110;
SIGNAL_B = 14'b01100100100101;
#100;
SIGNAL_A = 14'b00010111110110;
SIGNAL_B = 14'b01100011110111;
#100;
SIGNAL_A = 14'b00011010110101;
SIGNAL_B = 14'b01100011000011;
#100;
SIGNAL_A = 14'b00011101110011;
SIGNAL_B = 14'b01100010001010;
#100;
SIGNAL_A = 14'b00100000101110;
SIGNAL_B = 14'b01100001001011;
#100;
SIGNAL_A = 14'b00100011101000;
SIGNAL_B = 14'b01100000000110;
#100;
SIGNAL_A = 14'b00100110011111;
SIGNAL_B = 14'b01011110111100;
#100;
SIGNAL_A = 14'b00101001010100;
SIGNAL_B = 14'b01011101101101;
#100;
SIGNAL_A = 14'b00101100000111;
SIGNAL_B = 14'b01011100011001;
#100;
SIGNAL_A = 14'b00101110110111;
SIGNAL_B = 14'b01011010111111;
#100;
SIGNAL_A = 14'b00110001100100;
SIGNAL_B = 14'b01011001100001;
#100;
SIGNAL_A = 14'b00110100001111;
SIGNAL_B = 14'b01010111111110;
#100;
SIGNAL_A = 14'b00110110110110;
SIGNAL_B = 14'b01010110010111;
#100;
SIGNAL_A = 14'b00111001011010;
SIGNAL_B = 14'b01010100101011;
#100;
SIGNAL_A = 14'b00111011111011;
SIGNAL_B = 14'b01010010111011;
#100;
SIGNAL_A = 14'b00111110011001;
SIGNAL_B = 14'b01010001000110;
#100;
SIGNAL_A = 14'b01000000110011;
SIGNAL_B = 14'b01001111001110;
#100;
SIGNAL_A = 14'b01000011001001;
SIGNAL_B = 14'b01001101010010;
#100;
SIGNAL_A = 14'b01000101011011;
SIGNAL_B = 14'b01001011010010;
#100;
SIGNAL_A = 14'b01000111101010;
SIGNAL_B = 14'b01001001001111;
#100;
SIGNAL_A = 14'b01001001110100;
SIGNAL_B = 14'b01000111001001;
#100;
SIGNAL_A = 14'b01001011111011;
SIGNAL_B = 14'b01000100111111;
#100;
SIGNAL_A = 14'b01001101111101;
SIGNAL_B = 14'b01000010110010;
#100;
SIGNAL_A = 14'b01001111111011;
SIGNAL_B = 14'b01000000100011;
#100;
SIGNAL_A = 14'b01010001110101;
SIGNAL_B = 14'b00111110010001;
#100;
SIGNAL_A = 14'b01010011101011;
SIGNAL_B = 14'b00111011111100;
#100;
SIGNAL_A = 14'b01010101011011;
SIGNAL_B = 14'b00111001100101;
#100;
SIGNAL_A = 14'b01010110011101;
SIGNAL_B = 14'b00110111000000;
#100;
SIGNAL_A = 14'b01011000000010;
SIGNAL_B = 14'b00110010100101;
#100;
SIGNAL_A = 14'b01011001011111;
SIGNAL_B = 14'b00101110001010;
#100;
SIGNAL_A = 14'b01011010110100;
SIGNAL_B = 14'b00101001101111;
#100;
SIGNAL_A = 14'b01011100000000;
SIGNAL_B = 14'b00100101010100;
#100;
SIGNAL_A = 14'b01011101000011;
SIGNAL_B = 14'b00100000111001;
#100;
SIGNAL_A = 14'b01011101111110;
SIGNAL_B = 14'b00011100011111;
#100;
SIGNAL_A = 14'b01011110110000;
SIGNAL_B = 14'b00011000000110;
#100;
SIGNAL_A = 14'b01011111011010;
SIGNAL_B = 14'b00010011101111;
#100;
SIGNAL_A = 14'b01011111111100;
SIGNAL_B = 14'b00001111011001;
#100;
SIGNAL_A = 14'b01100000010110;
SIGNAL_B = 14'b00001011000100;
#100;
SIGNAL_A = 14'b01100000100111;
SIGNAL_B = 14'b00000110110010;
#100;
SIGNAL_A = 14'b01100000110000;
SIGNAL_B = 14'b00000010100010;
#100;
SIGNAL_A = 14'b01100000110001;
SIGNAL_B = 14'b11111110010101;
#100;
SIGNAL_A = 14'b01100000101001;
SIGNAL_B = 14'b11111010001011;
#100;
SIGNAL_A = 14'b01100000011010;
SIGNAL_B = 14'b11110110000011;
#100;
SIGNAL_A = 14'b01100000000011;
SIGNAL_B = 14'b11110001111110;
#100;
SIGNAL_A = 14'b01011111100100;
SIGNAL_B = 14'b11101101111101;
#100;
SIGNAL_A = 14'b01011110111110;
SIGNAL_B = 14'b11101010000000;
#100;
SIGNAL_A = 14'b01011110010000;
SIGNAL_B = 14'b11100110000110;
#100;
SIGNAL_A = 14'b01011101011010;
SIGNAL_B = 14'b11100010010001;
#100;
SIGNAL_A = 14'b01011100011110;
SIGNAL_B = 14'b11011110011111;
#100;
SIGNAL_A = 14'b01011011011010;
SIGNAL_B = 14'b11011010110011;
#100;
SIGNAL_A = 14'b01011010001111;
SIGNAL_B = 14'b11010111001011;
#100;
SIGNAL_A = 14'b01011000111101;
SIGNAL_B = 14'b11010011101000;
#100;
SIGNAL_A = 14'b01010111100100;
SIGNAL_B = 14'b11010000001010;
#100;
SIGNAL_A = 14'b01010110000101;
SIGNAL_B = 14'b11001100110001;
#100;
SIGNAL_A = 14'b01010100100000;
SIGNAL_B = 14'b11001001011101;
#100;
SIGNAL_A = 14'b01010010110100;
SIGNAL_B = 14'b11000110001111;
#100;
SIGNAL_A = 14'b01010001000010;
SIGNAL_B = 14'b11000011000111;
#100;
SIGNAL_A = 14'b01001111001010;
SIGNAL_B = 14'b11000000000100;
#100;
SIGNAL_A = 14'b01001101001100;
SIGNAL_B = 14'b10111101001000;
#100;
SIGNAL_A = 14'b01001011001001;
SIGNAL_B = 14'b10111010010001;
#100;
SIGNAL_A = 14'b01001001000001;
SIGNAL_B = 14'b10110111100001;
#100;
SIGNAL_A = 14'b01000110110011;
SIGNAL_B = 14'b10110100110111;
#100;
SIGNAL_A = 14'b01000100100000;
SIGNAL_B = 14'b10110010010011;
#100;
SIGNAL_A = 14'b01000010001000;
SIGNAL_B = 14'b10101111110110;
#100;
SIGNAL_A = 14'b00111111101100;
SIGNAL_B = 14'b10101101100000;
#100;
SIGNAL_A = 14'b00111101001100;
SIGNAL_B = 14'b10101011010000;
#100;
SIGNAL_A = 14'b00111010100111;
SIGNAL_B = 14'b10101001000111;
#100;
SIGNAL_A = 14'b00110111111110;
SIGNAL_B = 14'b10100111000101;
#100;
SIGNAL_A = 14'b00110101010001;
SIGNAL_B = 14'b10100101001001;
#100;
SIGNAL_A = 14'b00110010100001;
SIGNAL_B = 14'b10100011010101;
#100;
SIGNAL_A = 14'b00101111101110;
SIGNAL_B = 14'b10100001101000;
#100;
SIGNAL_A = 14'b00101100110111;
SIGNAL_B = 14'b10100000000001;
#100;
SIGNAL_A = 14'b00101001111101;
SIGNAL_B = 14'b10011110100010;
#100;
SIGNAL_A = 14'b00100111000001;
SIGNAL_B = 14'b10011101001010;
#100;
SIGNAL_A = 14'b00100100000010;
SIGNAL_B = 14'b10011011111001;
#100;
SIGNAL_A = 14'b00100001000000;
SIGNAL_B = 14'b10011010101111;
#100;
SIGNAL_A = 14'b00011101111101;
SIGNAL_B = 14'b10011001101100;
#100;
SIGNAL_A = 14'b00011010110111;
SIGNAL_B = 14'b10011000110000;
#100;
SIGNAL_A = 14'b00010111110000;
SIGNAL_B = 14'b10010111111011;
#100;
SIGNAL_A = 14'b00010100101000;
SIGNAL_B = 14'b10010111001110;
#100;
SIGNAL_A = 14'b00010001011110;
SIGNAL_B = 14'b10010110100111;
#100;
SIGNAL_A = 14'b00001110010011;
SIGNAL_B = 14'b10010110001000;
#100;
SIGNAL_A = 14'b00001011000111;
SIGNAL_B = 14'b10010101101111;
#100;
SIGNAL_A = 14'b00000111111011;
SIGNAL_B = 14'b10010101011110;
#100;
SIGNAL_A = 14'b00000100101110;
SIGNAL_B = 14'b10010101010011;
#100;
SIGNAL_A = 14'b00000001100001;
SIGNAL_B = 14'b10010101001111;
#100;
SIGNAL_A = 14'b11111110010101;
SIGNAL_B = 14'b10010101010010;
#100;
SIGNAL_A = 14'b11111011001001;
SIGNAL_B = 14'b10010101011100;
#100;
SIGNAL_A = 14'b11110111111100;
SIGNAL_B = 14'b10010101101100;
#100;
SIGNAL_A = 14'b11110100110000;
SIGNAL_B = 14'b10010110000011;
#100;
SIGNAL_A = 14'b11110001100101;
SIGNAL_B = 14'b10010110100000;
#100;
SIGNAL_A = 14'b11101110011011;
SIGNAL_B = 14'b10010111000100;
#100;
SIGNAL_A = 14'b11101011010011;
SIGNAL_B = 14'b10010111101110;
#100;
SIGNAL_A = 14'b11101000001011;
SIGNAL_B = 14'b10011000011110;
#100;
SIGNAL_A = 14'b11100101000101;
SIGNAL_B = 14'b10011001010100;
#100;
SIGNAL_A = 14'b11100010000001;
SIGNAL_B = 14'b10011010010000;
#100;
SIGNAL_A = 14'b11011110111110;
SIGNAL_B = 14'b10011011010010;
#100;
SIGNAL_A = 14'b11011011111110;
SIGNAL_B = 14'b10011100011001;
#100;
SIGNAL_A = 14'b11011001000000;
SIGNAL_B = 14'b10011101100110;
#100;
SIGNAL_A = 14'b11010110000100;
SIGNAL_B = 14'b10011110111001;
#100;
SIGNAL_A = 14'b11010011001011;
SIGNAL_B = 14'b10100000010001;
#100;
SIGNAL_A = 14'b11010000010100;
SIGNAL_B = 14'b10100001101110;
#100;
SIGNAL_A = 14'b11001101100001;
SIGNAL_B = 14'b10100011010000;
#100;
SIGNAL_A = 14'b11001010110000;
SIGNAL_B = 14'b10100100110111;
#100;
SIGNAL_A = 14'b11001000000011;
SIGNAL_B = 14'b10100110100011;
#100;
SIGNAL_A = 14'b11000101011001;
SIGNAL_B = 14'b10101000010011;
#100;
SIGNAL_A = 14'b11000010110010;
SIGNAL_B = 14'b10101010001000;
#100;
SIGNAL_A = 14'b11000000001111;
SIGNAL_B = 14'b10101100000000;
#100;
SIGNAL_A = 14'b10111101110000;
SIGNAL_B = 14'b10101101111110;
#100;
SIGNAL_A = 14'b10111011010100;
SIGNAL_B = 14'b10101111111111;
#100;
SIGNAL_A = 14'b10111000111100;
SIGNAL_B = 14'b10110010000011;
#100;
SIGNAL_A = 14'b10110110101001;
SIGNAL_B = 14'b10110100001100;
#100;
SIGNAL_A = 14'b10110100011001;
SIGNAL_B = 14'b10110110011000;
#100;
SIGNAL_A = 14'b10110010001110;
SIGNAL_B = 14'b10111000100111;
#100;
SIGNAL_A = 14'b10110000000111;
SIGNAL_B = 14'b10111010111001;
#100;
SIGNAL_A = 14'b10101110000101;
SIGNAL_B = 14'b10111101001110;
#100;
SIGNAL_A = 14'b10101100000111;
SIGNAL_B = 14'b10111111100110;
#100;
SIGNAL_A = 14'b10101010001101;
SIGNAL_B = 14'b11000010000000;
#100;
SIGNAL_A = 14'b10101000100000;
SIGNAL_B = 14'b11000100010011;
#100;
SIGNAL_A = 14'b10100111101111;
SIGNAL_B = 14'b11000110001011;
#100;
SIGNAL_A = 14'b10100110000100;
SIGNAL_B = 14'b11001010101011;
#100;
SIGNAL_A = 14'b10100100100010;
SIGNAL_B = 14'b11001111001100;
#100;
SIGNAL_A = 14'b10100011001001;
SIGNAL_B = 14'b11010011101101;
#100;
SIGNAL_A = 14'b10100001111000;
SIGNAL_B = 14'b11011000001110;
#100;
SIGNAL_A = 14'b10100000110000;
SIGNAL_B = 14'b11011100101111;
#100;
SIGNAL_A = 14'b10011111110001;
SIGNAL_B = 14'b11100001001111;
#100;
SIGNAL_A = 14'b10011110111010;
SIGNAL_B = 14'b11100101101110;
#100;
SIGNAL_A = 14'b10011110001100;
SIGNAL_B = 14'b11101010001100;
#100;
SIGNAL_A = 14'b10011101100110;
SIGNAL_B = 14'b11101110101000;
#100;
SIGNAL_A = 14'b10011101001001;
SIGNAL_B = 14'b11110011000011;
#100;
SIGNAL_A = 14'b10011100110100;
SIGNAL_B = 14'b11110111011100;
#100;
SIGNAL_A = 14'b10011100101000;
SIGNAL_B = 14'b11111011110011;
#100;
SIGNAL_A = 14'b10011100100100;
SIGNAL_B = 14'b00000000000110;
#100;
SIGNAL_A = 14'b10011100101001;
SIGNAL_B = 14'b00000100010111;
#100;
SIGNAL_A = 14'b10011100110101;
SIGNAL_B = 14'b00001000100110;
#100;
SIGNAL_A = 14'b10011101001010;
SIGNAL_B = 14'b00001100110001;
#100;
SIGNAL_A = 14'b10011101100110;
SIGNAL_B = 14'b00010000111001;
#100;
SIGNAL_A = 14'b10011110001010;
SIGNAL_B = 14'b00010100111101;
#100;
SIGNAL_A = 14'b10011110110110;
SIGNAL_B = 14'b00011000111110;
#100;
SIGNAL_A = 14'b10011111101010;
SIGNAL_B = 14'b00011100111010;
#100;
SIGNAL_A = 14'b10100000100101;
SIGNAL_B = 14'b00100000110010;
#100;
SIGNAL_A = 14'b10100001101000;
SIGNAL_B = 14'b00100100100101;
#100;
SIGNAL_A = 14'b10100010110010;
SIGNAL_B = 14'b00101000010100;
#100;
SIGNAL_A = 14'b10100100000011;
SIGNAL_B = 14'b00101011111101;
#100;
SIGNAL_A = 14'b10100101011011;
SIGNAL_B = 14'b00101111100010;
#100;
SIGNAL_A = 14'b10100110111001;
SIGNAL_B = 14'b00110011000010;
#100;
SIGNAL_A = 14'b10101000011111;
SIGNAL_B = 14'b00110110011100;
#100;
SIGNAL_A = 14'b10101010001010;
SIGNAL_B = 14'b00111001110000;
#100;
SIGNAL_A = 14'b10101011111100;
SIGNAL_B = 14'b00111100111111;
#100;
SIGNAL_A = 14'b10101101110100;
SIGNAL_B = 14'b01000000001000;
#100;
SIGNAL_A = 14'b10101111110011;
SIGNAL_B = 14'b01000011001010;
#100;
SIGNAL_A = 14'b10110001110110;
SIGNAL_B = 14'b01000110000111;
#100;
SIGNAL_A = 14'b10110100000000;
SIGNAL_B = 14'b01001000111101;
#100;
SIGNAL_A = 14'b10110110001110;
SIGNAL_B = 14'b01001011101101;
#100;
SIGNAL_A = 14'b10111000100010;
SIGNAL_B = 14'b01001110010111;
#100;
SIGNAL_A = 14'b10111010111011;
SIGNAL_B = 14'b01010000111010;
#100;
SIGNAL_A = 14'b10111101011001;
SIGNAL_B = 14'b01010011010110;
#100;
SIGNAL_A = 14'b10111111111011;
SIGNAL_B = 14'b01010101101011;
#100;
SIGNAL_A = 14'b11000010100010;
SIGNAL_B = 14'b01010111111010;
#100;
SIGNAL_A = 14'b11000101001101;
SIGNAL_B = 14'b01011010000001;
#100;
SIGNAL_A = 14'b11000111111100;
SIGNAL_B = 14'b01011100000010;
#100;
SIGNAL_A = 14'b11001010101110;
SIGNAL_B = 14'b01011101111011;
#100;
SIGNAL_A = 14'b11001101100100;
SIGNAL_B = 14'b01011111101110;
#100;
SIGNAL_A = 14'b11010000011110;
SIGNAL_B = 14'b01100001011001;
#100;
SIGNAL_A = 14'b11010011011010;
SIGNAL_B = 14'b01100010111101;
#100;
SIGNAL_A = 14'b11010110011010;
SIGNAL_B = 14'b01100100011010;
#100;
SIGNAL_A = 14'b11011001011100;
SIGNAL_B = 14'b01100101101111;
#100;
SIGNAL_A = 14'b11011100100000;
SIGNAL_B = 14'b01100110111101;
#100;
SIGNAL_A = 14'b11011111100111;
SIGNAL_B = 14'b01101000000100;
#100;
SIGNAL_A = 14'b11100010110000;
SIGNAL_B = 14'b01101001000100;
#100;
SIGNAL_A = 14'b11100101111010;
SIGNAL_B = 14'b01101001111101;
#100;
SIGNAL_A = 14'b11101001000111;
SIGNAL_B = 14'b01101010101110;
#100;
SIGNAL_A = 14'b11101100010100;
SIGNAL_B = 14'b01101011011000;
#100;
SIGNAL_A = 14'b11101111100011;
SIGNAL_B = 14'b01101011111011;
#100;
SIGNAL_A = 14'b11110010110010;
SIGNAL_B = 14'b01101100010110;
#100;
SIGNAL_A = 14'b11110110000011;
SIGNAL_B = 14'b01101100101011;
#100;
SIGNAL_A = 14'b11111001010100;
SIGNAL_B = 14'b01101100111000;
#100;
SIGNAL_A = 14'b11111100100101;
SIGNAL_B = 14'b01101100111111;
#100;
SIGNAL_A = 14'b11111111110110;
SIGNAL_B = 14'b01101100111111;
#100;
SIGNAL_A = 14'b00000011000110;
SIGNAL_B = 14'b01101100110111;
#100;
SIGNAL_A = 14'b00000110010111;
SIGNAL_B = 14'b01101100101001;
#100;
SIGNAL_A = 14'b00001001101000;
SIGNAL_B = 14'b01101100010101;
#100;
SIGNAL_A = 14'b00001100110111;
SIGNAL_B = 14'b01101011111001;
#100;
SIGNAL_A = 14'b00010000000110;
SIGNAL_B = 14'b01101011010111;
#100;
SIGNAL_A = 14'b00010011010011;
SIGNAL_B = 14'b01101010101111;
#100;
SIGNAL_A = 14'b00010110100000;
SIGNAL_B = 14'b01101010000000;
#100;
SIGNAL_A = 14'b00011001101010;
SIGNAL_B = 14'b01101001001011;
#100;
SIGNAL_A = 14'b00011100110011;
SIGNAL_B = 14'b01101000010000;
#100;
SIGNAL_A = 14'b00011111111011;
SIGNAL_B = 14'b01100111001111;
#100;
SIGNAL_A = 14'b00100011000000;
SIGNAL_B = 14'b01100110001000;
#100;
SIGNAL_A = 14'b00100110000011;
SIGNAL_B = 14'b01100100111100;
#100;
SIGNAL_A = 14'b00101001000011;
SIGNAL_B = 14'b01100011101001;
#100;
SIGNAL_A = 14'b00101100000001;
SIGNAL_B = 14'b01100010010010;
#100;
SIGNAL_A = 14'b00101110111101;
SIGNAL_B = 14'b01100000110101;
#100;
SIGNAL_A = 14'b00110001110101;
SIGNAL_B = 14'b01011111010010;
#100;
SIGNAL_A = 14'b00110100101011;
SIGNAL_B = 14'b01011101101011;
#100;
SIGNAL_A = 14'b00110111011101;
SIGNAL_B = 14'b01011011111111;
#100;
SIGNAL_A = 14'b00111010001100;
SIGNAL_B = 14'b01011010001110;
#100;
SIGNAL_A = 14'b00111100110111;
SIGNAL_B = 14'b01011000011001;
#100;
SIGNAL_A = 14'b00111111011111;
SIGNAL_B = 14'b01010110011111;
#100;
SIGNAL_A = 14'b01000010000011;
SIGNAL_B = 14'b01010100100001;
#100;
SIGNAL_A = 14'b01000100100100;
SIGNAL_B = 14'b01010010011110;
#100;
SIGNAL_A = 14'b01000111000000;
SIGNAL_B = 14'b01010000011000;
#100;
SIGNAL_A = 14'b01001001011000;
SIGNAL_B = 14'b01001110001110;
#100;
SIGNAL_A = 14'b01001011101100;
SIGNAL_B = 14'b01001100000001;
#100;
SIGNAL_A = 14'b01001101111100;
SIGNAL_B = 14'b01001001110000;
#100;
SIGNAL_A = 14'b01010000001000;
SIGNAL_B = 14'b01000111011100;
#100;
SIGNAL_A = 14'b01010010001111;
SIGNAL_B = 14'b01000101000101;
#100;
SIGNAL_A = 14'b01010100010001;
SIGNAL_B = 14'b01000010101011;
#100;
SIGNAL_A = 14'b01010110001111;
SIGNAL_B = 14'b01000000001110;
#100;
SIGNAL_A = 14'b01011000001000;
SIGNAL_B = 14'b00111101101111;
#100;
SIGNAL_A = 14'b01011001001110;
SIGNAL_B = 14'b00111011101011;
#100;
SIGNAL_A = 14'b01011010111101;
SIGNAL_B = 14'b00110111001000;
#100;
SIGNAL_A = 14'b01011100100010;
SIGNAL_B = 14'b00110010100100;
#100;
SIGNAL_A = 14'b01011101111111;
SIGNAL_B = 14'b00101101111111;
#100;
SIGNAL_A = 14'b01011111010011;
SIGNAL_B = 14'b00101001011011;
#100;
SIGNAL_A = 14'b01100000011110;
SIGNAL_B = 14'b00100100110110;
#100;
SIGNAL_A = 14'b01100001100000;
SIGNAL_B = 14'b00100000010011;
#100;
SIGNAL_A = 14'b01100010011010;
SIGNAL_B = 14'b00011011110000;
#100;
SIGNAL_A = 14'b01100011001011;
SIGNAL_B = 14'b00010111001110;
#100;
SIGNAL_A = 14'b01100011110011;
SIGNAL_B = 14'b00010010101110;
#100;
SIGNAL_A = 14'b01100100010011;
SIGNAL_B = 14'b00001110001111;
#100;
SIGNAL_A = 14'b01100100101010;
SIGNAL_B = 14'b00001001110010;
#100;
SIGNAL_A = 14'b01100100111000;
SIGNAL_B = 14'b00000101011000;
#100;
SIGNAL_A = 14'b01100100111111;
SIGNAL_B = 14'b00000001000000;
#100;
SIGNAL_A = 14'b01100100111100;
SIGNAL_B = 14'b11111100101011;
#100;
SIGNAL_A = 14'b01100100110010;
SIGNAL_B = 14'b11111000011001;
#100;
SIGNAL_A = 14'b01100100011111;
SIGNAL_B = 14'b11110100001001;
#100;
SIGNAL_A = 14'b01100100000100;
SIGNAL_B = 14'b11101111111110;
#100;
SIGNAL_A = 14'b01100011100010;
SIGNAL_B = 14'b11101011110101;
#100;
SIGNAL_A = 14'b01100010110111;
SIGNAL_B = 14'b11100111110001;
#100;
SIGNAL_A = 14'b01100010000100;
SIGNAL_B = 14'b11100011110001;
#100;
SIGNAL_A = 14'b01100001001010;
SIGNAL_B = 14'b11011111110101;
#100;
SIGNAL_A = 14'b01100000001001;
SIGNAL_B = 14'b11011011111101;
#100;
SIGNAL_A = 14'b01011111000000;
SIGNAL_B = 14'b11011000001011;
#100;
SIGNAL_A = 14'b01011101110000;
SIGNAL_B = 14'b11010100011101;
#100;
SIGNAL_A = 14'b01011100011001;
SIGNAL_B = 14'b11010000110100;
#100;
SIGNAL_A = 14'b01011010111011;
SIGNAL_B = 14'b11001101010001;
#100;
SIGNAL_A = 14'b01011001010110;
SIGNAL_B = 14'b11001001110011;
#100;
SIGNAL_A = 14'b01010111101011;
SIGNAL_B = 14'b11000110011010;
#100;
SIGNAL_A = 14'b01010101111001;
SIGNAL_B = 14'b11000011000111;
#100;
SIGNAL_A = 14'b01010100000001;
SIGNAL_B = 14'b10111111111011;
#100;
SIGNAL_A = 14'b01010010000011;
SIGNAL_B = 14'b10111100110100;
#100;
SIGNAL_A = 14'b01001111111111;
SIGNAL_B = 14'b10111001110100;
#100;
SIGNAL_A = 14'b01001101110101;
SIGNAL_B = 14'b10110110111001;
#100;
SIGNAL_A = 14'b01001011100110;
SIGNAL_B = 14'b10110100000110;
#100;
SIGNAL_A = 14'b01001001010010;
SIGNAL_B = 14'b10110001011000;
#100;
SIGNAL_A = 14'b01000110111000;
SIGNAL_B = 14'b10101110110010;
#100;
SIGNAL_A = 14'b01000100011010;
SIGNAL_B = 14'b10101100010010;
#100;
SIGNAL_A = 14'b01000001110111;
SIGNAL_B = 14'b10101001111001;
#100;
SIGNAL_A = 14'b00111111001111;
SIGNAL_B = 14'b10100111100111;
#100;
SIGNAL_A = 14'b00111100100100;
SIGNAL_B = 14'b10100101011100;
#100;
SIGNAL_A = 14'b00111001110100;
SIGNAL_B = 14'b10100011011001;
#100;
SIGNAL_A = 14'b00110111000000;
SIGNAL_B = 14'b10100001011100;
#100;
SIGNAL_A = 14'b00110100001001;
SIGNAL_B = 14'b10011111100110;
#100;
SIGNAL_A = 14'b00110001001110;
SIGNAL_B = 14'b10011101111000;
#100;
SIGNAL_A = 14'b00101110010000;
SIGNAL_B = 14'b10011100010001;
#100;
SIGNAL_A = 14'b00101011001111;
SIGNAL_B = 14'b10011010110001;
#100;
SIGNAL_A = 14'b00101000001011;
SIGNAL_B = 14'b10011001011001;
#100;
SIGNAL_A = 14'b00100101000101;
SIGNAL_B = 14'b10011000001000;
#100;
SIGNAL_A = 14'b00100001111100;
SIGNAL_B = 14'b10010110111110;
#100;
SIGNAL_A = 14'b00011110110010;
SIGNAL_B = 14'b10010101111100;
#100;
SIGNAL_A = 14'b00011011100101;
SIGNAL_B = 14'b10010101000001;
#100;
SIGNAL_A = 14'b00011000010111;
SIGNAL_B = 14'b10010100001101;
#100;
SIGNAL_A = 14'b00010101000111;
SIGNAL_B = 14'b10010011100001;
#100;
SIGNAL_A = 14'b00010001110110;
SIGNAL_B = 14'b10010010111100;
#100;
SIGNAL_A = 14'b00001110100100;
SIGNAL_B = 14'b10010010011110;
#100;
SIGNAL_A = 14'b00001011010010;
SIGNAL_B = 14'b10010010000111;
#100;
SIGNAL_A = 14'b00000111111111;
SIGNAL_B = 14'b10010001110111;
#100;
SIGNAL_A = 14'b00000100101011;
SIGNAL_B = 14'b10010001101111;
#100;
SIGNAL_A = 14'b00000001010111;
SIGNAL_B = 14'b10010001101110;
#100;
SIGNAL_A = 14'b11111110000100;
SIGNAL_B = 14'b10010001110011;
#100;
SIGNAL_A = 14'b11111010110001;
SIGNAL_B = 14'b10010010000000;
#100;
SIGNAL_A = 14'b11110111011110;
SIGNAL_B = 14'b10010010010011;
#100;
SIGNAL_A = 14'b11110100001100;
SIGNAL_B = 14'b10010010101101;
#100;
SIGNAL_A = 14'b11110000111010;
SIGNAL_B = 14'b10010011001110;
#100;
SIGNAL_A = 14'b11101101101010;
SIGNAL_B = 14'b10010011110101;
#100;
SIGNAL_A = 14'b11101010011011;
SIGNAL_B = 14'b10010100100011;
#100;
SIGNAL_A = 14'b11100111001101;
SIGNAL_B = 14'b10010101010111;
#100;
SIGNAL_A = 14'b11100100000010;
SIGNAL_B = 14'b10010110010001;
#100;
SIGNAL_A = 14'b11100000110111;
SIGNAL_B = 14'b10010111010001;
#100;
SIGNAL_A = 14'b11011101101111;
SIGNAL_B = 14'b10011000010111;
#100;
SIGNAL_A = 14'b11011010101010;
SIGNAL_B = 14'b10011001100011;
#100;
SIGNAL_A = 14'b11010111100110;
SIGNAL_B = 14'b10011010110101;
#100;
SIGNAL_A = 14'b11010100100101;
SIGNAL_B = 14'b10011100001100;
#100;
SIGNAL_A = 14'b11010001100111;
SIGNAL_B = 14'b10011101101001;
#100;
SIGNAL_A = 14'b11001110101011;
SIGNAL_B = 14'b10011111001011;
#100;
SIGNAL_A = 14'b11001011110011;
SIGNAL_B = 14'b10100000110011;
#100;
SIGNAL_A = 14'b11001000111110;
SIGNAL_B = 14'b10100010011111;
#100;
SIGNAL_A = 14'b11000110001100;
SIGNAL_B = 14'b10100100010000;
#100;
SIGNAL_A = 14'b11000011011101;
SIGNAL_B = 14'b10100110000101;
#100;
SIGNAL_A = 14'b11000000110011;
SIGNAL_B = 14'b10101000000000;
#100;
SIGNAL_A = 14'b10111110001100;
SIGNAL_B = 14'b10101001111110;
#100;
SIGNAL_A = 14'b10111011101000;
SIGNAL_B = 14'b10101100000001;
#100;
SIGNAL_A = 14'b10111001001001;
SIGNAL_B = 14'b10101110001000;
#100;
SIGNAL_A = 14'b10110110101110;
SIGNAL_B = 14'b10110000010010;
#100;
SIGNAL_A = 14'b10110100010111;
SIGNAL_B = 14'b10110010100001;
#100;
SIGNAL_A = 14'b10110010000100;
SIGNAL_B = 14'b10110100110010;
#100;
SIGNAL_A = 14'b10101111110110;
SIGNAL_B = 14'b10110111000111;
#100;
SIGNAL_A = 14'b10101101101100;
SIGNAL_B = 14'b10111001011111;
#100;
SIGNAL_A = 14'b10101011100111;
SIGNAL_B = 14'b10111011111011;
#100;
SIGNAL_A = 14'b10101001100111;
SIGNAL_B = 14'b10111110011000;
#100;
SIGNAL_A = 14'b10100111101011;
SIGNAL_B = 14'b11000000111001;
#100;
SIGNAL_A = 14'b10100110100100;
SIGNAL_B = 14'b11000010011010;
#100;
SIGNAL_A = 14'b10100101000100;
SIGNAL_B = 14'b11000110001111;
#100;
SIGNAL_A = 14'b10100011011001;
SIGNAL_B = 14'b11001010110101;
#100;
SIGNAL_A = 14'b10100001111000;
SIGNAL_B = 14'b11001111011011;
#100;
SIGNAL_A = 14'b10100000011111;
SIGNAL_B = 14'b11010100000010;
#100;
SIGNAL_A = 14'b10011111001111;
SIGNAL_B = 14'b11011000101000;
#100;
SIGNAL_A = 14'b10011110001000;
SIGNAL_B = 14'b11011101001110;
#100;
SIGNAL_A = 14'b10011101001001;
SIGNAL_B = 14'b11100001110100;
#100;
SIGNAL_A = 14'b10011100010100;
SIGNAL_B = 14'b11100110011000;
#100;
SIGNAL_A = 14'b10011011100111;
SIGNAL_B = 14'b11101010111011;
#100;
SIGNAL_A = 14'b10011011000011;
SIGNAL_B = 14'b11101111011100;
#100;
SIGNAL_A = 14'b10011010100111;
SIGNAL_B = 14'b11110011111100;
#100;
SIGNAL_A = 14'b10011010010100;
SIGNAL_B = 14'b11111000011010;
#100;
SIGNAL_A = 14'b10011010001010;
SIGNAL_B = 14'b11111100110101;
#100;
SIGNAL_A = 14'b10011010001000;
SIGNAL_B = 14'b00000001001101;
#100;
SIGNAL_A = 14'b10011010001111;
SIGNAL_B = 14'b00000101100011;
#100;
SIGNAL_A = 14'b10011010011101;
SIGNAL_B = 14'b00001001110101;
#100;
SIGNAL_A = 14'b10011010110100;
SIGNAL_B = 14'b00001110000101;
#100;
SIGNAL_A = 14'b10011011010011;
SIGNAL_B = 14'b00010010010001;
#100;
SIGNAL_A = 14'b10011011111010;
SIGNAL_B = 14'b00010110011001;
#100;
SIGNAL_A = 14'b10011100101001;
SIGNAL_B = 14'b00011010011101;
#100;
SIGNAL_A = 14'b10011101100000;
SIGNAL_B = 14'b00011110011101;
#100;
SIGNAL_A = 14'b10011110011110;
SIGNAL_B = 14'b00100010011000;
#100;
SIGNAL_A = 14'b10011111100100;
SIGNAL_B = 14'b00100110001111;
#100;
SIGNAL_A = 14'b10100000110001;
SIGNAL_B = 14'b00101010000001;
#100;
SIGNAL_A = 14'b10100010000101;
SIGNAL_B = 14'b00101101101110;
#100;
SIGNAL_A = 14'b10100011100001;
SIGNAL_B = 14'b00110001010101;
#100;
SIGNAL_A = 14'b10100101000011;
SIGNAL_B = 14'b00110100111000;
#100;
SIGNAL_A = 14'b10100110101100;
SIGNAL_B = 14'b00111000010100;
#100;
SIGNAL_A = 14'b10101000011011;
SIGNAL_B = 14'b00111011101011;
#100;
SIGNAL_A = 14'b10101010010001;
SIGNAL_B = 14'b00111110111100;
#100;
SIGNAL_A = 14'b10101100001101;
SIGNAL_B = 14'b01000010000111;
#100;
SIGNAL_A = 14'b10101110001111;
SIGNAL_B = 14'b01000101001100;
#100;
SIGNAL_A = 14'b10110000010110;
SIGNAL_B = 14'b01001000001011;
#100;
SIGNAL_A = 14'b10110010100100;
SIGNAL_B = 14'b01001011000011;
#100;
SIGNAL_A = 14'b10110100110110;
SIGNAL_B = 14'b01001101110101;
#100;
SIGNAL_A = 14'b10110111001110;
SIGNAL_B = 14'b01010000100000;
#100;
SIGNAL_A = 14'b10111001101011;
SIGNAL_B = 14'b01010011000100;
#100;
SIGNAL_A = 14'b10111100001101;
SIGNAL_B = 14'b01010101100001;
#100;
SIGNAL_A = 14'b10111110110100;
SIGNAL_B = 14'b01010111111000;
#100;
SIGNAL_A = 14'b11000001011111;
SIGNAL_B = 14'b01011010000111;
#100;
SIGNAL_A = 14'b11000100001110;
SIGNAL_B = 14'b01011100001111;
#100;
SIGNAL_A = 14'b11000111000001;
SIGNAL_B = 14'b01011110010000;
#100;
SIGNAL_A = 14'b11001001111000;
SIGNAL_B = 14'b01100000001010;
#100;
SIGNAL_A = 14'b11001100110010;
SIGNAL_B = 14'b01100001111101;
#100;
SIGNAL_A = 14'b11001111110000;
SIGNAL_B = 14'b01100011101000;
#100;
SIGNAL_A = 14'b11010010110001;
SIGNAL_B = 14'b01100101001100;
#100;
SIGNAL_A = 14'b11010101110100;
SIGNAL_B = 14'b01100110101001;
#100;
SIGNAL_A = 14'b11011000111011;
SIGNAL_B = 14'b01100111111110;
#100;
SIGNAL_A = 14'b11011100000100;
SIGNAL_B = 14'b01101001001100;
#100;
SIGNAL_A = 14'b11011111001111;
SIGNAL_B = 14'b01101010010011;
#100;
SIGNAL_A = 14'b11100010011100;
SIGNAL_B = 14'b01101011010010;
#100;
SIGNAL_A = 14'b11100101101010;
SIGNAL_B = 14'b01101100001001;
#100;
SIGNAL_A = 14'b11101000111011;
SIGNAL_B = 14'b01101100111010;
#100;
SIGNAL_A = 14'b11101100001101;
SIGNAL_B = 14'b01101101100011;
#100;
SIGNAL_A = 14'b11101111011111;
SIGNAL_B = 14'b01101110000100;
#100;
SIGNAL_A = 14'b11110010110011;
SIGNAL_B = 14'b01101110011111;
#100;
SIGNAL_A = 14'b11110110001000;
SIGNAL_B = 14'b01101110110010;
#100;
SIGNAL_A = 14'b11111001011101;
SIGNAL_B = 14'b01101110111110;
#100;
SIGNAL_A = 14'b11111100110010;
SIGNAL_B = 14'b01101111000011;
#100;
SIGNAL_A = 14'b00000000000110;
SIGNAL_B = 14'b01101111000000;
#100;
SIGNAL_A = 14'b00000011011011;
SIGNAL_B = 14'b01101110110111;
#100;
SIGNAL_A = 14'b00000110110000;
SIGNAL_B = 14'b01101110100111;
#100;
SIGNAL_A = 14'b00001010000100;
SIGNAL_B = 14'b01101110010000;
#100;
SIGNAL_A = 14'b00001101010111;
SIGNAL_B = 14'b01101101110011;
#100;
SIGNAL_A = 14'b00010000101001;
SIGNAL_B = 14'b01101101001111;
#100;
SIGNAL_A = 14'b00010011111010;
SIGNAL_B = 14'b01101100100100;
#100;
SIGNAL_A = 14'b00010111001010;
SIGNAL_B = 14'b01101011110011;
#100;
SIGNAL_A = 14'b00011010011000;
SIGNAL_B = 14'b01101010111011;
#100;
SIGNAL_A = 14'b00011101100101;
SIGNAL_B = 14'b01101001111101;
#100;
SIGNAL_A = 14'b00100000101111;
SIGNAL_B = 14'b01101000111010;
#100;
SIGNAL_A = 14'b00100011110111;
SIGNAL_B = 14'b01100111110000;
#100;
SIGNAL_A = 14'b00100110111101;
SIGNAL_B = 14'b01100110100000;
#100;
SIGNAL_A = 14'b00101010000001;
SIGNAL_B = 14'b01100101001011;
#100;
SIGNAL_A = 14'b00101101000010;
SIGNAL_B = 14'b01100011110000;
#100;
SIGNAL_A = 14'b00110000000000;
SIGNAL_B = 14'b01100010010000;
#100;
SIGNAL_A = 14'b00110010111011;
SIGNAL_B = 14'b01100000101011;
#100;
SIGNAL_A = 14'b00110101110011;
SIGNAL_B = 14'b01011111000000;
#100;
SIGNAL_A = 14'b00111000101000;
SIGNAL_B = 14'b01011101010001;
#100;
SIGNAL_A = 14'b00111011011001;
SIGNAL_B = 14'b01011011011101;
#100;
SIGNAL_A = 14'b00111110000111;
SIGNAL_B = 14'b01011001100100;
#100;
SIGNAL_A = 14'b01000000110001;
SIGNAL_B = 14'b01010111100111;
#100;
SIGNAL_A = 14'b01000011011000;
SIGNAL_B = 14'b01010101100101;
#100;
SIGNAL_A = 14'b01000101111010;
SIGNAL_B = 14'b01010011011111;
#100;
SIGNAL_A = 14'b01001000011000;
SIGNAL_B = 14'b01010001010110;
#100;
SIGNAL_A = 14'b01001010110010;
SIGNAL_B = 14'b01001111001000;
#100;
SIGNAL_A = 14'b01001101001000;
SIGNAL_B = 14'b01001100110111;
#100;
SIGNAL_A = 14'b01001111011001;
SIGNAL_B = 14'b01001010100011;
#100;
SIGNAL_A = 14'b01010001100110;
SIGNAL_B = 14'b01001000001011;
#100;
SIGNAL_A = 14'b01010011101111;
SIGNAL_B = 14'b01000101110001;
#100;
SIGNAL_A = 14'b01010101110010;
SIGNAL_B = 14'b01000011010011;
#100;
SIGNAL_A = 14'b01010111110001;
SIGNAL_B = 14'b01000000110011;
#100;
SIGNAL_A = 14'b01011001101011;
SIGNAL_B = 14'b00111110010000;
#100;
SIGNAL_A = 14'b01011010011111;
SIGNAL_B = 14'b00111100011011;
#100;
SIGNAL_A = 14'b01011100001110;
SIGNAL_B = 14'b00110111110100;
#100;
SIGNAL_A = 14'b01011101110101;
SIGNAL_B = 14'b00110011001101;
#100;
SIGNAL_A = 14'b01011111010011;
SIGNAL_B = 14'b00101110100101;
#100;
SIGNAL_A = 14'b01100000101000;
SIGNAL_B = 14'b00101001111101;
#100;
SIGNAL_A = 14'b01100001110100;
SIGNAL_B = 14'b00100101010110;
#100;
SIGNAL_A = 14'b01100010110111;
SIGNAL_B = 14'b00100000101111;
#100;
SIGNAL_A = 14'b01100011110010;
SIGNAL_B = 14'b00011100001001;
#100;
SIGNAL_A = 14'b01100100100100;
SIGNAL_B = 14'b00010111100100;
#100;
SIGNAL_A = 14'b01100101001100;
SIGNAL_B = 14'b00010011000001;
#100;
SIGNAL_A = 14'b01100101101101;
SIGNAL_B = 14'b00001110011111;
#100;
SIGNAL_A = 14'b01100110000100;
SIGNAL_B = 14'b00001001111111;
#100;
SIGNAL_A = 14'b01100110010011;
SIGNAL_B = 14'b00000101100001;
#100;
SIGNAL_A = 14'b01100110011001;
SIGNAL_B = 14'b00000001000110;
#100;
SIGNAL_A = 14'b01100110010111;
SIGNAL_B = 14'b11111100101111;
#100;
SIGNAL_A = 14'b01100110001101;
SIGNAL_B = 14'b11111000011001;
#100;
SIGNAL_A = 14'b01100101111010;
SIGNAL_B = 14'b11110100000111;
#100;
SIGNAL_A = 14'b01100101011111;
SIGNAL_B = 14'b11101111111000;
#100;
SIGNAL_A = 14'b01100100111100;
SIGNAL_B = 14'b11101011101101;
#100;
SIGNAL_A = 14'b01100100010001;
SIGNAL_B = 14'b11100111100110;
#100;
SIGNAL_A = 14'b01100011011110;
SIGNAL_B = 14'b11100011100011;
#100;
SIGNAL_A = 14'b01100010100100;
SIGNAL_B = 14'b11011111100100;
#100;
SIGNAL_A = 14'b01100001100010;
SIGNAL_B = 14'b11011011101010;
#100;
SIGNAL_A = 14'b01100000011000;
SIGNAL_B = 14'b11010111110100;
#100;
SIGNAL_A = 14'b01011111001000;
SIGNAL_B = 14'b11010100000100;
#100;
SIGNAL_A = 14'b01011101110000;
SIGNAL_B = 14'b11010000011000;
#100;
SIGNAL_A = 14'b01011100010001;
SIGNAL_B = 14'b11001100110010;
#100;
SIGNAL_A = 14'b01011010101011;
SIGNAL_B = 14'b11001001010010;
#100;
SIGNAL_A = 14'b01011000111111;
SIGNAL_B = 14'b11000101110111;
#100;
SIGNAL_A = 14'b01010111001100;
SIGNAL_B = 14'b11000010100010;
#100;
SIGNAL_A = 14'b01010101010011;
SIGNAL_B = 14'b10111111010011;
#100;
SIGNAL_A = 14'b01010011010011;
SIGNAL_B = 14'b10111100001010;
#100;
SIGNAL_A = 14'b01010001001110;
SIGNAL_B = 14'b10111001000111;
#100;
SIGNAL_A = 14'b01001111000011;
SIGNAL_B = 14'b10110110001011;
#100;
SIGNAL_A = 14'b01001100110011;
SIGNAL_B = 14'b10110011010101;
#100;
SIGNAL_A = 14'b01001010011101;
SIGNAL_B = 14'b10110000100110;
#100;
SIGNAL_A = 14'b01001000000010;
SIGNAL_B = 14'b10101101111101;
#100;
SIGNAL_A = 14'b01000101100010;
SIGNAL_B = 14'b10101011011100;
#100;
SIGNAL_A = 14'b01000010111101;
SIGNAL_B = 14'b10101001000001;
#100;
SIGNAL_A = 14'b01000000010100;
SIGNAL_B = 14'b10100110101101;
#100;
SIGNAL_A = 14'b00111101100110;
SIGNAL_B = 14'b10100100100001;
#100;
SIGNAL_A = 14'b00111010110101;
SIGNAL_B = 14'b10100010011011;
#100;
SIGNAL_A = 14'b00110111111111;
SIGNAL_B = 14'b10100000011101;
#100;
SIGNAL_A = 14'b00110101000110;
SIGNAL_B = 14'b10011110100110;
#100;
SIGNAL_A = 14'b00110010001001;
SIGNAL_B = 14'b10011100110111;
#100;
SIGNAL_A = 14'b00101111001001;
SIGNAL_B = 14'b10011011001110;
#100;
SIGNAL_A = 14'b00101100000110;
SIGNAL_B = 14'b10011001101101;
#100;
SIGNAL_A = 14'b00101001000000;
SIGNAL_B = 14'b10011000010100;
#100;
SIGNAL_A = 14'b00100101111000;
SIGNAL_B = 14'b10010111000010;
#100;
SIGNAL_A = 14'b00100010101101;
SIGNAL_B = 14'b10010101110111;
#100;
SIGNAL_A = 14'b00011111100000;
SIGNAL_B = 14'b10010100110100;
#100;
SIGNAL_A = 14'b00011100010010;
SIGNAL_B = 14'b10010011111000;
#100;
SIGNAL_A = 14'b00011001000001;
SIGNAL_B = 14'b10010011000100;
#100;
SIGNAL_A = 14'b00010101101111;
SIGNAL_B = 14'b10010010010111;
#100;
SIGNAL_A = 14'b00010010011100;
SIGNAL_B = 14'b10010001110001;
#100;
SIGNAL_A = 14'b00001111001000;
SIGNAL_B = 14'b10010001010011;
#100;
SIGNAL_A = 14'b00001011110011;
SIGNAL_B = 14'b10010000111100;
#100;
SIGNAL_A = 14'b00001000011110;
SIGNAL_B = 14'b10010000101100;
#100;
SIGNAL_A = 14'b00000101001000;
SIGNAL_B = 14'b10010000100011;
#100;
SIGNAL_A = 14'b00000001110010;
SIGNAL_B = 14'b10010000100010;
#100;
SIGNAL_A = 14'b11111110011101;
SIGNAL_B = 14'b10010000100111;
#100;
SIGNAL_A = 14'b11111011000111;
SIGNAL_B = 14'b10010000110100;
#100;
SIGNAL_A = 14'b11110111110010;
SIGNAL_B = 14'b10010001000111;
#100;
SIGNAL_A = 14'b11110100011101;
SIGNAL_B = 14'b10010001100001;
#100;
SIGNAL_A = 14'b11110001001010;
SIGNAL_B = 14'b10010010000010;
#100;
SIGNAL_A = 14'b11101101110111;
SIGNAL_B = 14'b10010010101001;
#100;
SIGNAL_A = 14'b11101010100110;
SIGNAL_B = 14'b10010011010111;
#100;
SIGNAL_A = 14'b11100111010110;
SIGNAL_B = 14'b10010100001100;
#100;
SIGNAL_A = 14'b11100100001000;
SIGNAL_B = 14'b10010101000110;
#100;
SIGNAL_A = 14'b11100000111011;
SIGNAL_B = 14'b10010110000111;
#100;
SIGNAL_A = 14'b11011101110001;
SIGNAL_B = 14'b10010111001110;
#100;
SIGNAL_A = 14'b11011010101001;
SIGNAL_B = 14'b10011000011011;
#100;
SIGNAL_A = 14'b11010111100011;
SIGNAL_B = 14'b10011001101101;
#100;
SIGNAL_A = 14'b11010100100000;
SIGNAL_B = 14'b10011011000110;
#100;
SIGNAL_A = 14'b11010001100000;
SIGNAL_B = 14'b10011100100011;
#100;
SIGNAL_A = 14'b11001110100010;
SIGNAL_B = 14'b10011110000110;
#100;
SIGNAL_A = 14'b11001011101000;
SIGNAL_B = 14'b10011111101111;
#100;
SIGNAL_A = 14'b11001000110001;
SIGNAL_B = 14'b10100001011100;
#100;
SIGNAL_A = 14'b11000101111101;
SIGNAL_B = 14'b10100011001110;
#100;
SIGNAL_A = 14'b11000011001101;
SIGNAL_B = 14'b10100101000101;
#100;
SIGNAL_A = 14'b11000000100000;
SIGNAL_B = 14'b10100111000000;
#100;
SIGNAL_A = 14'b10111101110111;
SIGNAL_B = 14'b10101001000000;
#100;
SIGNAL_A = 14'b10111011010010;
SIGNAL_B = 14'b10101011000100;
#100;
SIGNAL_A = 14'b10111000110001;
SIGNAL_B = 14'b10101101001100;
#100;
SIGNAL_A = 14'b10110110010100;
SIGNAL_B = 14'b10101111011000;
#100;
SIGNAL_A = 14'b10110011111011;
SIGNAL_B = 14'b10110001101000;
#100;
SIGNAL_A = 14'b10110001100111;
SIGNAL_B = 14'b10110011111011;
#100;
SIGNAL_A = 14'b10101111010111;
SIGNAL_B = 14'b10110110010010;
#100;
SIGNAL_A = 14'b10101101001100;
SIGNAL_B = 14'b10111000101100;
#100;
SIGNAL_A = 14'b10101011000101;
SIGNAL_B = 14'b10111011001000;
#100;
SIGNAL_A = 14'b10101001000011;
SIGNAL_B = 14'b10111101101000;
#100;
SIGNAL_A = 14'b10100111000110;
SIGNAL_B = 14'b11000000001010;
#100;
SIGNAL_A = 14'b10100101110011;
SIGNAL_B = 14'b11000010000011;
#100;
SIGNAL_A = 14'b10100100000001;
SIGNAL_B = 14'b11000110101010;
#100;
SIGNAL_A = 14'b10100010010111;
SIGNAL_B = 14'b11001011010010;
#100;
SIGNAL_A = 14'b10100000110110;
SIGNAL_B = 14'b11001111111010;
#100;
SIGNAL_A = 14'b10011111011110;
SIGNAL_B = 14'b11010100100011;
#100;
SIGNAL_A = 14'b10011110001111;
SIGNAL_B = 14'b11011001001011;
#100;
SIGNAL_A = 14'b10011101001001;
SIGNAL_B = 14'b11011101110011;
#100;
SIGNAL_A = 14'b10011100001100;
SIGNAL_B = 14'b11100010011010;
#100;
SIGNAL_A = 14'b10011011011000;
SIGNAL_B = 14'b11100111000000;
#100;
SIGNAL_A = 14'b10011010101100;
SIGNAL_B = 14'b11101011100100;
#100;
SIGNAL_A = 14'b10011010001001;
SIGNAL_B = 14'b11110000000111;
#100;
SIGNAL_A = 14'b10011001101111;
SIGNAL_B = 14'b11110100101000;
#100;
SIGNAL_A = 14'b10011001011101;
SIGNAL_B = 14'b11111001000111;
#100;
SIGNAL_A = 14'b10011001010100;
SIGNAL_B = 14'b11111101100100;
#100;
SIGNAL_A = 14'b10011001010100;
SIGNAL_B = 14'b00000001111101;
#100;
SIGNAL_A = 14'b10011001011100;
SIGNAL_B = 14'b00000110010100;
#100;
SIGNAL_A = 14'b10011001101100;
SIGNAL_B = 14'b00001010101000;
#100;
SIGNAL_A = 14'b10011010000101;
SIGNAL_B = 14'b00001110111000;
#100;
SIGNAL_A = 14'b10011010100101;
SIGNAL_B = 14'b00010011000101;
#100;
SIGNAL_A = 14'b10011011001110;
SIGNAL_B = 14'b00010111001110;
#100;
SIGNAL_A = 14'b10011011111110;
SIGNAL_B = 14'b00011011010011;
#100;
SIGNAL_A = 14'b10011100110111;
SIGNAL_B = 14'b00011111010100;
#100;
SIGNAL_A = 14'b10011101110111;
SIGNAL_B = 14'b00100011010000;
#100;
SIGNAL_A = 14'b10011110111110;
SIGNAL_B = 14'b00100111001000;
#100;
SIGNAL_A = 14'b10100000001101;
SIGNAL_B = 14'b00101010111010;
#100;
SIGNAL_A = 14'b10100001100011;
SIGNAL_B = 14'b00101110101000;
#100;
SIGNAL_A = 14'b10100011000000;
SIGNAL_B = 14'b00110010010000;
#100;
SIGNAL_A = 14'b10100100100100;
SIGNAL_B = 14'b00110101110011;
#100;
SIGNAL_A = 14'b10100110001110;
SIGNAL_B = 14'b00111001010000;
#100;
SIGNAL_A = 14'b10101000000000;
SIGNAL_B = 14'b00111100100111;
#100;
SIGNAL_A = 14'b10101001110111;
SIGNAL_B = 14'b00111111111000;
#100;
SIGNAL_A = 14'b10101011110101;
SIGNAL_B = 14'b01000011000100;
#100;
SIGNAL_A = 14'b10101101111001;
SIGNAL_B = 14'b01000110001001;
#100;
SIGNAL_A = 14'b10110000000010;
SIGNAL_B = 14'b01001001000111;
#100;
SIGNAL_A = 14'b10110010010001;
SIGNAL_B = 14'b01001100000000;
#100;
SIGNAL_A = 14'b10110100100110;
SIGNAL_B = 14'b01001110110001;
#100;
SIGNAL_A = 14'b10110111000000;
SIGNAL_B = 14'b01010001011100;
#100;
SIGNAL_A = 14'b10111001011111;
SIGNAL_B = 14'b01010100000000;
#100;
SIGNAL_A = 14'b10111100000010;
SIGNAL_B = 14'b01010110011101;
#100;
SIGNAL_A = 14'b10111110101011;
SIGNAL_B = 14'b01011000110100;
#100;
SIGNAL_A = 14'b11000001010111;
SIGNAL_B = 14'b01011011000011;
#100;
SIGNAL_A = 14'b11000100001000;
SIGNAL_B = 14'b01011101001010;
#100;
SIGNAL_A = 14'b11000110111101;
SIGNAL_B = 14'b01011111001011;
#100;
SIGNAL_A = 14'b11001001110110;
SIGNAL_B = 14'b01100001000101;
#100;
SIGNAL_A = 14'b11001100110010;
SIGNAL_B = 14'b01100010110111;
#100;
SIGNAL_A = 14'b11001111110001;
SIGNAL_B = 14'b01100100100010;
#100;
SIGNAL_A = 14'b11010010110100;
SIGNAL_B = 14'b01100110000101;
#100;
SIGNAL_A = 14'b11010101111001;
SIGNAL_B = 14'b01100111100001;
#100;
SIGNAL_A = 14'b11011001000001;
SIGNAL_B = 14'b01101000110101;
#100;
SIGNAL_A = 14'b11011100001100;
SIGNAL_B = 14'b01101010000010;
#100;
SIGNAL_A = 14'b11011111011000;
SIGNAL_B = 14'b01101011001000;
#100;
SIGNAL_A = 14'b11100010100111;
SIGNAL_B = 14'b01101100000110;
#100;
SIGNAL_A = 14'b11100101110111;
SIGNAL_B = 14'b01101100111101;
#100;
SIGNAL_A = 14'b11101001001001;
SIGNAL_B = 14'b01101101101100;
#100;
SIGNAL_A = 14'b11101100011100;
SIGNAL_B = 14'b01101110010100;
#100;
SIGNAL_A = 14'b11101111110001;
SIGNAL_B = 14'b01101110110101;
#100;
SIGNAL_A = 14'b11110011000110;
SIGNAL_B = 14'b01101111001110;
#100;
SIGNAL_A = 14'b11110110011100;
SIGNAL_B = 14'b01101111100000;
#100;
SIGNAL_A = 14'b11111001110010;
SIGNAL_B = 14'b01101111101011;
#100;
SIGNAL_A = 14'b11111101001001;
SIGNAL_B = 14'b01101111101111;
#100;
SIGNAL_A = 14'b00000000011110;
SIGNAL_B = 14'b01101111101011;
#100;
SIGNAL_A = 14'b00000011110100;
SIGNAL_B = 14'b01101111100001;
#100;
SIGNAL_A = 14'b00000111001010;
SIGNAL_B = 14'b01101111010000;
#100;
SIGNAL_A = 14'b00001010100000;
SIGNAL_B = 14'b01101110111000;
#100;
SIGNAL_A = 14'b00001101110100;
SIGNAL_B = 14'b01101110011001;
#100;
SIGNAL_A = 14'b00010001000111;
SIGNAL_B = 14'b01101101110011;
#100;
SIGNAL_A = 14'b00010100011010;
SIGNAL_B = 14'b01101101000111;
#100;
SIGNAL_A = 14'b00010111101010;
SIGNAL_B = 14'b01101100010100;
#100;
SIGNAL_A = 14'b00011010111010;
SIGNAL_B = 14'b01101011011011;
#100;
SIGNAL_A = 14'b00011110000111;
SIGNAL_B = 14'b01101010011100;
#100;
SIGNAL_A = 14'b00100001010010;
SIGNAL_B = 14'b01101001010111;
#100;
SIGNAL_A = 14'b00100100011011;
SIGNAL_B = 14'b01101000001100;
#100;
SIGNAL_A = 14'b00100111100010;
SIGNAL_B = 14'b01100110111011;
#100;
SIGNAL_A = 14'b00101010100111;
SIGNAL_B = 14'b01100101100100;
#100;
SIGNAL_A = 14'b00101101101000;
SIGNAL_B = 14'b01100100001000;
#100;
SIGNAL_A = 14'b00110000100111;
SIGNAL_B = 14'b01100010100110;
#100;
SIGNAL_A = 14'b00110011100011;
SIGNAL_B = 14'b01100001000000;
#100;
SIGNAL_A = 14'b00110110011100;
SIGNAL_B = 14'b01011111010100;
#100;
SIGNAL_A = 14'b00111001010001;
SIGNAL_B = 14'b01011101100011;
#100;
SIGNAL_A = 14'b00111100000011;
SIGNAL_B = 14'b01011011101101;
#100;
SIGNAL_A = 14'b00111110110001;
SIGNAL_B = 14'b01011001110010;
#100;
SIGNAL_A = 14'b01000001011011;
SIGNAL_B = 14'b01010111110100;
#100;
SIGNAL_A = 14'b01000100000010;
SIGNAL_B = 14'b01010101110001;
#100;
SIGNAL_A = 14'b01000110100101;
SIGNAL_B = 14'b01010011101001;
#100;
SIGNAL_A = 14'b01001001000011;
SIGNAL_B = 14'b01010001011110;
#100;
SIGNAL_A = 14'b01001011011110;
SIGNAL_B = 14'b01001111001111;
#100;
SIGNAL_A = 14'b01001101110100;
SIGNAL_B = 14'b01001100111101;
#100;
SIGNAL_A = 14'b01010000000101;
SIGNAL_B = 14'b01001010100111;
#100;
SIGNAL_A = 14'b01010010010010;
SIGNAL_B = 14'b01001000001110;
#100;
SIGNAL_A = 14'b01010100011010;
SIGNAL_B = 14'b01000101110010;
#100;
SIGNAL_A = 14'b01010110011110;
SIGNAL_B = 14'b01000011010010;
#100;
SIGNAL_A = 14'b01011000011101;
SIGNAL_B = 14'b01000000110001;
#100;
SIGNAL_A = 14'b01011010001101;
SIGNAL_B = 14'b00111110011010;
#100;
SIGNAL_A = 14'b01011011100101;
SIGNAL_B = 14'b00111010111100;
#100;
SIGNAL_A = 14'b01011101010010;
SIGNAL_B = 14'b00110110010100;
#100;
SIGNAL_A = 14'b01011110110101;
SIGNAL_B = 14'b00110001101011;
#100;
SIGNAL_A = 14'b01100000010000;
SIGNAL_B = 14'b00101101000010;
#100;
SIGNAL_A = 14'b01100001100010;
SIGNAL_B = 14'b00101000011010;
#100;
SIGNAL_A = 14'b01100010101011;
SIGNAL_B = 14'b00100011110010;
#100;
SIGNAL_A = 14'b01100011101100;
SIGNAL_B = 14'b00011111001010;
#100;
SIGNAL_A = 14'b01100100100011;
SIGNAL_B = 14'b00011010100011;
#100;
SIGNAL_A = 14'b01100101010010;
SIGNAL_B = 14'b00010101111110;
#100;
SIGNAL_A = 14'b01100101111000;
SIGNAL_B = 14'b00010001011010;
#100;



end


endmodule




