// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 15:05:46 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nijkUuKbactz0qqkM4OY7QmZycL6LlyLFBzv2Qp1Kke36wSDoC2jX3T8QX65zpyE
PBf5mebtG3lxcPUOphKkL6CLFCwMx9yrLdEm0bRNAKoXbQvgeE/XES1AkwjJ33oz
YCsCkiRcw2sE3tNxa7GqK2KSmLg2xdAWOaECOnMgq3M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21296)
EDdN59aq9m7lkh8X0iYCj/KxTN4AZLy57OKvujWN/u6wPgaJb3kV9qwXbiWH8xr+
gF5gzWDB1v6xzbyv5iiaisEjmpqdHDSsU3IrBpBY7fvwy2pf9G1mzIbTVoV5yj/V
Hxsf0WS1vlWnnHgA76NK8oQzo3Fy9hx/brFNYoxdAMmt+0c2Po/k1d7n2SbA03M6
KK2ji1O/sYRJTWbDDYvpjkFjUiOBCqvNtZk8omakM18y5Ute0OnmRi+GlSqyUfL0
n89AAsIkFJZTVvcSbuJrHq/S619YCTc5dWQcsIQ0NdoIw77pViMDs7TnajRmo4Ec
cyjZ0Wje8SOSRnSd4DzDXdPLhnBdp/8owduPyX/7Qy/uuXiBcq9xgxGK2P4dXd4Q
Hu7qThb2/yGAqS2z4fP5EqKAyZQ+euqVdszXHfMxjrQUg52Fbon2aXrK2YRzYdxR
yu4+eusStlsmZVJo7XK1gIZfdoCW1XWbyGsmbe0XZV1yBTB5JMsuJXZ7YWc/ZRzT
8+xCdzE2xf5bUmGq9Mjs3rfDeszI/I+Uu5oN7sw+GpMZpXf00fB6egC0nP567u3F
7BZ9OgMAePONQalaJsqYaMPOSp09e7nlt+8C9lH07903/SR18cQC1+75OvHhmmZZ
PdAIjnqOVIBtINuy+coa+nlHDWy0/wbs55NZp2K9FDkeIxn06xVoU9ZdAFzrF+i1
BjX7bgcpq3hQuBkiINoFWT2mp/b5I5zTO9ngIWiMCX6mJeNmiUecSwAKnj24H6Ve
cJdTa8p9+kIW7IdmAP6ZGNJ630hVTksBt7rLCxzx9+n9KGcX5sg4qDtwzVz7uk1v
137fl7lNkUIo3GUsumrUB9D99YVCpLsD6FZUAhoFQ8had5ZAgOZxGxxrZ4m1liJj
OzYBUZNCPywpJT6RFve1agqlhDOMmc4DDjIwO/0coFIEondXpBk+CjEEEfhTbXCb
GGcrDYQrPRJAYZ+wLlN/ufyiAiJou0LFTdc1N6sAan/lvv1fsW7kE2ut1nyOrAAh
z3gza4EXCDNq7c28CwQtBYQyXJ9Oi32BpGs+3hNjSVnWyZ7FChePUjA/CSg2LtNj
0LFbM/6PvtNRRvAlEn32rHrwRycDAapBYGkL58b32Ohdp7qgmN6Sc5JwRICuvgag
VT6uFeEtUIR9Lxf5LsH4llCPKRz+oOpioVCLnwzi/8/EjADS14zXmdcg1HFX0eCp
9DSGLvl6lXsuhceOTec0S8LyJpcamXdz3jmhOWBR8hAAoJGg4UT1JsfVau5UIRzV
lA1mI3R4TCdsYiqdzaY+CIhofSxnUVlO55n9L4ixnZhezdwCEpbWHubv9nqzOVFT
bNL95ssaPQl9L1Vc79CSG1ZEB6F4zpsF54MvAx8GeT76Rf30AO9Dy2ZcwzMldPAu
ZhW2Kl/dRx6PuTq9lcuhT6/lnlQlVc4ttiu4BSXJiHx6dAZDHdu3WAunGWmPOhFC
fW2D6+3i/q7a9Zq6mtfP3IieJt0mOKlrCmYFcEj7147l/WlxrkXfx74AONZ5Mw02
MzMoiK/2oRthm8vQsJNZnRRENIsGESBGsWJjBsh3b3HE4VCLOQXdKAs8hoo3ju9u
xexoNUDH3AWmzO6mMDgjsk4ybJBjknw/R37o16qSryCluyPfAp7zF6/whr3baSDO
ZnMWlHlqGsVR4kex+RfJfM/jSS2z04/v6VtsQfXT7dPihFHf9vX9XD+FND7JpMoK
NUkrE0D/NxzhJnyutN85q6WT7y9YwVZnexh3IFj+Ki6pk9nN97dLDRXuPTK/XWdj
dW+QkFKKtrIuiVBva91yWgRWnyPADs2icpZlbRD8hLS+PCDVQOPOb2f0RwUCJZnm
Zh7r/SW0vJ1+fAGWy5yS4Qw9eCzx5FitxdWPu0Ngcv54S4fIdzVvWOfn/AMCWWre
t7EN/1xcG6gZolELoSSbuohePiBpHrxZ3l31VEwBpsZMYBGafp+zL2RHVPxIzjpy
OcMwF0Hm6RDj3lq42SaLV2BCUyOtgu+VGNKxG3KBeGzGrtvUtRE3iTSv/KPGBG9S
zHDegtRW6M4NugZMLlyWF61FaZVa9JLWX8TB5GBgNYBgmCobw89AdlMXmOtHKOoa
Ahf/UPnZxtWTKN+8oE+La9AUIT14nRLPg7IcbSJveUMQZLB89DFoT0m8IQzAaeIM
G8nrrEs0On/cPf7/zGZcbMF2DBo1I421dF5Tv0uIamNxaMz3DEn7RkXdSk+bDJ+Z
tB1iuMEQUwipkypZl0G1IfELdN1cxvc3bctyLME/m6fUBZUu0JHs4aPLgScCmZdB
5qWXpQFHioFr46M55Pnpz913w7BPYUZhIqw7J3mdZSWXi9ySHi6+tSfB5YV0RYEN
Vi+6g5wzL/7JT47qkN/Q95E956Z0No3rAC3zVf/6MVy774OypH3yBgP3GmvFvG+l
A92v+chWWyfCZdhnDlmmiTgiHuZ47j4tD4YwmVtgoj1FLycEjq+A42i3q00uvM9K
MTh52MaJ2sKb0xUdSZTdqtnJoxhiFq40cZWYCzSmVbXy+6LZlrenL+6VQAU0TmT3
Su7lbVRe07FlfpWWovUpCUMzSbplXOGoGMNp1ZMvuMGE9bcnyhlErzcN0iF8WWdI
g0Ke8R1Ef2QKQm47MUaLRilPhfn6LZrVrgZrzXjgtJttKB8MNdbl7pYHC3H4m5a4
usbNG4x04oX6ue9z9he0A4gYnyKaZfEKUEiK26XD6UXm5Ag/88e85HACnBxPpC6L
i0Qh/7vY97dQMmcVwneUFEhDtX79qqFa2j5+xhB+mHp2v31u/IS/qk4NMO24T+EA
lNasXBD/5lGSDiHcJXtk2kzAsGyVsmCHve5hVT75TEGs1YzOSaOayNxQ5PjUACyJ
F+LRCgli+1iBM0wL0h+fbGiZVkrtAFVrw1HRFiXa6AGkLvffh/vBFbfHzwn58tNW
4q3sWorT3XxSPSRtQSUV3OpwIdJzxhv4+f5mb19RZ3HYbR2Udb9tx5zTMHTBrppy
TpDbfnD0ebBtPI+jF4wOPA6kKOlOVRWTHOeVRTUQrS+WFyqv/cjVORA46uYx8buD
mWV9ghm0CYpzMpTOaBGD5OJ6sghQiGl87o1RHHQ1qLL2exDXE4XniipIz27166gT
k0PJa2NaB1+0x1uMOP9L0qOZE5DqXRPpTvMbJX3xRM2kpXaur0B801G/tTtB4S/C
vaH/7Y9XOxSa4IJlHrBwTOCoqmPYyidW+W6aqhavV3nMXPNXTsVigFC9GnRvRwKU
N/lbxsaD53/i6fAM6Y/+dzDaSFIh3rYVjMgMm7um1TYIof6yJZgRNJq+/37dIHa+
ZcaJ23/ftXO5ze52mTfTGtZZvbwdt1H+l+ccqzgJ5FLYw9csZM0xApiuQymhUI9T
XsPQaFqiVedDVe2VSa53/o/6IZ6ZzRgUcrv/Z/KZBtUPqBxxPUGmCtnPv+mD6daP
9geapqloEluud9WXd67krmU2Hk4Lu/B8QU/q6b2KS7xotfMLUSGDQf/B4ypR5uUZ
YTaGcenyfGblhjL7isjMOX9nrxV8VCFBX/S4RY2E7HtTVL73bPGBVIdqIOcw/TdI
Zxj05XsJKWpQyktyW6oG5TiK6HnHvQPJedpMReIALuG3oumDaU9Da5WCuIYVpkIQ
gWu0IbGDGUlT0EKJd8sSJTdA/ZKBdur8AmnqNiFPUKAiVwiNdILFTD8161W8gq2N
IkdTd1AwRmKzbleRVppSdX937VyhA2DC/QaWum/LbYNpp/XDES4uFhOB1qIkoH3g
KOV4QP0esxSJjKqkN1btdy6WpvRkNO1yBNeucgpC3Hh/Ih1W0pZB/1cL3QpRracX
+zSt+uO3f5E1/WkPive8gAhDUGPco8sA7496njoYVf2zPzX56hyutvEdhj+gqi0E
sWOk7fD3z/9OIChnT+Kh8+aR4AKZFyLvkCD8aQXq2eeb6p5sPQlv123Jfc5YmQNQ
dPfF+AwFgqsNFBhwl5emtda18C9iF9gJ5pHgQWcRBVB/Rt2e2gx8TmzS0Zqak8d/
TEVUxZGxRmQ8mPOEfMTgupIS6XOw0rGlNugDfgM88wEWFOwZ0bI7gaLqNgoXjihh
07n2cCe/mdT7UQL8RoNn+oPYVMzBiowuDarYlC0VaaG8pqUFlciRCn9UXAJlqS1U
GkcJeKXrsc+rtd4qYKfD4GF9yT38WdID+7a90RocfqJzS9eo9WJjNM2N6Xt/L/cX
lF9c+BR0v7vq0hrngI7bfp09qSXR7+1QwHqsXeX3IkmqMAt1LeWCKlpP6tNJ51Gh
k2dJqlaqd3BF2IhwJSoop4tZn3nzcIyKlPxJvEO8KhaoYM/LCJ8B5MWs9ggitvD8
nk7uT1lLHO+Vme5kFgvWUpCRnSKKl0gKiu55H3mWMvZwLZE/qk2ZTMnAS04Ezh5Q
AgtvQqxQar8wyMuYyRp9PARMKzGIY1oUc6iJ1pOhw1kDYutrWL4C3W5adBz4Ukep
IlR7TDW+S0J3e/uhg/Tu/H+sg0Yj4h9TJU6fKqe14P/VDMTjLiVn7etXuNnmICpQ
W5k5j9MAH8JxcXh15Rwbnak9RNo1fUG9B/t+hPJfBJMcslb48UEi9gLfLzau+wm6
Biz9e+1mu+/YmNH/11G0z/hhLNIi1tr99UiVu0GdXdvHNRFYYH4WevdjYm74i/BW
X/yk3M3N/GwDaFCEDBmXs89dscceDxTf1s8ueETeLCb/gDkGNO5mhzV7V2vrcXev
qs4hJIqSj+ZUL76RUquDWwGeSaCO5TC93sPRfLGjHAIKkkEYpTOjCKq4Td3+uYG/
UfHI+smLgmfF3FDxq6DPthTkPvq49W1k/+Gh7xApf7AOzkUjPPHu4EnTxXgqmnX4
/TF8ll0gQAGGxFiW6JIHddeCxGS1qPvNYfCgZogk8srvDoyx9Kjp6Z/ME3VFOb2M
H2zUsmu8mGpafLXws055kChBVIsXTRRvInP3Lh8cqOh7fHWvxZeWKl+CunO9qst+
SeHRlX+RD6kQFt4phh1i3ZhbfHOjivaIWgR7/jDlS5Y5VEGE2SAoqV/gJaBRXIGr
ltPkkaDa9EHD0axpXS+AXSIG74J6LsH1dsp9H52678loTMNavFCwssrGO0O7swD3
7/BNGNfrcQjH/XgQsVjagOLf2KYZtlMGgltCyzkkSxG3jDWTAC+NIs1LOWbIEUye
MpRrIF0VjaBKaYAFv4PnMPD1UxP6Fl8/Sv9q9rJHys/W2+STlp17rOOTLc6d/1CD
EafwMFD6fxVnhASyZWI1OYCuRUJ7n0f9dUkKL93a3Pi6HI6TLhgXbXC/HQdAtTmE
UnLRRNQqGMvTWcQNdvPtR0BcWRZrc340xSPziU7MlysNE8aZw735HRM4sQZDogxT
A/afLMMd5Ua7FXAzM3kuLIngvHEjC6dCs9UJyjTLvWtSHTqowo4ezuDbi6f98Jh1
p00yYN/3IdITpxI/4J119nj9faGiw6r3tR/8LYv90FnF/3qwHQtt7cKuTsq3Q7Xx
OeaDpaL3AZadehsBSvB7BENxSA2SytzfMIlK9nEBj+1OQVcyy3VkjCEeRK8oMUPi
ylIaRgv496+fbmyqYsnPFf7JJohKGVMiqCasiHdFsqENMXfIobvPwBCysONbb5dl
uaH8myQ6JSsJ4CZX3WG7RJ1SAxSoW6ZrERMYMrd4uEJ+u/Lu4x+EQIlEragEVGaX
JaVKhbXkDDpRXICmfRRu7X8gosP3p4EGN/NX6LtmlBFFDInDIb2o2w/exn05u3na
Yzj5/2Iq8V6dinWVfXGhLKBHLPQmPUMl4IAcxJBOBWRIMsLuWgs6+oJUeQe9ZbZr
CvJkwHgACaV0BREuh16VsXH3VStuh4h2oOsY3E2ykNHQIfGMfKYPewahgjB15ug5
+2M/c1mFGfwNq0lSj/RGcaVlHPoEABlyico5Z172somVpQBxk8zCnjC1WUNKtV9Q
9OxJEq+AZ9WESGbNsqSwf6vNZxmMfMSi+T40mESG7MPzlwMgwez5m7L17HJRrhCq
o9SuZWHQEPbxXE+8a4E6OqDiPujfm/hR60bp2rHUzlp89s+kdrBS0NL72AYGI2pO
Lv0N6Y7kdZngIKB1YGLeuTIARsEqllXLAIsfqo0VCz8KuK+v8iGh1qdBo30sJjGK
CITnEndvrBIXra1Ha9ipo26pqOQD6ev78VcRR0/WkhpuJKaJoJZJa/MONjtNU7bC
VeDu3lQv0EUukWHRiEL4hLUbUltpdbk93gNBnD3ewnlVklWRZ25htsZU5sPLFr4e
HQrZNwx0PVvam44+A/OhTmprNLxxALDR5pZW/bzjPs5iK9Dz9OHk3e+J002aYMfw
yc2yur8kDQhMhVz9dNYVU/b8r/KIbSxsv8zvQOO+7B6qNU1ZP1ZYEdZ6E1IvTPI8
dIt/eRKnZl2Ss6k9bCSHpktrfj0G6/fhhezAIHuzTVZjodsym71WzdfFSDhFCXTY
BUh9Da8otfMVHYUEVxsl5/58tYMR3VlFVHNIh/mRwhkLYa3QGpSMq+gcQlfWlvw9
mRxvYAk+J3OyU9dHXaAjW+3uGmhKUYQPM24yneDc7UA0E1AivLk1KqchS0v5UHV0
E4snwA80GKEXjDYCPc03hSTze464/eFotWIwvdhY+wHI71MKpf6XfNi8hG4CgfCr
U/8KMOyX8eN7q0X7V1gwLn1jvIx1HWGnmDcYNcmR7OICuiCRXZOWYZ9yTwdvUt4Y
aVCAEFcPmW3OWLsQgJMf9w4PI1A+5+M/sI2+m/Ec7ArRTXr+bVP/65cuBxioqQ/C
kW3DUouZFTpLyz8TZOS5IlrT5piEaFrJu0JBIT8wtm9qYKDG7Rn4ejCazvjIec8i
OY3TQTrZ614MPfbvBI4AgLPTSqz7zOjlyE2dW/tiiV4n/EWKKyF/r9+RqIDoi4e9
Zw9+gXX2gXp/y28m47Q5fGB1WgstyHUlq69BF+oMtnZDetLsAUoZNLB+Wp+/+qXl
Ar7IC8k8Ui/SEw3PDFFOYih2y9rj/vXxDlW+SeiNNMg5EJsngQnFr/A0V6UCj2Pt
g7pMFLbaIhEQlvJK9BGo2n0oTfs9jfgRS6Jdw50SFQLLqYXmptVEFv80YHWCT17P
aU+c/hxKNgScdMytSl3jhwkt+XijQU/nUOSBNQaRrG0TojjHBeu+6hhyXhZTANF+
X/SrcXCbsSS7Vwcp2xcEvLL7zK80WeBrYyWTAOY2+xaapqqeJW0HHTsFyz6vXD9l
iHNu/4++x1PSICU0sh2pz9zz23wXL7dXACGU53GdatZ59x1L+mfIROvTky8juZLL
ahL1ohs4X/ozuRhtuWulbla8ZKm0r6Aj5otikqZhEqxRq7HyzN394q8hbmqQW7wN
2LqAA6ORmT5pGh7p/nhtdskNtaUyf0RIeCJqN0It9ijwWpm73tpxI460CVVFtGua
E6FO6plB4GYgUap+S05fbAbAzulZc0mjN2IvWQorNd0W1r1g+ipg4SnE0Bo+KE0V
/9GrDLNpxviue5qRKK7yIoSIv9Yfhf4iEf/aLEeKwmBjb9Rt4Af638mij3w40Ibm
wpL4eppfYzm85E2lY60C2F7vhVFTMTkyroz2wpo3dxoVziy59eUqHomhNWGDKClV
jLkxmLmP0mJ03R44RVutEOolLwvPxbw6NO550fql//3Dewb7X3xRMH3LM6CTCuja
K+TEMefgpDJf1GePrfaOOoHG7QH+edqU+jVi76xduCQ8TWoH9PHsz5C1V+cQkmHl
sWZvg5ygOZGBNPr3+wh/24zgqM3Ud2yL6lnkR5ekdqtkiNYLjOBJm7Ta+ktRcQLq
VMihrwuxRvZMyHwjVcjV9IRVLZzQCj8GelgFONMNNtjj/I0DSXkO40MzLZQVghvM
+hFMBiQDAk87T03UAm/6wU9dnMaE9R68XVYRiUzXWr3n3LfhxDiKhXRXzK2WbxYx
xBAv2OrzCrN+9Eh3l0wUo0zLxMJrKI4nfcOdC2Il3owwqBQ2F7+eATLyFjLTc3Md
nStvUnr9m/rCpGnLIaQkno5V+JWm0evBzRACUw41cqGCGDUIAaWZ68iWw+7dQ0y3
Nqrnqdn14OoZ/8xwJsx6cYLs/YDEQD+f8o6Pmz6weq7bxqCtf8e02GU/V1CoQrMY
yXNXYl6jql0UoTPpzlM2/7oFt0n3CcGLp3xBqTfE43XFlri604z4caxlFFlGQ12L
l/M++R1T9TBS+iZBebxz6tr7cNRpZvil6EWbF7/S+c+kxYkPpfF4FPhte7+m0CxB
lpGA19EIguO1xDZE4Dq4kfgFnBUs57QgjV4FvRY5313v+0z2sh3lyz7vjZTSh4Ft
R7r8Aj1itcZNjer2N+w+osNJz03jgOOnGehQDNCaVVhCwjcIrTqIeKJnwNUBVpVs
pLb5aJC4tR6uRUrINCZ90qWNHcVvhePxV0PSecl1zY1Y+YZAKfqGvfM5yAK8v9JZ
nH2phwSzRd5xGFm0rSMdxM9JbIRdPPtuTKEInNSosTwTxTbfCdoilbZi9fC34skj
EVfVBJ0M76xuckr5MqYPKkU+E+RBmeA60BqnPM7HxSTa6OXQj2QSa7OevorNkTsg
f9fSCkKGfYyJ5YfOb/p9atX67FkmfTtcYrIdTWH3uZPlRmCqyxsTEQHA9zW/wL3N
igP3tVcxjd2QaYy+Htffe5UaNoobS4MYBVU1jIXB3iawDRpggQ/rCoAaIZ5iR2bU
U8R1bReuLKSEFSv76fPS7wkOJUnYjfHfKDx4piIyjeIP5yZkHfjH6T0o10WnZrLc
ADIW+mTQ8Hj0E6XsSTWNo7vCr5vb6laQ9rTd/WA6st5QHBi+7AXeMrLMvroxxUpn
34pHnPZVI2ziX/VEbKQayPqxc9R3OtgGPizVRe9G9o/AJ7JepI7cX15zY2rrQpfc
4ZTfaauX6qaU744tNs3jauKZQIBCJggMuP1ryMp0koH3QtqMH51jsHTOF/iO81Fq
T5jCfZbE2T7OQaYtD0j5PaeSDiWMPQlP/r0AZdjEsKkfGoBWAw7VzHsQClKBcxWw
colbamL5+H3KnkvbhnYsbl+VQ43yhJIAp6ao+v/CC/293a1GXTamLJcNEJGBa4ZV
gSAlLF1RqzNrRu1ibpa+SoxHd243VxQX4RQGDugpLeHSHEIkHY49b+OTWAutS2wl
p336SH6vyQjNGfWNYc/cTBJEdAmYqG+vhk+W/+lD94U8MPNunv1AI224LAcNammf
vL8UzLFdhckAVSmo8uCZMolcjOqSI7L/ucQ9sOBdS1Cv6+/jmIjzaqE6XK5V1tnx
h8df8K7ZPVdwPCGYnJ/a5li9v3cxEjHNPQpncqqJ7JISydLwTqSD1D+Y8onqqblX
deL6jnaW/1I69Jlz0HM9fpnM43vC2qhXhUvu0szpGhhTx8NzBXTsJRp5kzZ5E9UG
1GjTunA+2W8LWOmVDZRmFdo+/wZ26fFw1EzhOdoSxPUJ1GLiGIrbDTWrEPyO4wHa
C1LXzovBF+FZGHYZUauIRNtBAxbsQfgXE+K04Fo7ctHUC71imd4khP+2zGfeQflE
ymGmSf3R3qr5HkoXyh1ry1xHcSKI8SmM0Vqg3IqCJWuFIBrR+Gmp8CjMT7qSY1ZJ
I42jaXwJ35Blt8eYpcdKtVQpVYOQiLUVMoeZvDgvt2ixgv11a0pLfdYyvwTp+ix7
1fAtTL/IQjnoribUF+vMamLBQWnMN5EPOfRTWzueM6vy3brXdFx7PL8pgpalIF6z
zhTu/bGBo9ei17he/oyFm6Rv13HfD7fHuHIVJrMjgbfVywL49nlczNsPow6OlShB
UDLhhkVD5+sxu3K/+ZSE016421/2QJUdf8opWFeGtV5zKq1vtPQii1SuOmQ5Ah03
wuaS6E4M7TpqPT+93KHHVsnAhsDluquG2SLroME0BXs4RyMqQriQ9kjcSQJy0bdh
akC3tabhda8dpb56whsohglJOhAmG4hXkMs9TpSyR00EnCckfvoh3vBkK4XzEA9p
JYAFEjIFKF8PQb2khhC2q1WTMo74GwF4hhJeVaAieU05X7BU3/hcgK/l/cstEBj/
21GfPe5lWm7IUlDGFsy9VVvrF3zaT9L+lIabsLHN5msEB+Y07bDGwLg3l0MH80tg
XKOJoEM+EIKbKN7HOlF3ux51vTSCtv64aJupMB84zMPIlvvCpzHIszvvfeBXG4Hi
ugtSOK/CxKzl9NXh9hyMj+b+37zj2Rn3uBuHvayr2PYY+yhzdF0KzObuHE7LAwu9
fOTx++vhnUqkzUAZjlXqfAHnwRKzpae/IOapdRTdRU2jgXnULWyFof8uWp37uO+z
QSHY8qWMdqDlxp3PtX69rIZRO4trUAdmOSf7ohOQcCJo++ix9b9dBN70e6/m5KtO
TUgqJm7a3wBBjKHDo8ZoLdpHcALvbH2sCTC+dxLCnP8IixuHaFXyVOJFHILeg5Lg
LqToqCrkQuaqyJrkpGUhzMp7ecACUQxc3k7FfZNdTijzY/fE3Q5Qv1Y3hWtrcW2l
qi9c4okmSeBRUPBzPqARgqVM8jfjLhigxSCbM4MQaz/pvk6abXOcXDO7LefWJmrq
/zkH02tqr8SNxgwsmsi4ttg661DfSYPBOq9Oe+7bSn3uGKowRc9JB6Z7EbVQ6rjj
tLHmyVtObyKdJ7wCmOMPVq1AbtMVjtm19RuNH/Qm4xCEZdOM821As364KyOLbaq7
UfPxjgutoPsJwXrZGNhs4JYjXOgBQMnRfTJ4qhOjT0UdXGEBUx6Jn0HOIsLzbxNh
Sum0AvbWTGvlSR2r5m95EVafI5+oVSRatRMAQIOfEH76v2RuFIWpe3ZzMLumypcn
U81iamwuunJj231QwsqTZzw9AloA11VunmyCiHQiCaubi+SmljA/sufHkW0pq7FT
KoL2/OGjn6ujnEbVvyL7WerkEincTI8pWq+XzhGgdbzTZIWlFLvMHuDOlOSAj2RX
hIvfAeQ2fZksOLTLbAea8JJAWQttGnNj7oD6Kyeq4kmwRFY8fZtY8AEgmmVRzSg1
b+q7gHeCX7HaXYTg9ychbAmEDNblsL9l+Xa0hpYyvoMFfRS8brz2O/5snY+sz1ka
ZBKH500Bu8HB3OWqiHkPSJNhPz20CZsHmCkioumm4cgGONOFQU/Q4HE+CCZA2/VR
J9UHhOHhpXyzsnke7UZsWNOKTEEDm5fFMcESdoEi8gQEJuokIp7kaWJG6yIk7WzL
xLqFqAI88DWSdIJ1Xv42JhfqylAbhJAQN5yDjWn/H/jj8X6ihAougxMTxco8S1gV
eOg6ylDu4ypMc6A1IIJ//UxIloGxo8VG3ILjIos6jfdy22bS5FUfa6jJBbo03VIR
R1mLwKqiGME3otgy3xJdSMq7gBMxzH5PYDndR/NmlHLrBuQU2OsltfyD2e1fmSO1
XAf8zybFUXWCvqL/zb9/+NXNxmKKQ/fyVnUZw7Gfi6JoP5e+awccl3aTF1lHw34y
ajL/wEBDsTAtckSWhY8hvpDlttEF/nS5TAqA/Z42Qjrm12bORjhL7Zi9Cxh3FJcp
6KCdvub7zwEOrKs0tHmmmPH6hiwmYBeFjSDxpUYOc/cxRJ83F9yUOgNbteNy5ns6
xMyo4U0XYBOkpMVOT8ddM2HmaX36huqNC5ZiEQQn8RPZ4e8agyD7zkUPSCaG3RRF
1pDwsjbQs3w0r11SzF+pc5Tm0/zDYGGwif2OU4KhFh3AgWH6x7b+PgJXmB6X8yN8
JiCnAS8xb/x1S4CWWYeHKDey3J9nQKO1OW2Magp7S5e0BpGCfm7DOKfQmK7g/Ea+
f4NByteDhTKCuC7nARWniCzNYlI3FJ/aRxTn87j7X1scqdkh60QYNC+OUaiQpCgi
6xjAhwxfbmX3cT8QRCB7KkielpKWrhty28pZm+tkwP0iRU+ohmtiFHQm+QFEf6QA
q0wkwAZAoWWDKNaHrO5ZxTaY3zWSRgqc+clAt4A1vBlVfqbgpCao6ZpTcLn31gEt
F6zuX1Gr3yAdpYUGNxIss+pOV961SYB+AMXxYbBrnXPNP1lXMNH23jtstHin2C1E
XQHR7nwInLjMlnO4CZLwxkGY6r7DrivZiW6rIfQcKO263UQIZw4T0Qn3IHwaIp5f
EPOUaG2VHlL+xgwIAAmLwFEgcRWay9jmGeC8c1ZVmSkpMNmGQAfVI//g5S5PpTjv
r0WREot9A/mG3iuf91jdAy09H2DCIGUM27Gdf8t0YtOH9X3FazzLG2iegwHCVD+r
d7R8e8v2en1NzZWhxg0b3GDEP4ent1ZqKtrm5bRqKe3Swl/p1Fr4tT1cJ0dH5meN
H08bMsO5fviKz6qrD4u2r9jUoV2hycRKe+SYnk7dXyN8/EMqMAz+T3p/XmfLHrTT
WG07rNqlpaWzW2eG4/NTFwzBFXWD5CDmrNqfC0Swf7XuxLGX4jHdxS9+vElToLvR
svqTxjduV+NRidudD66pBmz68iMF9Oka2iLOVspLLzAN0waqUo27VCUPOmy0ztc3
927xPyyMyyPHgIGHIJbn5nop7adx9VNBJmbLiqZC8ACylvvx0MejrRK5FnZeRMZL
Tfn+MM2McatS5D/UpIJlregr8ycHH/PsMAeMsu8TohhIKmZuvHPsooRhRlGtuIb9
O3Ap2kpDN+UYy7i3MuPV+V7zhEYqJR2DsO8fkBfQPQVyN3akjovdPqEW+DmBoi/t
l2jSG7jHP+mvhoIvpzXwcTjnM9qE/uW+M9uJ5g8kFaar7gc0kzrj8OmMOvC0NDmH
FJsK0EMxJECW2hnhNVdbPIfNkcKMXjNvzN+X/TUvJwC8Ruurxc/d4+cZfpBW3CUS
eyLPaKQKNrlkvOmrIUa7cW0kKGrXIPv0owWGf1EMqIer732NAiQPOzE137jzfJYp
60wKqTCHoGsEffT5DdZYfM1U+fVZh/N5uUMhxh44+AWJMzO8Xb6d/g9xhQbdHphc
vCuTgOiW9DBK51V5T0BeMk6CN6HreE7yYcTt6WJy+ltVo40Ap/sA3hZHRVigaP3C
4LQqKTCrBdUGCfkKsl1QgsUBZaKeQ7SmZAi1gHcHHgN6YpQ+JQni8+MrhMaUWdgC
zxQOMrc0v3YtAAAL6u1PeAhl8q6V9WyeBfrXIxnnOHt/LIjuztxhWZtXEH9FEicN
k8p260VHz9bnQvqaFfX5+wzd6qOahrR831wUyC6ZdaaaWoBRr0V+/dCFoCmwdxJc
Agc4TVz5i6yYHG9qnaBsq8YFEPa2jAaQGlsTiwN+XnrGVqYN6LpjmmgPb6cssapQ
ngtAN5oqVWPMuVlC6bzlRcIf05LWF0obF9dP+DbE2q96T+dVIN0m/BGLvmJccUbc
HASesZbDoJsxH2QnHNyPCmK3oORQCoikA0fFsGmAr+IbfszLuCwd/4MscwPzLA3w
DyrdMmDcATfKEd88yQgH/jbBOO/rs4rhQTVSv337WfiPqI4rmY9kDYKEOhuf4FXx
2PM8SNzCmUEYlvwS7tm/lPalQ7BW5TBt99uikLO6vbvGkEtWr7IvK6JH0N8k1KWy
1sb+JpF/vRfTefsBXJ6R2by1DND+Qd1UFN/sPqmrzTLsK61BwyjzOMyuoXM/Ts2N
ivUhKPpX8o7UVxq3VYJQiVmi72gsmX4isE7XWfE+GvKOIkNVPs+LW9Ptm9NLe5ji
ok8vfEAXyemH1u+iOdW4C4nySy/gjdz4GrKkNI7n8ndyqFoLXCloq8IGrGCWxUFJ
bdQN93aplNPGD5rtXPce8cOWNFTsku1qAM+h+6dZWo7CXtjN9e0UpinoNV+YZUPI
K6dQ1HzG4fJ3an0wTF6rtz+Mucqwcyvy3F0QqNvZUNQCay/RoprO87acjyxgS7x+
QHrnFNjxFW5iFrry4CFP7zth/LN4ceq/wF2pm9Mbo2CEKJam/4TyRJFKT5G9q64e
XY3yvB3HWze5Zg6PYr/mkr8Wk0kOs0xboweWRTLkjzAp0dXpbYjrekw4lizrFWud
YnecCOZgI/JSdoG2yd58pyfRyg2wdBxfYf36xIRrQS9Ty7TnME6E0QiqUoptJtrt
5k5F8s+3vXTD+ixc3xkFUE6Bshf1B0BL8bS442ukx36MYGNel4ppRo2mcIfBTvz3
/rxT1cvO2UdB5bePtyuMFte0mk5QiTDJ0PkFCOPS2d+uNPuq6T474UoZXqJtayM2
WmnvYbHAVf9orghlTCwMOjHCAHYEfW51BXQIT4V4x8TSgpFaK420ICacDRYclbTZ
/LdJrDmInkHPoc5WRqLSKIJijqXI3YyPMIf8uDktRkLnvtr9yLpWFJiMtXY9VSLC
3LOHCFN5kuWZ2lUbdTwpNq/YIDY9J5MJgPeY8Sac3HjVxolrloLTh38GNOVpi19C
UZBYA0hfIDB4kylQy2YQOH1YMH7c9LyT7hRVF12FBmOz2wMvD6KZwzRFqvl7qqqx
9bkrG8sVMvdV6ttknJj+/9D2Ho4EHaacoX+tE92zsNb/pLaiLjLp6X835Ig/dAfD
/5ry3PEgFO7t9ESrxEN9tF0brQUMTIc/8BAoOMnlAG7WiwlZnKrxC5oRV0yAJowV
spvxYONU+u+wbP/YZgxqvF1ikKHfVoNQDofNg2fui373+i5mmMK/j9r8ejpgODaz
IhWVDP/y1PT2QIs7OIYjd9g1ZekbxXVztAqOHirNq3ShJpfWvwsc9Vxt2Crg6mOk
VUOfsNGQvdkpy+/OJ2uN5+mIWO/qa5e94VkZIDMCHZkK1BM+fnej4GTCGPA+Fd3Q
cOigs24MAtqRsTcB5Du+9t2dkxB2O4YTzaeSx0tNJHau4S5BolMTSuHT7j1g5O3B
uWn5WoLx9HG5nnsvX+rvHa83EjOxU27jzexVxJBAik6OEhd5AYWItkIo94fIqakC
j5SOeA9Urr/wPE5J5zzO6tGiGgLKAEj/cZrGDAHL6X6HicV22NYkyMN9bAZOV2e7
taLZTtzthbayqdFmLlAOc98X8SKkQUjxFSx56ZLSdEmkJF10v5fGqxVU48+bC5Ab
dVa7UTCUmen22oUO7DfemW5XbW89HJBit2UXJPRTvQ6RlkNd2KblZ1MYfPDHeYzb
rEdnTAfcPvzHtRLz7JPmxLhqUALJ3AnodPQxIeryVOBLMN5SmtqLg82f1votN7K6
itZ8Id4lH+IMJrMmnoJ+JfiyUkqW43LAo7K3vbVlDBPGhTQXF1voEIaIG8Ew+k9c
sUecWC3ammAi3YDeeTnDgh14cU4bNBl9ImoHMbyqWrElizu/KYhqGNplkIOZsNmW
e5SlH2+HjG/SLJw3OT8O2ekxrpkDWXFkRXbboolxualY5n5raTLJulzz5+AZmwgO
hGUKVTd4K1L5vD7dbPmG89rfr+X2Uje7a+pYK8LosIHdJcMH418fnx0PBNdUTgx2
6nptlBA2TARnCorM09OXRDU91g2mU2yj/MBrKiytXqN8GEC+ZGUM+5UnyVrMVxNo
LOMRgNOHx+b4fAtCQKOS5AISrfIAhE5XsqNN1HSsIL4r3ddzhCl8Kwfcq9Xj6yBk
3vBr5FMEzGvYYC6PLyKGrwkpYQ2cZzbzWav6NEn5QilNyIGIfjj0H537LoRDMREh
Jm0ItKs0VnJYrr3lXnyMKv5/mZWKH2QlugZGhsfNEzeJgTyukU7bgGq9cijNuZE9
Ln8htjMF2sXOz1Lgagh/jtZPUEXwYrZY/rXUlz0FzRYqgsjIj41HzEAJEuhfk3KL
CKM9V8wGH1t6n1N2IiSOiJzJGsYqJ0MIS+x1vQ23bSrnc5qJaMdRw1/gzyvFay8E
cYW/l/++d3DhMx2ptUe0lEDZwozfX1X/byFAA65WAJMHu4CVNsPUHVvPuBLDjSOq
mxt2azmZLXIboUjXjoHQwq4AePJgixKggpvLFkQTSdozkEuSTBQ3HwfGRbYc8AWg
7oGoibbmQemkX/XRr8D/+y+rSogdnunWfdpllSn3WWGP5kNh0KUIYIQQMPwObwmO
eiffRDz1Upv0zmi4UTwuSLpPEqOA6cHnv4ystWjstA2qKpx5hP+UH+2SGNy3+7f1
dBBlGtdlugeptOIuzlqzbEC+p/8kH08u/XXPVq1Ros2s96+NrogolB1qJckyh4bZ
iu/Pjhj6Z1Dv+GgC47W/d3Jnf/0TzYjWRslMf+vSLZvsALyAzHmGFVI3yUyN2vAL
zO26C5pIRS6IrRDzXLDGGjxx/U6a1DLVBNL23rv/Hu8Wgbu+/ycOVOF9vac09/1e
1hnyleVy1/4uKMY/ZxLRKozLGxF52ug7YUeWHmIMX2lLVZBN7NNaCyvCrw0wg0lF
Wv9qFSfPwAtjYWX8JK3JX69/1KT1n7VOaJxMK8pIZjbcCZli6Va/Kym6voHhHVk6
8ToBrlEoAG8lMJEI875f/X/xG+Pk8KfmIflIo2O15IEuGnG3VApWOVDsNhU28CmM
0WhVtT9sL4ijusFyb1pp79VKe+ltmI77k1liUqZgmtQDxgzedwHuDR7YOBjQtAjn
gty5kbe4Zba+n+nFJV+/K+isBGIN4vmN/6H3tBexvY28JpbKKXFLDHg1SHZcWdbt
UMfaUF5Fvp52EZxEkaqi1AOZmPjVHBZJh+bZzhDVjHtNHBOW7OEHUTv7D6Q8wG6T
Oo37DSShx+l3BBq4a6cYvqORy0GqOo5F1cgBSdQwDIJF4723K0T4JsnIbWGOkyll
6NxqjHayoENJy2NSjvpdxoMI3EBYoqWx3F57xrS4GVAY6exXDELgPV+WaGyRoqWL
eSnW+ek9+egtAZveT6MSGCofsVZ3sXbNGkgA6Sp7UAFs39s46aKrncUMwce4aFU0
DaprHJJpmPMO38q7aCe2VrYYXvsWdOJbbWu08CbANSnAiWAu4PjW+DCM8fhpNwJ/
CHanr/OKf7okrHj7a0AtVU+jq7E9DUm+l/v7K/JgCllwZVULGnXEe/lSibT9oDTV
R/FxH/ZS3Iu+3dBiRkVSZKDIdmqNmtFVWCc2LEil8F0HJ6VoKfk+CCK4DgEcRk5G
yy1DSXkmRxZzGCqsibIOCe76MT3tWlgv677EYUzwQoOwvJMA4czk1CZc5O0rg4m+
vnM752RtG//pfhMU8j2MNzmFRgTh4nPKmZzzkk9LTjRhLz70ihH10rLPk5GGIQAo
WUpHNEZr9cREYUaOYXm9wNqpkAvYNC4to4fCX61szTpmkCIHLnc+SVuwCx/PubwZ
PCP29CB4yfA17K4Xum98iB8ujwnDidW5kwbR3CmLVG1rS5MCYJk4IZt7aBbuEEcq
fdldPwlmZ7kSef4Uq5G8RYscbIMSN6iydK+3xLRlfR56GdEZi77zwdZfPTzwDZng
AhZ82UQMrL5s3w0W63a3jmCNyLuOkkV8vJnojxTp1M1inT73q83Nbg/ihtrmWO8y
qAmy4wRPCU4t9UPV5iwRz8QGC0HyclQDSscHN4y+xoVD05Tqh2CRUn7fXmpoxhsg
zz+rcqEIk3A30tO8gdsztaENPuR68FI2poLqVP8VXr+UHOFyFS7kGU686vexeTRS
gjlP4sYiVrxyuCkFTRQkydiI//DUEdLR8GCR0vX6/xRomyb1sVQqU5M3x004KTzm
w726Y+/uQZvtfP05U3ClInUOrqIzs4dNYY+Ks6lth07cAXPVl+gDAk9XGb76xv/h
lquWo3opLimbEuairuTP/j45Rk7/IXBvTrUVW7dgAvB6sOpxcNxierWi+AbP4keY
GBDFbO8sOaH0lXZtujeBXUFLjdz5VtTzqJhwixDze4XCpuLyRaaYoAeQtS72ydtk
yd8AKHYAdZDar4MsIfTyw02cYMvUqOoHQxH7MmKtx0iiLmuRvno/egl6SsCRqQzD
pgjDaP5FPTFrOiUU3nCLfuRR09FPxua86ZpvsompBpELNIdwy4AoYOGviGW1sfQg
JQRnm2V0KW7JxxNSL6xoWvHU2bfk+32TU9lEWci1P/wBAbchSA1gfUDRK77Q58JU
rxwx+wBGxZ2FuuLEToTAX4ckX91AWFbsKgpl0JBCfg5HNXqMPF80XCornC0PTmmS
2abC+f/h07QhBtPGBZHgTuztbVCcxxFOq6FbpCSZbRjwlXl4ho/MledTiMb/1q1F
SmkmfmqECdcQ6SjEZiatRRgchHmb5dtVtVTNMzCSq7T1yTvG+gKJdh5VWtZkKoAh
FOUsuxxjU0sKPUjSajSz02QGP9Ress3aBH+ecgh747nCYrU/FYAjseMnnaGVRD/Z
acAeRshhOSJITsxZC5sEoCxTeiyG+SYxCS3MegVYKFCMK5KY3tZFRfjMo7UbD/3m
+swUjkI8wyX0uTf08DYzSorl6NeqZcjHtHC+p8fBS+35pkU90GPyeWnzqut9HInD
42gqhp6/soqthwcBbvGN81IE9DuMoAdtnPqmitI6Aj6BZ3GVz+VEIpc+2SYVd2CQ
LfKRqkgUuldNeB3YCLRwqZYeJ3uF461c5d0vruMZz0BEe3kNWDgjTQcaMzNbel/k
hS3uiXC8qDKlW1VK7fWD8F1XnohnBiR0hxW5g68mw45FZA5ruvvkkUtVLTRCmKdP
FIKeFyHnptiEer2PO1EJ5i34aRZ2EbmYMiyNgdvV5Qd3fjR61qWyw2w9IqjVyj2b
+lZQH1cjn5smnHcSGilJ2iVaF8QXCX4j0tD5bTlriLpKb6L/CpGcZ+KD+EP+SEfp
70eCmWep0MiDk5SpdCDNqR/Viok45UHr/SZlEfcGA6Nnp+x2akjh3sgEJvS5xjcU
42wVkicI1LXDx9AY77O/VaHZDuOCcONsLTsx/oralXbmQnlL6MngeIvbIJztr/Zb
xX/vduuDNPqCbwng1KU7Zavve0+ssHWeymzrn7Q78xgQcU83x6ogbmL8M2M+RWFj
0Cvy3rd+dGqj8PNQjdDWdTHPghPcv/KAVWgiEBxZCbDIc55hiIij17BEyL3i6h7S
xLWjPBu4X8p2jIfi2YFVoz60U/AdfXkQDw7J7OMTLb3QgeJAUaDQu+cUkLCc6xvB
QUA7XGokyQ5iY5EmKiLV+0CBCulQI+yy6He4tDU/cgcHUKc/rMiZ6rn1Yyz5e9oA
1WVLEV7QDNSLcaZL2o+JUxtXPCoEnU9FtqgROeKvFJ9MiSr57IIvVIfxk3elDZWK
dK77HTEiyK1vG20Dhp/XxauCdI4LpQx5J54hHCFgXJO03hCwg2TI+m0qSFYaQu/R
kga0jk3uUNPonq69haMg/36ycJAT0A+wCwhxr33cbZgDLEPyi/M1QvH0w7kBL/l5
SAJn5MQcVKI7yw+8pXp/nAgu5y++hKu8FDc12u+iLu1UXpLv53fwFYRhEg1rW6JL
i9paWFSH33U9Nu87D0u7497XyIWvAvcQ5HRxOCA6L3dXp0Zi5nJh/Y9+4YmsP6Ws
7EB72GZnEaPrptkFnx+VvXAa063AqiN30eb+Q4QXvJAOmms5BGSHYh9cP4mCVq2G
JmAx8sgPTebPgKQnYa18TYrN5UvbAnr4/wegAeez3BI/BrzADQvztXrjUkMayYDk
GuVeBd00E88cWBZBMWkA8Evgwx0nT7B3SsJYFSUpA0UknR3zNWj5O1ciFMogCfQt
q6eOWGeQkQu9m5WmRq60REAApyv8OZuCdP9UwewrPwRoI+tpdYtYUwA6Kjh9R8i8
0SnfGAVNT7yp6Ak/zb9ixS+rlw2QvI8egPPDpakSzyS3eR1o5dKwr3AnZD8Dt/IX
IM15HtldHnPeTyctmBxR59Sozmyh4RvSLbGvHJAlhOMFOs9FJz23bG+yqW2L+eHU
a2nvqNemWLQqgXxfwHeg8kTir8hPp0WA5OAzLDl8pMeC008OV1IDox5p8T2POSjH
Muo6F98YL+2u8XTwP82TB+KP3KPB7Rteb8IKdXxfr5200ZzbWCtGGmyoabTRxBMz
1Qq7SoKYssGJU9/SyBFzGpauCUxyrgA2N8+wFoisJ4RpXlUARz+9YjuLAMROImXE
IGIDbgz9M69fK1CxGCF/Cpeo9wOwom1Ywk73f/ilnPdSFYz4UD/cxWxtomS30ao/
vgS71aVWFEjdIAfAEO9nE7JQt1Q2zM9ClGxwEKxpbz2h8tzG4d+ifFDRanZ46k/2
G0PXk1XKErSAWd2JL+2qVRwqi/g+VaWHNFmGDXY24ae3fbChNrNkGFW1tQUbs+C4
rwr7EwAr9QfPrkj3f7T6eYdQWfKa0+4F0/V1rRgkAz5mGoloG6HQNMx6y7vupuR6
bnBrjfC80MVDVm1/PNMovEWQaU62yLniRqcr1BCwP41WH23Tgb2S4/lCRSnidduv
neVnBJ48dlSY0i4AjOmsEfQNYmRkS9eNFeq+ny6+Pg5pAguOP+WdNIMk1Z8+UXag
E7YUS/OHzE0JlbLn/kMV/WjsTqiXY7HGyuYUSyZ/5UroExbCxl/qOgxKUDtzu3oN
7fwade9D6KEp8WTbPehT02HxVSNjp/q2b5RUoPBYyZggi/Zq4MUyBm0OqLMCOvrU
vVSJlIQoLyKJKCrUC22JIplZgah28weNRxF4clrr/HsL+WB8FIZpfL716CPVFcLM
RJ2c/y+iTqEeQu43hGXK9aD/qbvFViuntTOj1ziftjl1Aggt+2JGU2nr5BtDpJe1
KkvlOK5zxckui+E9NywawKojpS69Y1jNM0hkHF2NKkYX43KotToVaiJbTazGRyvi
h5X2tUgspRWaSQ3scrdaOrEj0V7IUW2JUCPeAeEdnnKXEuB9BvcNKpX10HIxF0qb
+lTMuvtqkJfcLrNMLwc0Tu3sIealghyNgUonOPCPJEADaye/svKXA8XpW/YwDdbS
/R2tFr2klxkMfbtYa1fqoriCaKdLIDi51Y6Fsmlv8/5pNCXSdLJDiaXndbkwiI++
q6QsvS2zezFyDdIkJte3QuW63+TYXJzBTmRt+qZ0/CgwzOVN+gCX0V+OoYhsYWu2
ndmC+EaVjRz7GoJRimSVrUbHqhqVklPdWvaDL7jZHY2f2SdBdPZ/SHc9cPTIyeS7
hnVau0ZoQ8Xxn9/GoI8V1Qy6TzO9HDNZz5ZvRuwsKG0pr2N7n2u8CHkd3KxFnHFq
jXQx8XzCT6I9HWPNY8JTHULIckDuC1gzhp1nFI0+WRXDNeGDouqPrWlxpduf1aHK
BmNpfWgRScLY1aNSTJYuLjiZ/Aifvqc2KHvH0WIdDWP0F4cHi1lTPqh+iemPFkXx
VJ+4GIMLuGss8ncQWLjD9Fjc/6l7LzTySfs83YA2bPKyKgGbF8ZFSQN5aaZLI4yC
HSKh63z3yNxDIaw5LbCfynt4OPgBwCl1gAWHLa4KfO+jXhdEtZqCYVlZE1F5ozzc
M03A8BTnjUX60hhbLU+qP3A/E6q6k42p+qYPZIhOqwt6vQ0WZZWZp+ZmClGKAudl
Df1caqXQVcHE3lGgitJj/MCFkmORAXkTYr1a534/TkduYA9LPnsZXuFrsiQesIrp
A6ZOEKcCSB8XdJGoL+J0N4PFNIY5zjK4sAJUg+ynzvOnThpULNw/GP+T4qhCP+xb
cMNGZJrYdQrXdd5Mn9agXaqlsxTmpFrs5iDOWEiEnSZ71yqLTdLjfiAi3beRYpqI
XEJbMpBnf7chTcgyRgC4ur0NXvW8rm/BeE8e8mx4iUzUuzT+ABgGLswBLWEhO6vj
J8+IYZYcbWkgQrf/k4xEhx4srwmy1pkBv/qxX9iPNIcX6Q4u/8KM2EDbVqMjKDx+
i8a4psngNC64qCMOnH8JfViAhlXR6pAl61YZbJsJ6wjEiUfKh77X1gQSGHUcBrQE
Jwu87L6A5gTgk+/JflAuAAHtXsWAqrUqxaYJdszYYxh7HT/9/i5Fa24SvifHV6lT
aGFgrwul0rG4WPIpURoMsIPzbGl6obPhzfvwbUhrLLH/CRVuicb0Yuqsvt83D2ap
9Fv6r6cwk0a2XBHmiNPlyVPlc1beQH7A80yDVazt3Z2ajgsqxeed7P42KrVuUAT4
7J2nDw75bNDtuYRo6vZ1/EW9G6NoLyONIpIo1J5vb4g1y6BtwIeKbYpAAb2W7Qi9
WOTenp9Z1nn5ejvQAH3anC2munstkMKgCi2fv7gtR7KpqYwJ5ZqroLhlYzlDanSx
46ACZXDk17SdkqxDoKxHalUHDORR2I9qtAnaVw1c17EpFu32zoU5kXSNnVVSZvVo
5BcI5Zny4HqJWUcRgKg8MDl0LBqaYJ88P7gft8pOZOmB5k5OIEsiEX323QBAg/T5
9SaYj8R4KAIFoO+i9NyqKc2wd+4b9SBM6+NS2ENq1ZKhOvoB35tL0fv5Ug/tFkWA
8hI6li6wYmV8/E8Lba5VUgscZ5cww8x2IAPDQ1gPhhDGsQ0W0SQSIGG8qYXAfYzW
LME9JKdwr9oV9oiAfmbeQFl2qustlsWOWGVQTARNphBIW2vcjfCAv8OEUl0iAHwZ
yV0AiEZnfI/Rm4wA5jkm6NjAiUN4BrlMT4FskqJlE65uVMWVu8zuJhSpvBWWA0Ll
3hHl9+sEuV5mPP7r51f5HgekCc3kFcIs+vzReJJ9XotBZRNAwu1mgn9Bk5rAD/XH
DMWloKEX33mmGNHIbsumE61R2p/TY+5bRawczlEUKG2Z/y1TCEhi9UmAnyYAIcoB
L55arm4GFKTvdBgJMQcVh3XZcnwV/2bOGAN3zmL6eVpuumBVoYsQ/t5P9tugbZRk
ROX5RKqnYz/YQhHCwiz6PnUnV/hO2EZ24PVTMuVfmpTSHgIoX/fvQySLOZ8H/Uwe
iVQdrBzVZe3ibFryqtehnCiUGy+WYrWmxv76T1lyKfoCXCYl9qzuXcJ4DQNrjFSc
aJdh29mcBmDYtfKPw+bQgnpZSdaRRI2agL+DItzokIqp/G1AhfANcEiejZM4c/QA
eT+oARzaJXdjTP34SwycgErMI/50ShVNPgIyaeFUiFf1LJrS77hEHAFNcdvMTeS3
nYG8OiC+WeaSGAWv4wFkxKwTnsijKPWdMaQ47gc6Zr7wHeufam5rZe0uyzsOocwS
JL7ghvb51eaIxCJjJJEK6+e7q/UjcacsxxgVX9qqi+wPLlmP6/c9YBgKGoOw4XC4
ZDgUwZU329IDdVife/0KlZimJRoDiVBuyX5G52139A5A4nIwJm3b+UkuulxGGfKp
Zbqsel/7K392leTcnUtM8CIJDAZuFV2U0rXF7Rhr8cf+rBWH0TnIwhT+E8w5iiip
Z5gz+aOMpvCDOZrBBWxhSHIVLpoo1fsqBebVcjZxJfrjEai7UAk9S03xtbjS/T/l
OtPQ9zOyt+XjbOnHPF/K/IBXQVLC69EYfEF/KCPe/p5Fvj8Xa6hyFg5lrWGai4hE
S4iW7HjUv6l1f9/+G+dk9aVZppFZYZQx043MPesMXw3Kcm6OJy1a8RXdXx4jhiFn
+sge3xdgrBedsctFqlr2hADl3TzHrcAQoeSnlKzUUM3/MQtb6eo4xeqxoj4FJJsI
x8gEChPDAMh3/yU6nbwi2ehnpyxvqrndYrF4+8+VSz+/Zx400awcNi/TM5xKIMjE
LOaRl5rNaIDbIGUyH0r2nR3kHiWvU9Nk7BE6DFFd1vYfrvJ0dAyy7yhIMGsU2BLD
fUIGP9qaTYp/ShAQMrTh10VLzhEbvd9wC6j2f8hvDINhCdKfWsCWOo1eCHKZzBkl
1LjfeNHgjVKUas5Si1atW62wX9SidERvi1dTHWk/F+MyLFpcqvxMUUMEfV0emdL2
0CJ215bkrx+ngXywROSl+cX51mkZx70oTvDBtlOn3l0jNgNb92O3W3VlH7PeQ/vi
1GxdumPHdmLZax9TdfhEh25UPqzCkNQh3/wG2MCqP3ZAbAVTAPwZmZPoR7VxNr+P
EcrRGZTkT4WnGGJisJB6hImRv8MQCM0JoUiNgY0XJENH4o7iiZOMzxn+m8EYIrcx
vX6Wm3vOzmtPfp1V+vbMNEAm0rGC/tbwtYrItCKeASV0VE4avCOLV99rILXQFg+V
O0r9Jm6U0fa3bUcZDIWAU3IFUxOYm7UWVvzfBY3NGRIXUfgpk9amgHOgBRDUS0AU
UMlWxoWLhdO98GIKPztHkfArDTtR1iUqQsxjxUhUEnejOgliRhwZYtCRe9JyaJ/k
R3aauuQLa1lhMQ+VchC4lspeGflGYvVrTo8z3me9Hhs6MIuxolMK/fSG+NvoHFxT
OJMczQ7T9hPsEbuDiw4x72OQTiIzG6FHl8NZ0SEpM5+NG1Ly7vMoaq1WtusiE35v
3E18qvQ0rOWesgW5FJO0sAbII7GHRZj0yQeZaZqdp4OZLOi8NjXj4ZvnxwZaQ0z7
oMR3rLYGdqelXpClQL//gjZ/6KiwYJ4003D8vtsJf3nNLihUTms1JP23P47Qw4Xu
FSbkJhKVBLvzhcVG9k3iv+CBBX+DJvw4HTbzw5Dq6DB6EROif72Frqc5LcKv56Y4
125/YEFdNLFw8y/QdDI3qwanFi1V9o2d6fE8DPW+8ovgvlaA5FYnjuZKpn9uRn47
otrrwoU6A1oyutHbAxzkPb2mRaCf7X7F8/oTgq9m542XxbTOOn4kSbdEbbJ6Q12e
HIyKnUSmjmi1jZueVRKAMAxQypvGx5df6p4JhqtZsVxYMDh+DiWSuM3EVweXn0gL
JVckODvfOuQPM5sxjcVz9V0pSOUZpBSCl7clOB1dKyJm1zy4joWyYQrJBx1qztfe
BwGatbho0cPXvPsbTtPv5dezZId4WtVxgrIrgqWCsTX16w6kokd/HAfxvh8/6TRR
0MGlyP2knwrNyh4U8yuewjPYojv9LkMPzMsXkVBzsLsqE/UtFvVPLB4QqhajgBLG
mdoGAP5m6A3UjensjT+e2Lq0T7ymMdl6SpO8LUkNk9Uhoi9CIvgexGN9iFPaiFUU
30ozaaWWodaVZDMkx1dnNvE4i3ZOU01v/8tAh88S3jItuln7z2tcwtLqir6720uw
ExlnaGLQACK0tSkEPbk7QixtRHeiDueQfUzFls3qlKq+TYigfLpOyinK5yL99o4o
IyA1YlOBM7tm6utgumkV3ISyCs7x7dN02cwpo/+SHhiLJwSZA6jGrqK80NevnKFc
nLvGvSqBHbPU+Cny8qLLVI98ZjjRH6QAvP0JotZCmfkHS1RYHAycP8OjivJLL+lj
O1QoOg/mlGdJ2mlj4MX6IaU2UPM9vPn1HrPjQFNxiJ9pHfPq4PDk0xzkplNqhwXJ
T6C695ZOq3Htdza4SePERKIy8z0bEwgzAk5ZJZlSyrSvf0FU+CXqcg3MGrxNczhe
h9VkGvLXn4VgWpy/50Ap1lTois1G2vBg45M4WWRkxlHYnm7RxjK0EuQSKdgb7BrI
AnYaWLcxa3hZ0MY7lwadIfKHJ+1YAEAX7nYwh2p4+2GRIaC/YNn4fIrdXF/zycac
Xil+RAa4rmDaHm76QAa7P1GEcDWNDxwpY8nl7IpzzWpo4lbwDQ+24zLFbPDuJQPf
kL5+Ll9Q7RuEp6ffVXTb6NuSkXlQyvr97aSmpWq0ZqFr2uOIufCi7fYYhPCniBYu
5iuogDyx/FqrZrp6OoGbaPBM4Zdr+TMrsxn9FhOOJRBXO6N9czF5KMBe6QihVa/p
pVxZWFGrpB/T9Z86bg4+9VWSzjxrSMScK9INXaakCIdrmt7ws3T1IkkI6F6YWIqD
EuSwYPMwGMHorUskMpU38dZ6U5ZlvQTLM9OqiiF1qz3zRPP9Vn9kDW1Pfzwl0/Vw
xy+hrJt3EwETZhVd/nBVIwOPYZLDO+YF1bPjijE5qENzS7LfkE1VrPT0rdun675F
allNIjCtRCKW0Lf2pQGvKvUAyG0GleP1Xn5vKEAHOWLvoL0SOxO6cIjlrXrYvtuq
uRqld0yvpzhWqPTM1npVTDk3TSImSNIJyO7r/AWpKe0kTrEanl9mZjUBrl2uMER8
/gRVDvbAsB9WFEEwAhqW5/Z+vNskv6XdpKjsj2s/KopM4nLjeZ2UQ9FlXg7/vhy9
vQpG+Wmw0RKvxsxvEi1FgbPXwWwQg2ba/I+8MThs7bszxWY0TqM1gk7Obp4T/Z9W
vYui3rVXenRxGJSmko7oxfiCgqX0UX6G7tu6adA2eJMzrvhd5xbkQzETPJqZNd/s
Swk+4dejL75dYxZKfAVmBKhVuUq8KXUcVmvs3J9AWD879mvffq8lNPtIP7qtQeIh
m5/8QCleQhj+AvbY1aF89L9LhVM9FJlR69uTV53DELV21voi9Wci4Q1vtVzNc+kf
ggtVlShsBnD4WxD7FlM+fHT9/3TsjbGZzoTKzEnibGoDAbeWqLXc7P1769z0lJRB
zeUgqXOfQEIUXY2ZpSBvLHlSCBgRHILiR39blNM3eZr7f5EKP+Ob6sbAJWYSzcge
X7r2aWUBRCqgY1aLIlcdIvErGh2Z/fJss+OqUFTOsAkL9TJpatHW9EIASJS7iifJ
o5GzA0+daXkpxLDqJMG+h/sWvwM8NmiRIl/GkfkcIG362kVbMsllMn92hDRrDdf/
qwKNhigd7hFMeF9qhZbg/b0/UFI2PIW9QL2D6gY/tGSgqHrWqUibKAR0LUUcrKDE
36y2XVDtYnrwQB3sMyTF1qGUXzRnP51J0xVnVlYJjD0wPS/qs+bcHq85w8wAfAF4
MtOnUmwX3jkKz0e2VZ7Nz/OZMrvuWe+EltMBbMnWguuhDkmdZo2WlcjkzNv4tmX/
FP4kaRV96Dag7w7KZXpalM53Tw0z/8k1/BrZQ1yzRwIcIl9lppAsaMRCkWHscu4K
0eurYEFLKRPAMmJEFLQLOFXnmkbX05poXnHi1OpbC04s2kNOhFBKypX1ahNLdE6q
S1Q0SmJqQwoOscQGRjwGzImmO7lvUec2Dn3iIHJsJrIWFd20lymO4Lw6sDnv/U9e
822Eo2GcZcHpauVGUPGgSUhH6+MkoiCB22uu1x7ppBptTPs4iQmGuWaUrK7cKg9H
2/+JJZ/Wktg4OCkC8TuIJXo60v5CyD948gaRYVTIYtCl1OSs31/L8tZQ/610/1oN
3FphKB+reFZeEhikw3Pj2GARSBwW5chrj9OmC3IUQ9b3wBfeOPJcaJyHpc+vwsQL
8IRqLyAplcBcpXDHWQAIv63BHQm+EgAti5DEsiOX+kdQQebu0WgeNF7vqahAM4S3
TMN1tukx+nSENCLl42QRg5C6KsH6JpTVPqEnqYHlwpCQQw9OiXOg571cILIyV2F7
ZA0/AHIDTRW1NuWC9zt4Y0bTne0m56gUzIWIhH8J21dcpj8aCWuk4pvTKo6adAAt
JaxzMSpx/Qo7G9/4cVYr4KDcY3KWWO87623WLVGrvADdURIDRTJ1IV5zBN7Tivru
Ib2xHf0uwvNOdtQzYTFJGpY3gDxcpXiqVVW5fFdmX66zcHVazFgVEMLaz6qby7Zx
uBEyWVlZb4wzLswIVJ5egjUdKh3oHoO53SRXMcnyWZzS2oN04eMsNw/xw0R328Sc
BYh5mQJe7R5VCjZYbwigbBkN4FDKB/fH/Vt4qdpk4fHBZdLsVLuF4L8uIiDZ9LkM
RcbiUPlpZZGyyZ05myKdR+WV2yK/vrsNpAcRXkyujHqhP95qyddDb/JmdDz5/+l2
CMsIes4DTND22soECJRNgyCTwh7x/K9pJzkEGsUSuD7Rz5nDBKrVsLgoS/HKl/HT
c2duHAwjJtoshq3KkPFwCw5tzy5wA2syTbpauJV3324mY0+1iC+4IS/Z4DdTc47L
b/Py7rafOnAcoDxwnx+DSqT6YY2wo9qfyfeQfvA7h4VNrmYfmCytn6CKqzs2hnKD
EnTuVkt+ezEo6nYAIVO/22yDnvhlSMa8dhpOjdmn6KPhi8wt6DBsso17z4yJCpzM
crqEy/dNI4bDnKpugkRH1F8ei9WT5GaRdfcOKf6DNv05d14wJHQg+vj/K06PpgQh
LDb7Mnb/AcJifvPA/VnF9gmTOyAC29ik1Ybmr4Q9BtqqvrWukxKwcAbNEAznLJq+
BBw2snm4tpdwwyekykftU0XHFCKCOtvw8Q8PWjN7/uMz3/HmfhfPs3JWY6YbJxX8
l7Gf78J6L8ctId2BfQ0Zrj99WPVewOIq/+2VfNeFvAMDBmifTO+iV4BsGkkFpOMq
4DhBSCJ9fZA2VVd/Lt+9WKoFzWfz2/NBhy5tRf9KvTaxXCezLiwSsp9zjMqwT53E
DnSEyb3pjr1+fxrUMtaxEN16UttHpxwf+eaHqlt/UGY4pQAiuXXMXK3suxP0Pc6N
xETA0MnZutYvMjk55qWjjnuQsL9UYI8hphzlu1CYaSDUt5XA1Hmo68h7WHD3wQB0
ERf+0k5v9wNwteRTTiLWDDfWRT+RmsM+uu5KLXjx1ljc8ub+I/khHjZSZD+dwaK8
NvMm3IzG0+d0D0Q2Na5SbHlcwL3kIAodFKnhfl75e1+vqXRahtkmJx1FEMl6L6lO
CJmcBhMZP+L/Aye9qFM6Q+lOciJlvNnbgoO3gAs13z1jVfOkIxpuIue6G4CLJ2eG
2UuWeKSHaLRNo1/ilXV5jhKTupXNlsCpBtHt6J6dcFk=
`pragma protect end_protected
