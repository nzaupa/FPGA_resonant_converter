// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 15:05:46 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
abzu3JqEydHy7SH9h/EBVeEjWsLDLRHf5EK3JyZhH+3l2X9Ap05DhyW72n3atxcZ
ackRz5w5iqt83NZEgNLjZiq+z+UZnDJlFjiV3UbJYl9kX9dauIo96mHX54vjrmFE
TvUrjjS7kCf3pJoojh9PRS8SfFnT28bmdQ5+uS9BamA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17360)
t5TzmFviZDCY1EC0cU1YWG8Oqu5Qoo7xOwTDsdc+vayU9GScA+BpUx8MuSUPsA6U
GbKmbEjgiArFu8nXpEn0/+NETA/fKcWnecTJJZvw5zJiUxRpubB044sZ3PUfM4OH
edVPLwHDm9zpUqxG9WNfkOmQvUSG1zgBXlwS7jF5rZxA/+F08+RxzWCISIFGzo1C
s1mzu2IbE0nMA5QvkoCsFbosu8wa7zOkjjVIsDNBsHQXMt0h9k9Pb7dlQdRAnIGK
M60QhERrL8+6byEMTbtX2OLyN7D/Bu+eU7btxhZ/+z/VI8LRbRIALZVJL6M9zvwd
QmJrhl7ERLMfbFKY69w79/xpOTso7niwWHf4ExCUhgaGMy00OysofK4QBx95dMe3
ZwXGnpO7nUjUZtZEMcbujNPy10r+vcvY6dBvNS2qvoipnB4+9AhqC78ggEf5LVe8
OODQrQUKKEAadQDvAhHljeR+XtAVazvXQCyfIfVhgppn1zyoSTM1jbDjRMnIhRsY
DD3wc5magrUu+UrXp0ve3MvQnUfZsDeoG4Io38qYX7g4IIZdozeuhEik2MW5TojK
TkvDypLQ1gFAm3GjmgX2siqQMKEvV8ydP5UeCTFgwqbQIE0dXtjlfCJ8cLXHjf0Q
bxWeFLX5R0BlG27mIVtrVQi2UBNbGqTjyv4lQt0E0dCJqxn+dvTWt2LAAtzAvqDb
9iVWVOWGg6JY617Aq8CL+TvKhIMVe+gShmWky3E1pyX07TBeEgPiTMF34c+bqeGk
ikGEATZdDQ+Osz1he71k+Nbk+Um4Lr8Mw7CnL3Kq5NeZz3N5g+Fv0A/or0LXkCbs
BnqWs2N2OFRZihiARet0LRw92urJx4R6iV00NNog+MhOy36KyNoHdzbIDOKRpN2/
XL4CpeM5sprDTs1PFqRty4rVo5+ChmpanU6NN/cE7WIxh5TB6fNq/Cl9hclzO8Wj
73rCBuCScKyq8oegzM2TZCysoODEdvrKEt2xhBvnuanI7nI3h5T9nt6yu7xYJGYa
0uMFeqGT2BVi0lW/uv+oU74jxyyqJRQOC2X2/bFs4U1sAP/rBNOAiebC7mQOK6bb
k7AkM0e6xnmpg4/4B6knYCjDpO5JQ60/tDCh6pVXcxhRoNTq+kWK4xoS+Az0GLH/
DZTIoN6qHts/jI/4/lLezwEtktbQAqUUS9F+QWWq8ehkcfmcOT69jHbDQdwmxS4+
uCuVkvz16B6Qo/CGWQ0yXN4Zx/GjNh3eKVEkrnbQdLe4zMtMydejwcGi1+jpIWkR
oUQdm5vxwKKfJML0/++w6I3+kqDBvJa9NYEaLSAF7qT3jWO1BSalvUeIGCfjzcSt
Igg+lNdkoN0MJufsd2xFLPSsf/vi9NV0ZMubOZZbcQNwz4w1rtoJ3etzker26Jsx
hKsVtp2fDLI+4zZ4SzBxF3mVURTl3FvQeXv7ehSQy/dvkIcuccdZb3tM6XaPPpdN
JL5EaPrnFd8xcaQS0AKQmwivGuYvHSHxaNDwGSV6NcKI5WAmWSRwAl2lsy2Pq59w
9nF3+Wg4xfCvuX+61gDrXA4yiQVORvA3j1iXcvD5EGWcNr0u0YLeNWvxUhx4I0YM
Hsm34Fef5EvUAqHkeD9Eur8Gf8r1KHyYiVB07eeWAIBttYXsr48FBi5KLbvB+l2h
NohxYLv4Y+Pp7ueXW9TaBn1jkGitLHsnlV/b8JZ3WSOVpOpLexUhaf7VdwhVSIM+
R+7vnJSbKEq2blENZqiIOXq5Wp1X4YKBLS298U5+q2EIagMb6JJMV7/jWw0l7M4V
uHTg04mvadqEFDusvXxr+/LFX3KA3xCQOWMSl/2/vq2z2g2SMEpqVbSqkYbjUsIg
Kw3/sTTDA9f1No1IkSOgZykvgOchXCWNQTkBtObjqrRVZpv+ibRgL9ZT25MWoSTr
YEVD9M48DqZ6Wa/I9E/aaYP3yMOrwFD/cfP5tiOKEI48oVLUuZfPj0XVuo/xCcDo
wY2pW37Q3Kq9ln7cF98f1Ltf139lrAOdSrPzNAM0rpPktrrAL4U6yRwmHwtm5xNY
7OtuIhbLsbxU+b5XUBIcUF63qoQP2ctWxAoaa+iQwVewQ+My9p+pdgKTwOLpPuBv
x2f1cRb+lkmgZrBMwmu+T+dU+92n1zJ4gUgQgj81CZNokzj/+CzuR+w20JN1lWzq
DRX8o1Cs/JycVCFRbH4JAZ0IomKpBWDcjxZTWCLCZD7wXrZzM/nPItW/BEoioHo1
9vR+hT5x81X/sPw1WioqRjwb5mXEx4HORED4Mqyxg38IDA/Y2hnZ8WO7MnbXcA3F
6J4/L45uuGLIjZLVC552R37Js+EySmm/LImnu8CMRZhczePISw0nJ6O4KSEbdu78
FV8DyjOsVNG7pgnDLTY9qywTQgf8klxtwj8aVCiNYltzdODefgQ9PT/k6lwlrPrk
yEpRtSJ3+U8BKwiMxLrtfpxl8STMcYaoH2jRfJGOE2rKEqSMIHRiSDOEhH5eqGLb
8VdJJUb4UtczGwt3L4ZFNr1Ind93m0IAAYJCoY3e1nHT262bxut8vnsFNEs/g4QT
1nuM+76WI08yWfxvVNlzM3Pf9sNZFIljDYBeM00qq/GM2V6eOrdmvhCbZKDOXWvS
6UD73QuseUWfmdz2VLpk+9ObpKylWR2lVMFOHWu43Ir3jEVScaURujPQxqa7lvLM
q7JcQTY8PMpMxlGlHctBL1R+6C1lf7N4tFPoqyTJELl8rZk6cAR/278nrPq1CSHX
xBeYyXzrMWLq1JhmY18e2s9cw+0zonDqlZiGUkmSqNwny45sUUIwvKLwVsr9+ww0
NIf19vl14zoaZlhbBK9mR2kgTVAHN11SwYMccDUJnsZIYWDZW+7OL/kjp/6vNbFQ
7ML8IahrAbeo3I3V7Lb0wscdnlxX7xAFdXXK1rWr8PdaPCFeBYlKmU+VChoa7YIr
PLTgMSpyMnxu8xLemAgQDHDXDI5i8VDhMVeFNYcll6e4B84xevJcBHpMnIboS5+Q
Hn1CQV2PoK0hvm404IL7lNzZ+nDkN9PnkQIEqW6b2EqdSn9xCL1vOvBOqDagzpGL
ozhWYjTfYc8J5t6/yH9azN5NXmGU+VQ3cHGeyvB3bC8ymTgReacEdecbv74+SiRw
5GtypL1qRDh0o7TOE9tjpAXEh0OY+Qn4pq2llWea+TqXZDEqi63lEQ5j3W11xy6H
66b5497W9GNnSTrvzl0oH+ifEYj5QdMbNQmgpF9txN1Wv9tNgLLVe7iNH6iOxQMP
HrOPABwrCxQTfzVFSS7XzLkY7JwfbzzMhBSqhvLxOJZZyT+ZFx/BTzLqfNBgvYp+
PrQ8p5QoKIzZckIu0pN83ULJRSOGrcpySTxU08Rt1LNyRfqGc27B3gkful0kF527
vyvBeJUkT3Rdnr9S6rEqP5eqqnKp6Vyjpy45381/1qHzK+3Dq3i6r6+llnAqH41L
znpnERH/Y4xKu+UMbwjWfeTG1x7Chdc7hIu08cn2UJKGpFH0C3HIb7gE5gXkvq17
IJz4CwsfngLejZpWyCunDcbMbAKHWqJlvWDIjM4NWyqXypVeEsg/GEvRxq1kgO0N
e7NMFi1mfT2reI6foXJRMme7EIAtsF2c+kMi1iBbXt1atuhaO3a0lE1sFjrJuCoB
o+FrrAmJ1EMUqLwKJ96ZHHVg4WnWOnWQV582C49Y1TvkshC4LVpvXfoO1jphojJ4
cC8hNu1s1s5cqI7Xmt6ZweKFqpYnSrZQCR07F0SYduMAma1ZLEnA/Q/OB66R2mxY
u0+eByGkuM52/lq8wlkHVF3sDrG7nRlnNWbI0HKnj30tDa3scmV2157UCGFPkSBH
/SgMeuNdM+Nt8aB6A4z6H+Q8s9GumQ+AwGEhbK9EiPeklcklC1wcHe1QMUlr8NBz
dJoq7QE379vlq1NvtcnVW96cOxzRFX/7RW3ym4PLDmetQeHX2bO2uH7nYQXjZAAp
qFwd5JLmZXZVGDFL3cnRbp6zH28LJwcrum6BVJITKQrzEB7cxfq6hb0P+046/Efu
JD8S31SB6CohH+RwkGv7NlfO21UmuE3qnlPYhXQdOfxC5mj6l3Bvr8SMQ+qQtIZ+
zsJ5NW+7/TsBLrZLpeF1g2FLBKmNSLAkpW3RykQX6ODOHGnhrLktqPtY5HazCYiT
lJL3dBuiLucKmGQXjSu4Up2Fy6qFZcC/1RrJsVe0Mjre7Ni9ly0mAC3uOLUtE7y2
d5A1FcH7WJOCUwQoomEEXMjGR9QJXU6rgKnoYi09uN8a3GXTzKHTckqLF0vRZExd
O6uxsW0aLzODOPdIhKSW/kOeXDS9vuiLgpQDZkp9MDEuNr9z92eUY455LDsoV+05
X2gjI6ZZ+Z4mFWQJXZ2Boy1+TAbldXCNYo2B7MQXrpn8rx6GYvtCWJXoOR9fSAql
ZkWj0Amh8o2XTXcYFqa8ikdH2ao6Y2bJpWf5kVVH/BM8zIdOqcHVaWuDiiJKP9CV
uVrZZGBlcvZNt74urQIlJvQUZwknnHwU+2HxeOyiF8sQS5IHMwrhbc4S3gNLFr0X
Fk54s2j4AaTaza6Iy5Uks2FpP4GhOy1sqexIiYJk33hjjdlDUnfsYH/EZnaAIGYD
1Zt97qTAYKlKir9wRTj4nf+7YXbqpDgxOY84iru10b/7D7WVSbl1Nr6gkZFSNt2q
xSDYIbCku82OFNoxsmzGjnCP7aBEZWY7Dc9MzoFYKC4VHHSidgDwXAcpU9zjaNmE
DPFF17GKPchbc4+GPA54/V5dUvF1qTNPJfjSqOdGyPjiUisl2yYniRw6GPwePVPx
PsrlgcZv7b4hiR6XwZSrUzal6GFEXwMbdXbfCezEZSbPSZEOuwHozs865ot5RnLH
ggHUI+84eXNm1JQQ8VhkIF5Jau82Rr9cZEDRjVmzUi4jSX5eodA7QSdkGb76dhCO
RTI6rJLLwEvSvYrGpY6EYwwIzwJX6jyL67cme0+6YmEigzcGs3jXWnTaoHBUhFBv
Bb7mcsDOHxP8iK8upIG6Wt0DzM7mkXwHj9+4EZ+pSDS3bWv+YnKcVIC14g0peKx8
lInaBHEqSqv4lfNNJdzwOEqv39S0+6SA2sfogVM5G8yznAmdayO9Et3Hxtxcpc3R
I70hVfarimg9NSDjzARyRj7OGWrCyk035QtVWShTzN270rxLt4fYkfwBbaOx+9KE
tDzpiC4uSuIyazDTbFqKOHD0QOiN5zDySnNjXRdJhY+HLvfns4h2Q9H0pJmNNnkw
Wo+9Fs54AUxROtQbN5P95gnU3Q0ouIkOWt5k7PHbubyRQwHhvwQvcAxzYaxSxiIG
8YVy6hd6Mg3eifW7vNINhqZjPULrGPxIy36b8EDpoS7kySPm3tNGhNeqJcWcJePt
Rw9D5zMsNr7D8WZlR+OxU2xCuNb99r5H0wcwTMwFfz7lHFygJna2fgTBj84BkMZf
N69k+n/5qSW/5d6r5jgBF6ilDmS3iFoL1XAYwpBgOAP9XjvsDmFxIu2T6ag04MHV
yok9PAQ4aoaLwpKx1hqMAPm1SW2HcylksjK5iimztNB1LAGHc1/1VV6gnGpLXfk9
NVl+yEs9bLRpFNn4P/ZeuQMa23i246PKONcELlQKVEi2TstsNdYKtMd37WIuFok7
hWWv5V6Ki18JA1sVWo1RAVBCvylanFxZyl31vGG6kQVksSS9gpITFNn9Qwduuq2T
cHHOvtidbYFdQD7d7JnntTQDIneMcHuo4nlQZvDc4s+u7toWBbLIdGYavqal6kvb
iC7ZBrAvgvCcj9gaqvJPgNIVxTXMoCzVSsLul4BpqG96bTnrGm+zuZy8NzKdFdan
y4ierPLbtjHDSFZJFIHXn9fBBhEHTi1H7oSICXQvRRbifSs1nWKocUFcPKPaMfak
YQGu9m8ACr8xoAjPtM8srZsdu0XFjVxpTtphCXDIk8DRp9l93hMYfCtGw4j9Odjk
J6n5CoFpFcgUnWg6nvZMR5HW1dFpcLd1AN6lxvmribYsuGaqz1k6ZiA/Er7UE7th
mfh1k/n+1XKrL2M6aHSefbdAezEXXlezgUFpPQGlfCBSXu78Dzi899+px7YnKpQw
1f2DIQVYZQ86/LAu+JN3v7BaoDyUUdHL598K+KK+2ZkEVQg3UYTKPgzxHPFiaaOE
kWq+nWjV/aouWK1xfjOBNimcPS8QOPs6c7ckfQT/qGkzNkm21fVYoVxKPVnRUgoY
kpN+s7ENPn3rCMbxuIZV09h7Y3jD50OXy+4Ws+/ZhwlqdKrxttB4fBJUDyoznDCs
G41+9yeA/7doAdQxwiGJy5t94SbtGq1UerplxgJTwa5F7El57rOSeUyLDC8TBKIA
KJGMhSEmugqj6yW2hinqMEmuPDrQuhCCk0IHhD59O/6ps+bsmVYdLpkKfaqmWSNu
QTpNAZMkYMm+B9NvbAW+85e9lf3X7I4xRwDtK3C2KoXXvdijwMzZ1ZWNsustkdu+
oNPCmSqnikwyLJ07it80ptGmVc8iAqffJ8/DYUVlVJkI21X8KsynyFZS4hE1DoKC
HsqjkY0CaPMEev2Zi56Pds8oL5R6N4PXfOHxnF76++gWnHegpU/KoUwmonoSJIyJ
fp5/NeG38Ko0qnaZ4u4ydYHh2K95anwJ+rNstw06fib55w0dPQJhOTHz6hXq86O7
ws+bI99de0l022XtWlp6FkzCbXSo6ynTkCio+HA74u0NDM5tUffcsfwTBVwzz86z
uA9eu9/s3eVKzsZB9+UwGQ1yEUNmdkdgbH63koCeie8zOeG3QpZ7lTEVLFlOVSR1
X+ZuMWvUUCKndMnnqKjWi+2H4gM4v4PCwerVQAUincC4VEIBml9Dmw/5aaKznx3I
VUL6nzltoJSy/KSlaWCu5L3Y1EtAfoThQuFUDjh3CXBaVf1DxD3mW8y5Bf3psZOK
XFaX+Q9JRTvTZ7TysReaYa2/ggkb5ugGrDYM/b8y/WDZG83qtqGc9NdYt+HbQPxn
VSMClia3LX3c6H88a8Hh+sz30AIjbKNtkvAHGB6I9H9DBzQKPKXxPnX3oD96SXLk
P5O83RX7EUquRNSLG76wpVVEeOp3AxTTA5DoH25D2ZkMYXHvNtaZJq9ee0+1uH9U
vu/tmVqTXRwLEIKIDD+fL+y91r/0pFe/rQt/7f3fY1iLw5kgRmB+/DZPbDH9Ddls
pdtS3exRHzF4RCQE4XshpVHMos3fhNnkvQfB5ocirbpjUQ5K+LLW0si/poyEeva5
oGGgxRZCZ0cj9PLiCUrHG/4kE+0QijA0ROdFtjECihuUrDn7YGrynjhxELD5UWWd
knJEs0tyuxL+4BjUKD4S8lOxqs8FMcdeBokzS9bMbxiKpBxIO1Igd+TdZ+7FfQkA
hx+9Du8NpuYvb5d2ybrS0zWbIpyTPxNnyZapeJD/aIwlFKs2tKU+2ikSh06vo6Cp
SXiXBzNLMG2p3oPFpCBlfrWGTtbQ8SgMvo3/c8aoRTABo1Aebt+5r+971fIXedMj
o7FCTnX7OEqR+co2YXjBOeP1BAJYonJZLaE8pczOnhJ6L7wZ9YwMWtfw2sbBBsq3
OfGrMXsnEqDOHApTL3P0mqYsAlk20Ubpm+hgXqoBPCba3XTtvM58zygkkQyUxuJa
BUCmNpwj9W6Gk/Ehz9X7lfW41vnUKbCas8Fyr+w8uCDqeBjHyUNrGKc3+ERfTEFE
ZpdXHQZEw6nzoQSp1lHzcf15NWi1n6QTq76s8YjVEwPndTXylkx0AONlqVJmNt7x
mfP6YZlqj/J0/ORonprKP4VsLy8nVEfzWyNArPnSpswdpMqQx1XHc1vyBBE3rqXH
6phSAvKB3VwCcku26CIgNEFe3qcmxX4buwSzSZngCc5UEKgoH6a9Q+gbWR/QPGgz
skyw/DzULKSRasHJDTSKdH/XVc9KRaIiG8ODBa3H0+BZdTpu1RGDXVtEBTgqHyRt
uNUH3H96r0rj9Irm7ynyT9LbgycAxDsRBU/cuiC7Jlng0IK0x7cegstQOvqldjxu
09NYu3QYBVjm8yLr3KwpHYbbt96gLiWQkujnEvmGFi4W9h033ixlh+HSIKgONqPR
gCOub/bWwyIfJCnen9mzhc5EhGoynVtW5eA45T63aXuPQRG/YnSbMlkGpkjs94CF
8kprntDf23NOOeZkNmgKV3ch03tdigZk1kbz5g9L0kbdd+Sos62mWuk+sv54SHVr
RV36kTzyrZc9B5+cnqAnE8x0kizisxBsIjizhHOh44ju3zxevkUiFMqdEgIvMXDd
Fqnu14e4eM4KPIMAC0K1V2XiM5MH6k/ezBFE9RPMc5UvXR25GMr0LCkJTAzuR38f
Mf1J7elcFpVduaiAHPbSE4DQB4wglpfmPMFpcjW8H3BpgO1mS3uas3c+JV1ZCnyK
hVYDMGfKi0XgXP5O6d2SBS33skT1UMP8PMCBaNHup11Epxmwp8HqT/Q7c0wSN7eN
b+X+10kqChAmjOJltU9Y63sQgW5suLiWNcsyhKqDvegm9WCc99KzBj+/RDcziwSa
qbdy5OGs/gTK4tx7livrS3909g2GpDRlCFIapKtAxq/uN3QxflL2XQG3Y6fKdXye
6tiZmaHyc8ZMX2mMI28yaVkatzTbDntzTx0pA7VP/Oz+eccG5TOY2b/6e5LMd2iF
3dig0LConVIU68GhsnJOQVtPzOFz0Gosyot8/6cWKZaECn4YxC270V8aP8Y3wd69
Wx7Wjz/tqPSHbLLT8r4yJR7dlee50rm9/vx9H5tJrtJpw0mApDn6WMT8Trpr2j/M
QA5D8jFOMHDcXw4HFS2WjW1gH4j/uD1Q7NXZbcYMM4WsYgBBibQaokpUyYm1CBsl
Rk+TCU2B5JRbsc9vah3A8bj+FE9Jl4LAsMdGPAhSR3VQ8rWBJdR9huSlOwPVzMan
XUblYlqnMKhGqrpCB4ZnImUNg3H18f1/5ZRlrf+rdPXp0k8ofthlIYfRr8RqYgbo
IuECo8Rbun0Pvx6Lk6ObbljyiKP47pzFxVyNWS25gqhbUGvttiXSuht5n6bNqR/U
JPgDmPym3dnqCO848hptjGbyCIXGHeyD+cIm+UTBymjjT9DUCxfzY8DhCsf42EWc
ShF+gCQNG+2rISUv+bavSWjiQNRLCHpco4+fPgL11FszPX1Jg8L//7/Huo2u/EdH
SF23WDHdadh8qIscm+BN3wGCf9Bk8iwt/pHcLlDybtzMO01mI5RsVTwx4bluvO42
GGELb0cQboUuhHHVO8ItAfjkTnAhL4e62Y8Ol+FUbiA4bUlJQKPyO1Oe1gAOSisc
JRii7lgbaYxFom5hyIhKtiIgsYMJ1r+jKmvMh/OUdhFRB8OzzhjpwNSxA6cuosKX
M+8YjlBZSAySYwdYavP1B47pZi03X2Tr8pgeQt4Ejd2hrWZDXzpzMAplk+/I4dBu
EU0Fw0Xe36yExybL4ZgDlYMwbQP5GGhiohEANlcCPSy2YmKp45EWmNrxNK0oCSgI
U4fxQoeC4WT1C+ixSYvmtkmOqQB3kXID9xFa0fOER8J6P5+2IOJHbTQM6fb0o1gZ
k7wOT++DMlPXo3vJ/mVQyQ2AhU2d5w3R0znbIdzRMQduwJciCe9hY/1XgLVB1Kok
Q+gn2HF5xWQ81Ww8tswn/7gqGjbOIFHJE9NePemNizqkgyfx7oqaMRo9h0oEssE4
LO9Xpyb5Ccl9wINTfmKdbxrmtiu61Kq5Nq/HlzRXINi2Fzg5WuDlnX1WSBPAaILw
CrwL+oKfCrIWfjKHx15ldxoEdJLUim6gl1BZoMUr9gQUsE4zLLVVIRx9VPNwVvB8
YBRXY6fGp5JgkU6KDiGLYEodrh+W+YodnhT4pOEODKBZtRwFN08zhkyV0oLrBdaE
rER8yEF/sLmA7kjmVQqKPhhTDlB7fyZTyyKH6Q3CV6ZUBdJ0t8aq/acb6JZZxkH3
p8xfX9AcnZ4fUS/FQC/s+YZnOUWrDTIbkQf7qjz72gaAApibbf39SLsrjiXc15gY
lTtzNpBZR3XtOC/pz8YoeMU77Nchm4I7HML9wbqLiITkolXXkM//QWWBAublp/Ud
4t54jvvzb+EAGuxyDtwEhxRzyC3aZBH7tw2VQbF6jc4VFz0jvIAJ+yGxJxxy1yXv
9sOirYSzbw4xEyadUg9n664QP0lHv4eHI+akOCcGIFVEfquvA1q5rcYsUmM79Mvd
9DCMrwSYToxo3WZbIE8pkKBWsBVSAJz+weJpmGbqt7EmSkyDbmGwHtr6umRn4fRz
ww6+GNvpAO8nbMZ7KTau+YPBXHuqtE5HUMr62DUlF81PZscZqvcIL9A96QxAkBgh
kMRiwb7Png4ybJCRcV6aQi79aU/hbJAEJ9BPQngm7F1rPU5hDt8P3vsJrPLWqlIt
8XZUDV6t5yu/XWEzOXo9yBuzXzf8PWzba8pWUeKg5a2ycXlddPrDeMYCXoBQSw2k
twoqkUZrrmQY6K6lzvtD2e40ztV2YWXmXhLwLr3VptUE+xMQz9NsHKCqN/XJanlI
P5c9KMliIWJo/kRpUSiO5QRhsLaGk8euqsWUVeiL++GqWSqlVXc3bwgKTgtQVeJM
CpngeCFd/W4rptnHbfVSMSf0jzdMi2aihG92iEwn+p53xejlgtyKnnmqvfgdTvkg
hGRpvgmEky2XbJ9v71D7Uu1DZZLDe0fLzNjBDcYMS0VqJG8keSTowA09+vQYBCoO
OCLbexcf7wB4PMpLzDxiwJjYSDFO9BGAN4MPLg6IHEO/5+aR1hdbyAT+VamoF01I
JKQQVt3KqI7GdXxr4sY+XLCl35k+c0xdqcYb9X4NIuxiyzFNtj2lQxumNP7qcR2z
Q5nmQ5uxuuiara4LKxyHAFdclsYTlphaIM0RdhX5z80lEl8Rsfac/S1tCvTNbZZl
vot3JrsVQ9H3B78uQPjrWraWq9+s4TiklRSvh+sM1wjDixHZm1AkU+3K4Jl0OvLO
GD9GtLbro7TD/WTvddFMSlUSrt+W/FnoHSPDdyNz7UV+M/cbnbyP/TUt+FHyvU0P
a/yV/d0+TtSbQxmuGfWzdhhX3mC3GhPFnpO+7RAe6VTdvJcG/ftfesEG7v6reFpa
wVFjjdWrZyPgI6Q1l4SPvbzxT9f5XBGUjboQP8FLWjFrdfgZmqJfOzDTAGYYI9tn
3Ew1J9u7Id3z2incdZ4MGCoNJQrx//Ul35cYlVmv67SJEt75M/zYtSKzmyPe4OoK
A8aZvMl0ghUlakPGD67aQLWngP1OVXFGizKlAnpyg3QMMfxQelbpb3nPz7aET5G1
DK8+k+VLyCQt2pyohucUz1EWmOvLukNNMQUfXabuby2X9g/E8QmAJ+H8yfhbGdSM
jZUQDZpEBd6YmzcBk+egHh5oIkdT77PhxR+AQPC3cWSbTDhEHLrcmc7/4Z3+WYx0
5fsZXSoNXPBu++djxaeKQXQq2MQ0ZdfNaUFrvRYPtmGITuNuyDkAB53r8B4eIQvg
cvMTuVujx+PYLZw1xJ2xEs5Ehq3AOK0TGF1Njf6hLyVkXIglBOwMcdf7Ione9vR3
WklM33tggtMqh0bG09MFuQRydLw4nwXtSZQosqQz4ISoJG35bUY0vIoOVRkUnp+W
cTNiq/UZ5RqYZqrbbfUsZypMFElZL+5PntCMcRZiHO0JRXDmDXRIS9HvZ78RCUO3
ZGEuBfiEkg+ksEyzhwmqMjjeA+UNecTKzuVv/NFhwYHKi4f57u4WVoM2yBYLKmAV
o6GMtnVt0BjRPhVKMW/W1r6RMDRM7tS8zZv9xEGE8XvkxIVEKgGD6JnSsdF8c1H1
oIZ8fCvPrCw5dr4iHEPxbr0RIhLZtEaJNDYMwrs5rh6ApBYZQk0HlG/MYFBMM1px
luqbUjpWssgBE6k6gR7aDKgxAbohCtpbvvezTdTtsKXh55DnPCTqzvnZXDBIgUAh
DKyA1ZuWoMFCahIOJpOI/GiYtq9zzc32R4J4l/UnmnL2zfix3Fc+vZHVgvCcY9ur
uz/6m58vzZC80lROZTEq5SCzlVhUqf8Qa1V7wtZ/xwKwpDDk2US+Xh9qGHzlIG5f
cSKSAXHBe6H7PVVR/PhJ/i/aROLtARMieysRSJrMSObBQ9lnw5jjrLURRunHDBUM
VVr/b+2lhcMXv4x8k7B+3ceIs+DSJCIcLjUHzLtDkV9lXZZ5T3uNixFF4M2rWQbT
5ZwXGa+CEpGRGNtKmdaxygGNBz3aAyxDWwyjI2L2IHUz3+y88/Aj6Ies1jycS/aw
0ON+zZpwgCKEIIUSQpgb8C6htzay5Lhq1rmvfqLnNQtFPC5+FmCqH/nhBtffsnkR
12cIxAB+kgmu2HfuNjsro5psmlU8yiIyJu6LOfS/w/X5RYSXIye+Vz5N/66Hf6xw
TWqLc2pp2K7ao73g4cjtMnV+4YZc3dlyZe7rq44qCbC8cVZzeLD9nDSY+bUCGISV
pwpMQ/BiacpiOYbxrDZ7hRn5ngQCAnQYBsif5H6e6DlObU7u8t6BnPTWPpma4TU1
B0VNq9t9g4tKlIIBi+qireuZvVfYaTlqxq+tbydqJa9/EqHK5nkns5d7OLu2e6T2
55AvRtxfj2bUwHrnJSvH3I8PVB4gGN8nU0M1B40zJdHtXh1lPfni/K37N7WIUb2e
Qz3Bt0/65Kdhoea4ZRAvw4PUmDWC7hEXPE01uhLnP8QPvFZxxQGawGZ9BFN4U7gC
A7gCEspHfg4lNZ39nrF9doea65zw8fXifnIhTNVM/rV8cFbC7qoFP7bHFRiD/Fuo
xW0o4ilk9mI/2ZqR5pRLDDtIS7KXsWqZkwM+8y1megrmDXoDryFBwLk58MLdLjkF
cahKTwIPgVepd0mMEWfBFK8gTRrVSZiI+1MSXActG9c6LIEpE4t81t8A7ym3rMnY
n0EWif7Z8k1f3wbBMWFtqh5JhHTnJypBr/KrPOBv3TmVqrkmxDlCsXf2Pl1EDP1W
u1/f6K58zSSyRAJvzGpIPpyNsU5x2UH60yUrzyoEyFgEBtHAzKvs+qQYoCb5l8ad
dqg0S2hIbaQd9h7kZ6ZW77FYXLA7E8Wjuy3/L4j2puk/Dw6C6ZS5Ikw02KD7+ucC
tS+maLu64txZYAQ5EsGeWtvn8LvpbKs28QpMXIlBYfKSRU9J2iUYUy2O3iIRRA77
cVliBiCZsxpZFynsWSi4LkoVsEpk3TC1+y6VOt5jEsalu1BBnB/DtMzMlA4PgQAl
jGOiIxrAuRLMDYnDoVy+3kQ4YJixIGSYwY3DgZj+ehRhLCkQI5ECVysuOSQVnAfF
8FDAVURCfVPDL7xE+BPD7OQJMeCvETi3TcOHpBtC8HgJyGg9T2s+vbUQ4o47w+bo
VJ615HTLFEgJfza+1OI6q1LSJ1Ycq3qqtwOoSt5hmoPnKqPjde3cJvc8J/nOU/bl
aOBYVQdH6fq/JE9bkRpLHNKRuuhgZI0zgmVIaGTRwZ1BtFFg/dx7jd1AVq2dZ/86
POgNaNizKXfjluKBHeaBiP5iWn+APK6Ai/r4HGboaAmzSQA3Q2C9yxFIWEuuBmzj
eKnKUI4f7c5PE/4S7DZrdQ/3aQGdGek7mMBhMZudzWNljpkRzLmSkR3aQ6GD1X5x
uLttD6j0A4N4p7BA8poxzdmm6ooPu0FrazNddJK4rLlLNFuM2XFdWopYoBcSuhGM
lyPT8iyao/L/Z4N9fHnqd+0FSfqEUhGpIW74Lgm8n5DrnWFGPCWaWi8Nz0eU3C5L
1vJ12tQI+AggTP4jeZgti2er2g+HyT9fbB/96gRAuuxGzZ6yqfzP1m5RgOs1GVV6
pUcFF2mAvy5x8MFdzhEoCoKZ7ZBsXWUu1DpbNy0PKKzqBvW0u6pl/JHnfSS0I2Fe
teyy9k6M5HeP4r7tZlLOb0tL/QN2GGAb6SQ7Jl301k3Ve4HcPr2ECbNGK3mJdyKE
HEv1cIllbH7qXbha0GBpP+2ri9H9jcmHN0Swbhz+bnicAB0fUfUXohaJW5Uu8SYO
jObQmmcp6bvvNFXgbSoqVbr6A/2AdZmTUeCpIFAL9eXOkiSOD1cxVUnf0E4nQWI0
1MJLPhTuM2M/EKU9JU7uJd/DTzlsPlLz/1V9wzl8c7imfg1A1jabH+k3AU2PLLi/
5n1jjHfwQ6l7HTtpxBbEWFwrYa9eheuLXB/81jxLl2jEraHhddyFGY28k92ij14/
YDAB8g+kct7k93t30J/NhI6AVNhhcLHOEPSGylZdepobPu2TQj1i0ZTdnu9cPLN0
zi8FTLF/bkTENwymkA36yq2fjUHbTEg8p00NdE81rQdvQEKs2vA1GRWfr/rKWfKy
Cn/wy6xW2eVzeTnFFQHpGVstorhl9Y/irpOV5OSIiy9R133XEo7IaBeNA1rv+ygK
TpPQ4fD9NIGGmsCbT4OUBEec9ZgVVVes6OGiuXxUiUffsqRvafPgiIBuDrvQw1ne
8va0v9j/DV5HnGXHr9bK1leT6KSO2E0YVEmUB5kfNbtaBLII1ptvQTzmnRziFo7S
jV/1XOAo33DswmIUPbDATi33pFi70bkhH85nlrRcbUu8Ig7SuMUVYke89+eCyc8P
qYa0m/ihH8Dx4A0jb/dycFS28FV6FA3F3BJ8p9b5OGYD1K9lhx8J47ehT9iyTyG5
AFDZG2cN1yX00Q8tqYTRoCMu/D6VNsUyptxtGn3ozDXcw1sA1xMf/y9xZ/YZunmg
KGmWv1SuNMX+binkrg0v2a2BD0jFgGjdMBL9SGfL9S6lXywPd/FqF4UMT/a1OWWV
Ljr/8V9AJcZJILL4Xg/Cjnmyt2zPfgh+R3mcpLrcLxUB2rWChJFij/6j3VgDujmi
8QUHJX+eXlIS0q6wLPn+KivTjM6g3tosRD0OsGIv6LX41b2Fm0S0cRUTAzLJEQdO
XfrG5/LOHnRS+t/WxgN4lsOkkOHk0BWKdwYkjJCOrWVHi/gAcTbamsBZrVHtwQmn
weZAewiImEO4N2wpkQzEQYxA7mftAaG38UM5yAgB6+8sK9kPFnLbxsAxEWOUO1ab
unS5mWqtGE7k/xZzk1bq1YSF5ST3vF66r/TuUm4QnwftQcGFJpiJbo2P2cQL1oyM
1thiHl1jXroYae0rdK6iegqebxjdHn0vKptBH7V69n/+VjHxdJwyY1+OpyhAjvnm
TKwKLFMLX+s8+6WpEPIX9mt1uEDeWj/iMA+73qSqnUy2HQ2YUXur3GePWQ3reyiU
ujh4pVvmEJwqpNceQi03NG/cO/P+Xfrb8XNePkJlMvlZGYGxEpafsJJishiAubD0
gbh9nfLi5kW2faghIF4savCOhX6G4dFvjjEUmN2wMX+AhIcBU3/yGBCfa2xhvWKV
xDSM7dLjF203aMYFWnKC7cy//5QSDDJH+ZNGHbeDgvohVovJq9abGNn8OJ/HnYCa
PsI05c6ACuMvj+vP+Rj/+ClJXuk2cVvs5Xv3jgL5GHS+oH577WwrEBIZCQ19kyvv
WjV0mbSLB1kQzWhk3XvOlfcZ2C+4XNWk2ma+vIBGNwvGFkkaoa5xg/taP8QXmnXw
EGYLL9NliMWgVoMb3i10WCarJiWwjlbBz37P6WRqpqR3SBlc0XuljUCLgRPe/UXb
2ywNFBwJVw5Af4cMgSdjUxNoHRA19oApiFr9VkLk7wDf5jaf3nk39TUJP81YOUYc
svpBbWzcHAW0i6N6JhnpY+E49iFoBbRWkiaZcCWJVpUauVmpDFQUSqDKcwHaCadb
aOtqSw8kwFN3DRcFjJWjzzeum5ySsJjs0uMHUNRbfXvFH39wC+u6N2BbTyFouYmg
LcsJU10jUhtlqil91jR6nGyCthWLCENmO8G6UjpiZQ9t3X+ZP0wpmw9TEAhb0XDt
zLbGYxbF1l0Uh4QmAaZWhB4MUS0ew6Tznw2zTgjzNliESxApNmgcTlJFBQPNh4M/
pVFfskYeGbolO6bsPtcAOCqCWBFMEliRSzUaN0R0QYTtUsa5RKoy9BPKblRz4/VN
dMr16dh5hLPmkLnubsCs+Q/3Ezthq9e2WEhL2DqOZ+VPqKvGandD2Vcubb9zWWvB
KiA7Ud/e5Cl/nJ1rT1DUg2KIVBGMwbqhTCgXs3s+AVWNiKhIEzyKsKa5FNA3yQnZ
2qtOWSXIXlLUG6I7x3HGA3xV7vecM4XQw4IdRccczf7DM6dOyS6+QJAggckyDXQk
FA0qP81jrt72CtzWZjoDexFtBUj94xNv2SWrtJ4qmGFImaRVFXxVvQozTuG/s5mX
9jVvYuAo4zYJfuQjwApKBTiQzTYsznarzZrWWo1Dc936E/NfP6kVO/GLQtYVxCJR
NRW8Mu99CDy8ALnLIzlIEq5psavRYcMkMa/o72ou39b8ldobfbcVj/Bkk0F4LxRu
Z7CHgQ+WUpdUMnTeIpOZAUjdneik2UQMaX43cLchWOoTjllrw060BCZQwS3tk9Kf
f45Z9U1wh91enFD4uDLlod/Acp7TkQ3K54PpUPAF18BbeWJHHiZH4KUgCJRNQxZQ
UfAemaUwC2UD59hm6a16Y2v/asQykUC2M3dVYyCWdPo+s5iYqtKJ2NENliPUxO5C
oGTwV4aeY39w8AjH7iVc9CoCOBwz/j3Gkgw8xUh7Nidi5ML2Qcv0Dq/l3dOxi66Y
owveFzfivpT3y3pIfjCyB2f3dk/V/76Bq6xrNQVjL752dAIPjE7OZSYyMcAFneIa
J7reLsCTRfw72CFbpNeFvF4QgS9nkEWkMcUYO6ZDHB9+OF4hs/03Qsd9WhwRo5bW
m1juBzKtj9QBUpE3bOMcwrHdWvedm7Uw8mXxFUVtzfIvJ9LP0fQO7mxFqkz7F68h
NYKAAtt2j0P6K9y82kvFOAsjmqtDvHsAhLtmykyHsXu27mZt66L2Q8MHF0kv95m3
LSvMkAYxDDgbBbxJMrdnpRJctDxsHG/gYFcHq0Uanz1pj7Df/fQe35eRL2qR3/W8
JAizNkRE168Eds4lAj2hUTKbSywp4iIlEGHcalhyHr3Po9KdLq9/+5lWZnaLofD6
u3IzfO5SvKHK99qelyjeDf73NEayyPiGH87U6i4Bg3jEvQ72gATU+S8XTSyZMWTw
l0qGUrz8O4WYgjVzFxUZzGzKD76yKMlxX/qMwd270WWtFWxu7Qx1QXa7CgMdXr8N
rX3Qie8HaSyNvZyeJNiLMcRUYN7IMusKRv5oSepJ6yTBioRtIc1wSA13SNZC73hv
AsI4wk+HVVkhsZLp2oPdzLOLEKhI6qCl0l9feZwMsXR3vroIZytcGO5qGwcrEqcH
h5Mc2P/aOyAW68M/FeNEX2j9/n2slXjDIVGr64vhevdXSXSwNQXjjBG3AEyNxGYf
aYb1gacIExKSZYArYJwVPTcjpMlhDFCDGbrhn86hDrjOMTMJ3Wxn4smN9CevLTa2
MGUTrp9h04H7oOhZuB5YwYGVrK+05yi0DQTz0KWBXauJYsOgjIRzHlQUpvmucRSD
CyuD8D+xo4Q5RrRmqlAtJqQ2OFpeR7nxTc+EtIyFaubBQhBDYMmF0u2wZ4ChuX1z
XAd3ODPoC+PgK1QbNQgmic+dJZIUYh2yLwftAI1PY8+CuX8oJVsTMmkbUN6I3aNJ
7aBSu3QuwaEIwEbel9sHz04FfdXSGm6l52ztBFIntCstGDCIB7FO0Q6Iqi4ToCxE
kJtFGKt7nxYFIWMp6yOC8Trv0F82Akc3Ul8SYQKX8+MpIGWdvyTirNrRpkLhJZny
y6C4baBHT9YZHFP8KI9EqmVS2+vrKpLU1weNt4vxzSlY8UID3/ATQMAzzd0smRwX
+0ox7mu1st4El5laSnWceQ2DteLhUGe7znEVAksuzFPnTBltY9qXz+3ElfYYZyq2
h80JqWQVj58QKBf/I0sib1WBXw3KXabyyUye9zeH06o88KfhU6uvMbZZKhksQsCS
oqj3PHPG73kaF1GLpFJhVnRQGuIPqpfUvic9/XsOU3OLl/Kf9wCXWNDPYoGSK7EK
PHLviI3yV8yLGj05DlTvWDm73+z151DiQ44LnxEsNkNsmjV1pRy/J1wSs7cMeFjk
1cq8lzh+c+LzLioBsoOI7XecD6IOW0X3xP6KrVjfA4yM1x8aqdfsurES2wqNFLOh
hNbiaS58ua5aDFPNpl8dpTC6+fkP5V9OTIEw3s5xUqDCaGieLq6+NpE7i+PoCRaU
m7y67JnCLTCKwwLbAvvz2s3jMLZj0hZqvPqk8sONLidYL9lfpldlsPSXWZ5Hxs0b
vXCSLoCMXO3YHmPVbgjRN9UVJffDs+qRprZNueLoHtWC1OFSmyJd1I0y4fTm/iOJ
RV/zDgPpJmx9lXvCJzMXz9Hh4xOdx092u/6soR3ji5pU5ZHq8IVLIes+Z5nQf3qC
13LoI8svi9KUdfwALms7YR0KXNIPO2QA2iG7rrKoR2J4THtzbHxAFnpu86C1hxD1
opDf16/uoQIWZ+aBHRWEZSuq5CY014RJ+J/XvAfcUqCDf8G7PkIsG3SCwlQL6QkK
MzJZetUCAjDLNWdIoXZ4kWo2fnygbjVaui39P8J/VRtN9pxYZC/YTjkHaqSvIgTi
PhxNOmWsFMl49utcCtaxhdFmX1yr8NaTnfZ0AAVluVZ/SL/+SLgk9uYZKTlszJpL
ukg9cqSJW057VGtBqtx3BEPA+0Qr7TfjUsTckZwDtaFKaE4vPH3W8+pZuFcoo6I4
3P/BXb6SceOITfN7sl2Pr8/CLzjpHF5EEr4zBEaVVheR8HfUyzc0oB3g+0M2mIFk
WXIHpWI7I4MSsRC7dIT65uVI3WtZNkMDUWTDPogz1FXL6I6t7HLHwloUALARftUL
tm1XIumgazMCP97vai62YhKXR055RgybIfpGan0uGxp/HlkWg1iuyWn9i3MXf8Us
lE1H//X10WR3wZ4/euqKdGmz7ifmJGF/DtLi9pmB/o+gxDzkdn52o8NFLY9ig6l6
8ZxzmACZ3/NC+ZWZJSOqJlLCKoRcPmAb3UwSNz2Lenel4a+qgSRG4cClfCkh1Wju
8FpzwU6P530amTbQEzUy9GLMHRCSD6wAU7nqNRXlhwy24+9RzU1BXr8Q2mIVkJOd
7v8QGx/NLHv4yy96kvoY3E0MSpwoCdQZr+itfeKNFELZB+Hq09rtxC8ki1I/nPZO
SuaYxKhRf+sWmzaYOIzFBJ/VZ6OEo1PXlE0Yq4AYxwFyiQ7WJtK4XIZXDou2Cv+8
TvKwRl5kSxWIoOTUm4aZj21Sn1+W9u2NL5h9O/GSvoun1mux2Cf6qcapIdQmRl3m
cVepU7aHPtWOPq/3NYa3li32znhSlKeGSWt+hJO6/0YG2J6hINbK/GyECQ3pd80j
Nps5HqiVxFO38iQfcW17XPsKqfH5OSWSICTksQyQZB3u3OE16mL13oKqkUQBKqdn
q/CuWwx3OANyjjrQVC8dLeg4YQiBEqMVoFOJ0bpCqCSEtVlPsrDuF0G3B9gyZ8bA
OeoBJMkPtHsK+PhciHinqk8DCJLtp4nv7Wv1x0xaHPlHQVsR4HNi3KYs/SanNVNn
PfmhkQaF4GwcUAa/Vcb3Vka7OwBHjfbC+Kjf7JecmMgv59OBJ4EgaCap3QRbuo/A
TpNqDBxQ8kWWzcTPFwTNChTQN0Irf6EwTMcVrSAAqQ7codiago/tiHNVwBCXJSoJ
agI/uATGjK077tM8Zuu+2n/HrJTQBa9m0Ml/N9aM0kc8ifs157k0VttaSbI0os/v
Ooqb0fjxEecRfBDVIxbQy1gOoA8tOej0JN/kEYKReRxH8W2kOJt4nj+I/pfiWQo8
0JUiod2/6Pg9Jl1ZL+pxfIURV9L4x8ffNhl7Sm6MYOdNulVr6SgefDMD3g5CturM
Sr9kNDOuf4FlnE/MyXga3wOS2kLIxq9Lhx+tprLgPOqxEv0dbU9F2FcWYEFAIiQq
v11lgC6NgRGWTmLe9EANEzak7RyR+BOtAz1t4Zg2PKePFvfkRyOXJUygiwM21Cmv
2bOACWijPK0OIeqHOzb05aN/RAKaPQPD7IRV9iMdSB5yjFZhlIWYoPGK3C6O8xWf
EgcjGGZMLrQvs8P9MY3RfDLqA4OQC5QqyvHqHS2FBzrMq3/S1dufzojf0Ss1/9Ud
csduo9S9rLMhsMPSS9DNjZ0fa33nVbKiX2w2TpK9L1jiR8UQRJCiWVLc5ZbOGfOA
7wgm0h+dCe7JWmUOog/LwKnen3kWYCNbiTpsjHxA/SfXRSc9kqy0NZ81TCusYhEv
ant7LQS2nThOOLAiEcYNGJeK1DXlauLHsu5r5+zN4dbcXIAPaRk90Nk3y3LyqTbk
T6Zzyqu8MLn1ZFowlHqhI4XV4r+GMcf2j1pDzzXG+syVjZIycRAvKg2s2zbhanQM
16+L3eHz194m/CavyIPNUtEJLR2tAXfqz8/iGA4h/8VX0tWfGmlXzC36R//48FL9
xQjj9N5kNHA2ew6801dj9u7TN8kRZGrx1OJBzVQonfbLtLABdiyaVDRDpX7uSLyn
EFzvSoiWlqP5Ir4SJQidBqHxj0RcHchDhqm5UrOkdSzO8wkQ1iygoYWY9gRSeZIp
yrN9tmrCVIB0ckYzOLdSgbYLjjLRc/DDhew+zZRXByffYYC/55nco/Qg4qwngAtG
qlsM8rl8NM1pVLLOOXuZjsC+iYXrLQyRXNrVtB9BK22l/QLyxN9GwSUya0BGvX0z
3YEnR8iPmXqioJ4hGfHThCW/HOl6ACLagY40ye/2DhdJ2s4FAgsN0IJ5otWihq+y
zZvdE2A1odSNb6mNVvtdixBAMtQJd4T1QMsMKZTNDchbTst7Y6GGpwccg3WwnKk7
sq05wwil8kHGHGHxraAFIY+x99VlO2votFAWvcYLQGWUNWb4KD7gD3GPrLOz1hyE
rk9mo7V5LY6Xq8zU2eKU1SaW38YYiVEqqbbzgwG9KUQT3eaboqynz47NcqfkmCrj
rH64G/Ym8ep0uTe6qTso8ufQphoQcntDAzP7ClZxinWQleNxaA8Sl3rsnx5/kMU2
v8wpJfSHM2YhCwTIcp9tlD0me0pVchhLyD/WbH7e+vsrxB1v33u8p/i371SCnpeQ
L66MevYsMcdaGL9enqfUnrbfk1lHwbLI/BaAXCrc5ApT4QPfD4DLGSrVZYMneqBl
4IO5iLGYkWm/ExF7bdMGeVLsvz4SBiSIMUDVXRnPYQbMp8nOqquXPfV4UF+YF4Wm
Y/MuWs5saOwKPUots1Mb8l3sOHvGBeBUDPiuEifxvO57edoSyLdpMfpEdEYZoL7u
lhR8tXfPR7fQvbTMvWfCHedLY6XhMPnL5XGR/QR4Iy0GivsdR7IHWomkpZWBffkd
NIK/Nl31usPMt7OdURuMp5uvwBqfIsOXhX+WIryLGcxn3llghFemSxvIssj7T3Ei
fqFmCYv2tyR+t5UwBhl/pxSc/119U6iPmtT+mWCF5MxmQxwU7TOSJsSb6k0oLcNg
f2vEihltxB6MRDvIHjSGqtVX5+bp8bxEDGIdVJkAZ4YWcDEsy69hJSZx0pQoQR7d
1zEvi+1KY+vpcWJyURXZepx4jFx37qF3Grr0wsfr+JbM/3zFXbZtliOgB5fdxECL
O+D9nS/b5pI/QSH9Fc2VM0VHxTv2bvnFx+jXNCXcSC1fIPSo5hGoklHu38p1cIsv
dOVyKPZMR35DLAI72ALXF2BSF5T+NzzmL1VdFLPCmK6Bgr0ttM/WrPlDZwFg39rE
b6QmfgRGOGEcxhNik9fb94Cnh1nSu+VZtAnorP7jzusdU8aPOUpsaDBQKIFi4/bG
AUblnnrGeeoMK4U3J18X/dEBm44U94M/m8WV5bVj7SKoAKz6LpgINzUnJBylBovz
RKszuVagD1sT2WWTFmdbE+5PGSoJ0s9uMeweX0gbwnUPIVFqsCku0w7kXDPLh9ql
6U0mu9UXcFhjQ5Eb1b1+MGMzvENXxnJIY/tDidN5bhWV2KLtFZTxnY2QQx/RAxoo
1bE26WqwJyLdAiGz9LtPHx6JxuELQh3C2CIuOK0QRlCqFez/QV3gJW9b9nvcB+Ul
C91paLRGcDEv2NdhhY0x/wD0Qxej6o9t1Ql+MdA9sw4dTBxzwLZ5HzyEdnXcZUaT
db+zGkxNVmi596QE2QjkvUWzYOsNqsJe3J0q+DEoaAmEOsgkLCuFozoeX1Ep6SCu
V9jkqkDDG8oG+2nGalUN3PhrMp/Pls6DlPGOnA8QAKG/s0QJQa22zUwfGmjVPhPS
649R5MHZe3lenrIgN2SkTOV2PKjL2kWB9LKxXD9u4qBsFhkYewMhEfE+MDW6dn2S
NCZH/lTx6QknrMHDF7zf4Za5+rTrIQYtpCtigYDZ+RP3AjA+hOFomX5QBJcpxZj9
KCBtuIKqeWbuIMqU98/7wBFZv7nKovuHMkL22urEc8bCY1qfJlCaw64rjQLeDEqJ
S83xZCyBSwTkM2yoROdMNCJKdUo45uTj5UJcBMPtSE7W8x8FSDrcVlMMnOaFYyTB
jRG1ohcTwu7OuukJyuRVFkfQOnoyhiutuJV8OBCCexfzsTgve0/vSVOvw0GcKxTH
nymaNbrBdWLokzZ2MYlnmDmAE0KRSb+RhxRIanx0sEqBrCiGzgN03AO5g7wni9B+
VysL+IGzhZWfaBtG4sUHU+T7AUnB49lV7wMVpllBfyhxB4JUHZRPvu6WjUjBKgGB
t88iyPSFQ/Ubw2JKzg6e9vRdbf+M+r+KuC3ngAVLVxGpAemXLXBtgVWYXBgtDbt+
P+VVHvW2MonKq3Sc/q71W7kKv6i0iqUlGUym+ehk51kmkvU8yvs/pM8Vb1PCFY0H
7INjnQoaoe5Iu3equjZlFpk0slz4vYXZPajZ7Qa4+eOzJS5xfXvCv0nULLsJFiWF
YOBWrrHBJaDfwzRduQxYgNljkGJbXp4ILmBZIJ0pwugXkc/xbgfJ8a3ix96ioHCl
SR+WWgBN0nq2lSeUTfYkizyOU13xa1VSZk1n3QTmbF54vPLRG4CedH+U1Sc87GmN
ZiHCQQXZV1PfwP67MjaRmEneOo4gR4oQ8NJZeiJ01m+Cgd2n6oux6SnVUSt/2Rm4
JArq+KhM8XTNfJaNnHKFRn5sodDBzmgUlTcpmm2wcqA75kaOT2PNcmRAzy9zNur2
X/47GSP5E/sPzrR8HUfTn/l4VT+dfKitv9nI24NIRY4swlvGRTXVj6kaXfpShN1z
K4KXiO1/w+dhdfffMzlHwtKnev73voWVj4ACE+swOwk=
`pragma protect end_protected
