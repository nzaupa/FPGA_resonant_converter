��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l��ӡ;h�>�C�0��-#R�&�`8��2�_E��6�kI�n[�{e傭q�wҴ� u�j;hKb�>�$'���a�찁�l�f�^��xGL�Q�ɸnp��݂L���nڜD��Ve(z���j��ǭ%��H�$e��~~�)��/ޛnI����ܯo��{�k�yl�	`���#•�<#�`��L�C]�Z���B�Sq&�$o6�f�_exa�0���B�\j�kPؙ���wB��z����	��O����IJ>όXT %R���yX�7\��~:�F��4.����7��3����!j������κvٚ7^�����U�)\�m��{vW@ �fYT�5�����󿪱�lU�s���� 7�3��5�9(�ʧFk�]�6ҁ�7&���l?*�;��ұ(�q{l���A{��4��!6Y��<�}V� V��XW����2ym��C\lq.�z�18�G�~�N0;��k�;�H�L��)���Oɣ� �7��x'�8:��D$�s`e��k��M�;�I�����b;����və��_>n܉x��J��Y���$�I��j�	�ʺ�/_�x�;?�I�^��mL���S,Iw���K��M]���Wf"��MT"	oEC��Z�l0F��_�����?
���|e#��*���9&%�@����kH��;Bl)�˱��[��9Ta��^R.z�=z֢����%q'k�]j������-����0�&�T�S�7p��-4����z��3ױ@fN���jC�4�f����9��.�aJ2�����_	b6�gA���_��Mc��us;`l돍UH�Z��6/���/�X�T��H����Y�M�3��h�j�kڨ^�m����(�������dĴ� �˴"i~Y��BaU"r�u>�i����4�����U�RO��Fy�VGc�\8@`���(�	��;������� �_�)u��j_��>B~Dv�z/��MXY���؀S�-�{�
1�=!�ԍ7�������,�X��2�Z��<�2�W�q�Aj9jN���āy�T��SBK�|\�r�2�깜�a|P�ƯwY����C�E ^k��y�9g�6`-��wZa(~���\=�dm��8�[�ߴ��=SDP��Ţ�C���|��_���HDE�r���c��7�U_�]Q5��g�)���)��;�I<��|n V��M�#�|��Y�� ������N;qO�i�~�bqQ�$Q��x��윯飒���*j�*k����̂3�S�N��"ew� � &�/�o8���n�卍s6gk�ɵ)^��W�7j[m��Kff���B�w�V2�qa�?����>��y,	R�j�a�U���{i)F�����2@� �)$�E�_x�*N`���=--*jEW6����D/� ͜&�B���'�㡫V��q?��a�;RS/C�J"��͍��h��n�k]����ۂ����o��Gg{eV��\����H�7Yjkx��Bf.�7>,�Nj&���Z;K�,S¼��h��\U��U�l��(�옢�M�.�GKz�ݘ��J�����u�	C�̮�C�O� Lb��ܲT�I�ݳ���G�����`���`��s�t�yH����_'���y��诏�@P�ix-w�)|EL8 �w�+ p&�+�B�zG�{U�Y�\�\��j���ꂤ�{���+P�"W����� �mˁ��["�`�mN��k������/g�8�K��&�$�?�^�y��:�������*�Cou���d<t�����s������`Б_h���4GΑ�?Mk�V��
�꠱LS��H֟��?U�3�ϊ��ʹQ�}��������	n�����>��>�i+�}<S2_�J��uu�%pĖiB��//7�:7J�˟bM�im�B��Lz���䜚2t�#� ���B܅�Ԍ����T=r����"��cn�7R`.�f@#�)��1�y��sl\qZ;�}�yr���h5���_iD:N~���O&��&j0\��.�熙�-Jʒ~�=�ƍ�ٺ�R�5�>��6()z�FQ�� �%�i�Ò�@�ҹ�1���H����om�-��d�:�ƪDY�$%��sY�SaK����XD�Q��_=�re	���zqA���h�P��G2Z��A�5�����p��6��*O$���a�c8#��]Ys��n��γ�������MD����։���F&�3��	n`R�F��r'�0�-�ݥT�1��4G�%WP�MqU���E��4����`�**8l�O�:��Y��vD� IGj~R�)Ġ�A����'�cJӊ� �]��4x��T���w���c�rk$.�`�� ��;df_
��?||L����9z{�}e�yi����E���]���
��wň��b6s�l��JwJI��٣sY��ix�?�������gT����"�ʙ����:��%%���g���f}K�f��$b�=P��+wNª(����o���EW�BS�ċ*s�؈ܶNc	e��� �)���34bf_a/p�qO��}���Y�ZU�}��[�z�e�*0����̊1�12<�`�����a���TO��!��q�'}�`f�h��tfi�����v&'����T֭�Վn���(.�M���7��u=)�Xo5�HT�'n���*�x�D!.Uņ DѳD�H�O��#8�HD���=r(�a��g&�`߬X���x{�ː��
h�ֱ�f�ly��vUdK�If�Z��"�Sx�3�	���p\�<A�Ot�c�3���hB�+M�h'�d=��ͳ���Ǝ��_�}��wM�okĄ29
�x$���T��8��1?>I�/�:e0r�Რ�_&Ox�OH�c�Z2\j4^�W�޷���F��p�{*fT��,Z:C/��L��Z
<������Z��A!�+4��q�٩F�sP���(�`jb@������ͣKH�~f)�dc�%��*���&��,�>��.)���΂�K-v6�i02�R����с�kg+�%�Gd�Ȓyh�r����^�����u�>*3��|���y�SC���*^ �T��3�9Ɛ�B���Jŗ����$+N�f�+Aṙ5��]+O��z�O���5.��'����e�n�VU�@���pکz�Q�(&��A�n�mR��)�9e__�ʜ<� ���ǹR�-q���د����T�..F�n+�X�Zؠ����?(��:��\o�>��#|'� ,{U>d�(bF�o2��b]#��O0���CE�D41p�&�71�TR��y!Z(�n���bŬ���{	�ղ�ǎ�{���~�|����:V�oMM�+���Nk����e�(W�8O27�����Wbk�b������2M��3Y6��s���QI�q�N���0½�k1,�6�k���V�LbE�(w��g�Ư��vN}�tc[��JBe��)���q����6U`�2@8&�{�WR�$H�V���u��ۣ�Є�m�ď)�;P�]t�䫒6� �G�}L"k��1;"��,&5ߒ�W\�ph��y2e4��E]�%ns2+��(�(KŃ���m�z�ZV+����v�����e��>ۗ�ՙ�|�S�55C������<��+k込��g6<�����v9=��ǥF��o�[�~��:C�y�Ƌ}��fW������(.��%�-��K�fK?pU�d�^wq���M�[���X!j�8$DD�;%�3,�B{ȋ���Y˚��r�m6����娆����d6��2�Ia/�ӆsL��a`���wl�������v$��tV�Ɇ�� ��2��ĂVjQ?�ݨ��s� �N�?@���T9m,6l,C�����T�TPTL��{T'�8*�q�6��hH��R&n�(��^/>�/���� Hj�xd�Gz2�O�Jj��B�U"�_۽��TZ�w�X�Bj��n�zCLL����ۍl���_7X��Yc����&��蝻&F�S���$�{^��fBХ���1��.�2bb�~B@2Z�|3[�Vo��U�=�ߝz�A97��Z�h��:��ZǊ֐�l���QB�<@$MKGTi5z���3Vw�Ű2�y-g_��~�c�l�=����{����Eo�.QʯMS�VM�
A���VC�,�VX�΃&�q}�qݡ��JX��N�Hc5߮�����JlP�ڻ6�pԚ��p��]˗�����Igf!)bm��F��0b�/���s�P��o&�lfJQ9CL�[�$@�����,4K��ž#�A��R^%;���_�(�Rꨕs�7ł���Nw�Ȯ*�{�D�Ifu@�µ�:���eph��,FǍ�1�^sl�1��8_b2=_������8+�Z�Խ�����,L�-`�>�-�tɧi��5��0W��۾T��w��}�ڳ�L��z�Ǹ|��7g ��e�q��3��z{bB��J^@%�z4;(V��{�*��Ñ�i�_-ސF7��+t�5�Mso��J��4�jeE�������I���(l�]}K6��|3�t�f���5xX�W��엏c|�=�%̈�S�?8����[��| ;d݇��>�I����Kum~&$����Y��e���
/�-MRV�����d��x}D�\X���L��?��#�_m櫼Z#�64��?Yp��~#�~�g�mnq��AR��y{�K�6{���")�m6��p�#��V�8ßR���_?�.c��5aD�·$��Px�b�1ԣ�j
c�o� ��,�w:�Z��^�g��!�fM�E�L�UBb_�f1w�  ��^��6��i�C��3�3 {<s��87y�/��j�xx�d������$�8T���S5.�e�t�Q���1���!@>V��20��X�`ˤ�+5�㮘dy���8^�����|�G��;�9x)2M�jE��o
�mj���Pw�V{���R��K�"2��'�Ӿ>
��A�0��y��Wm�Ŝ9vs�h�����1�\GS�c�h
��Z&�Z�A�)���q�1�"��%"Z�գ��p���%��'"k:X�v=@gHq���.:t��0�"a5��b�e7�s�5�4��f2��Z��M�7�:�8�T��_�X|,�H�^�� s��3��u{v1>އ�����juS�J����?�f�ŉX��;�bo��Ա�NAݶH���P%]T��������������[��]8ZN|��\F��F�d�
*&
h�ᜊp��f��U��¦H�(�����A.iR�߄�ά8T������w����}�@��qQ�j��WJ��U�ː�чjBoO �`��{w�X��㥃eRů\���Ր�ô��)�r��,p���I5~s�,�W�L���ߥ���n��kpsjI`K�H�!��3���7��7yY͋�Rw��-�+Dl6�:�2��!5��Pz5d�
[�ڡYҘ��-^�f�*����\e�}��WB��3�2�e�n��F��l��Ջͽ��	�O6�}�~��7�Y���I=X�4���h��<F�"'f�&ؽEy�)g���^��:L��=O��T��[�10�O�*�Уk@ ����#�nA7�䃩�^n�X� ]��E�X�7��