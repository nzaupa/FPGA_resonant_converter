��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_;�"�Jg�4ʏ�k�.b�Y5Y�1ۄ�vWˈ���Ȩ��=HB� �������3�Z��l@5.�1&��5�ꏓnn_��W�<�^��^᪪��Ѻ�$�[�𢚷2L���I?�l��I�?��6)���;��f#��)���O6�
Y~�|��+q���&d�TD
����A#^��9��h��̢Z�ܬvySUk�;���/�8�E!K�q�e�I���n����X���s#ʶy7&6x9/R3��<P�L�L�j�0�P���lm1�HJ��S�>��� =�9Q�F�
�f�ХN�:x�C�r=�����t^����U�M�ݟ���TA������׹ �zU�K`�s;���r�����Ml��a!�?���6X	���Vz)�w�*�
ɱ�����D��k�gdK�ys��_,� 6����C)؇�Rmvuv����M���5 H�?y�?U��B�������.ג%/�tFЫk���f��e�
���f(���� ����\I$_�Y�Y��(a����2Ab�)�!G{'m����+�t	�IBKf��AK��
�M�ߥb���g��݄Ɯs�oQƮ,��|��b��$�(�������g�����!J%�Q�7ғp�+�ֶ=��q�X���@E ��tb�'���P�F7X�E'���#:�XCG�s�L=�5�X��X����s���H�n�/��4�;~���a����*���m@M���8J���)Z���x�Vs�l���i�|q˙�����E���$Y��K�-̎�Z�J|��~3C&k�R�)�-Q��Is�Wpw�a-��t8�@�������Nz��-��K��P������i͞�ͤu�v/=6��@��;��p#_C�>���~���5�qK���Je���4��Rb��Yc�qj~���Oզ�מk8#a�@��a�	n#up�Y�x;����l�k��2�� �7����æ�
T�:����k��b߸n�j��6q�k�N�}�g��g-k58!���;�O��P2�0�P]�=w�򐒤%7$.�=��Đau����±��'��0�� `����
BZ1 �+�T�{;���~��s��o�,F�1s{dĖ��yg�1r����n}>�p�Y��L���T4Ή=�����ً;Τ�?�&�)n"���ܐ���
��Ee��;���tw=�ܬ�]0 $RO�P�������$k䀱�;��F0!F���֒&Vh��5��{{�/y~�x��MI���������X<��+B�	�����pSQRAF84-<-�����?�j�><5�����>B��U�D7J'��%x����4O��{
"^���gƲkH����)��
�Ĭ�l�ζ�0���H/A��:>���!�!43�G�r-�dZo4��H��ةG��[�L,��զ�$Um���xLO�Wi0����ƑF��n�FK@��l j,�s~�Zg@�V:IO���^��_0���0��XX�����#RFz�m0�j3�� �.즪��ba.�`���s\"2����H�n�(�݌l# ��5�[�k3�Dx��8���Ђ�g���zoL��^b]�"��p4(^���`�ke���d8�%e]��_��3/NmT�A�.]���N(6��հ�]���[��o�&�i
�́�g���'[���QV�6t��ZRQ��e,�6`��u
ZO��;j�}$�sd�l�L��!�J%ߞ���8|*�f�1g9ڲp���ة�p':j�DӸ�nߤvU6Y��O>b�?���*� 9^��?���;Y�����T�b�y�ޚ���GA���[���]8���$�X�E�>��c:�U��\fi�/��*.Ǳ����c��V�ѕ3�������+��%WR�U�T���.�;}�A$"a�oP�M�Ch:Uȷ��V�V� $a���E����C���-��J��,
��i=��E�y0�lZ���(D�=�\��P��#����#�V��u�I�+�=�?ڢ��T�F�!�a!EY�����q��U� ��n�z��t9"	w�{��t��dM�Ɩ3�d~(c���ܓ�VrY�O=��e5,�H��褪�nʩPr|4	���h����p^Nn�3={YJ`���y�cwq��c�l.
�P$���:Gj<�3�v����.ߔ�rk��zQ������/��cM�����]��E��"����>�,=3/�"-�[+�� 0��fHV=���)��Y�8��I��`mM�ķ]�b���i�&�bqy�O_�ZR��Ḍ��?Oa���V��#^&j'/�!� $7�>P�v��9m�g�΀��Y_��DP8*K�V��c���ɱ��	7r)ܰ4>gp6��3�����LP�g7��Dkt����E�[1!o��]�}���Z�B����h�����$�V����4���,m�{+����G?���wet�Oո�n_�- %��!�m�PG���n���!��������Έ*�o~��H�(e���IB]�Y8�4n(ک3�zIY��|�fdX�💜��q�n�~�ݕ�ʤ�&d�F`u^�����r���2������s��6;��Sʠ&!"9��6!��!-���(�ᗀg�e!�;��a	�l�ld����3U-���=!� �ț
��I�����o �P��dJsy��t���΋
��Ë�&��;J@�a:�
g�z	*X��O]�n�墈A�=Z�U0�/��_b�����OZ�VT�\�����B6�SA@���A@�щ%'��.�t�y�ڷ�UV�I ^���N#{��"!}R���g+=�C�U%����3f*A�&�΋���c�A��ᴁ���J�M�&���ȉ�ɚ���R�65�����s�P%Et�T�*��/��� ���8D^�Z������ÿӢ}C<Z4������@��!��#f�mX��/��Q���%XCf4�5t���� ��F�� ��ㅳC[4�a�\~P�/b�r�}.�7EB�ۘ�E���؅:��=�ё_�)(ruz`���M�$,m��Z����D��lkTf��e]OF��J�;�d���`�����4_����x|1١�u���⣙5�ͥ(i�z��ԕ'�QEeVF>��3
�{%H��u s"%�4d���L�K0c�m�s��d�,Z��Ж�|k���Ş#��UdЅ��|�i�e��r\OHł�*��m��m�*~�$�;v��#�-������G���5=�l�������E)aҏ=+�2<l����[�툐O���t��]"+�i����`u�4O(tr���av-h
Bu�W_�~z!u#����9����ԁG��T�S�:kwjS����d*j��"��p+�L���k�?cT�e��$Z-T��bg��5t��3Ө+���3XP�)����
0b�%�aP<0_W�'+���ӝ�`_�S-!zg���� �?�c�����;��׹nGJmUf���f��<�
S�k}���� ����ؙ%W���x��&V��gI ���*���l��cw��<��h}���?W5s?UJE���
� M}F�M���߃�=��� .��.���y�&�)A t�R+MZE��v;�7�fD�UD�ݻLk��bh��0:�� #�ν=%�I�(�`����(��V�I��s��E�����=��2Mu:�SX+E�e��U8)�9n,u�z>��rm �q
m��f�U��t�G`�>��N|���Y�mp2��Q
��?�<&�>���KB���� [�՘��+�"��K��*A��m��Pu� +���9�����Y!˵W�9lܚ)�t)��wI�E������YW ਫ�8�֖�H�Ze/�y⿘;f�s2��x�M�L\�(�饱�d�l�*�8����Eo(s��Y33�zVf2���'�1�eõ���\:�	��0�9zNv!M8,%�x.����"NF�X��X�;�������f�'�38@:F�$�6�T���$��f�[Iʣ"�	J��^�Z^��ٖ��~[�5�����s�K����/)�2�l�G�#����cy�K��(d��J��� Ӗ<d��梲۪��D�5�VRe�h�F���Ij���yk|q Ѡ�Fk8�O��J�H���.���b�Kͫ�q+�4���^��%�R���~w��_�S\{z�v��&� l�Ñ�4CDx�����p�̫-jg�E�~���2�t��Z���O���r��cw/��񥞅O�J5AG�ee7��.[u���.��/�O�Ճ�a�9uK�=# g�3����	OL/�!	4��}���6Qҩkƻ~N^�3\���w��?DW���)ѯ@8H�֞�+߿��$��rȧG�:;3��}�@������|�a>
,�\�cEY.,M|�E���9�Z�C䈾D�n�$�� ��g�wz�y��� Up���-�Xgw���mi��U^Â�MW�Λ~�� ���`�6C�=�_-�,qUK��C%'�S�L��=�=o>��Xs��b,�r�hm�P�\.�G/��a��wٯ��o���8���U5������P���j�|EG�en<Z�_����Ϛrx�!_K"�=l�#f�j�p�����3>G0-EroM�ԫx?�ۼ7��7{J
/��c�w�I9��oDM�ò��' |}5�g�����/+�}��@@���og`�B�Z����y`�ux�	��8������'����ș4�n��}x�?�8h#^���O�	����2��U��8:��Ϣ�����}L��Il���=�ZV\�p_��HoJS�%��[A�W���u��l�x��?�d ~K��^����-ͱ�6#sc4�}tr����^���;>s~��EMo���f�d`���)��L���A�"�xm�L���VUΝ6L�_ӻA�{�7o�[��u���a ��-�������ØS$�I��ΐ����E����Lc{��÷�ˇ�;e���&�m�gl� &D��R�.�|�H3;�6Ĥ)�8�ah��V̲0[��.���ܒ�_����p�"�E���ge@�[d���f���>!�����+�h�,���&@4��B��/�
�>)������
I��|�cH	��Tx��^Ѿ#�S�뻾!�2JV�q4�����cPeϳ�vx�\�qI�U�3�U��ĽR3�v���a��ܨ㕭�}	��њխ?�.\��E�7>?MÄ���q���
4���	�=@�}Gu��1�x9�݂ ����9It�u�=/�-����C�i�!n��!�u�R�le�k��R����?V�۵�<�X��Ī3���s4��Z�8[ֵ�u�6"븞ܣ�M$H����(pY�U*O�D0��U��Ѡ!m����R�(�K[:_��T>/�܁4~�$�(��PW��)JO�=�H/�,��`�O����0�7�qS��ҡ��c�Y���������E#]'���+�KtK�$�)2��z�-�F['D��M�|~��)��wh�B2��8Wg��,P�����H8��i�L@c���!�Mk�aeU�vM�ݨ�F ��%�R�_��9�+W��Vxg
�K⥬�r���eW�|���6�g������`+�;�X��[��"Tk�jk�<�E���^�י� gfwu�������~�y�	ݕ\��+�:���d<�N.�����w���u�H�,3�����^XG�Z�d,���K��T���]�3��<��i��tȋ"����p��UI-S�2|�+�l内kt4�{��+J�D�,���{���4F4�Z�'b�.N�����߹������*wT7����}�Bzq���⻺1��Җ�S_0T8_�4�b�����Қ����w��7�w�,��!7���1e�� /[�Ue��J���d�"��%���W=#O$���#ٜKC���J���`��^�N)�ZܖX�Mz^W�[�k�χ�YI�?����0��S��/���TO�Z=�k���f��':W�@��Όo�(P˻	HO9O�R�����ؗs7�ߴ�!#��PT%/7�(� ��������L���,�W��^&������x2B7��"7�O]����-��hh?Љ�݅��0�\��5s�$!���"{w,�
������ 9]�/B����{H��k��o�l$7���)cU�f.0P+ �1�Z�K�]�O
�Nǜ�Y�y�vy�����j�}�(�jW��k�Z���<ݹm���x*�t�8'#�e�"-5����H:+.� uqa�ѫ��_z9xtƵܹ�Բ\
*i��2sc�^��_��2��p�����^t����J,5��m��� �s1�o�g�EuՖ�;�!�xel���zR�񹨎g"5�K�3ɻ	:ޟ%ڭɛx)����i ����Xp@LĒ)\�:���tժ������KJ����������������1|�� �Α���\@��"�b�;��-���Q��j�#���o��r)l��^& '�ƿw��mh�t�UJ����Y���u����f�|�?�Ȗ$�&��ʥcQ)����*W�����MWPXEdI7m�*=����Wq����B���l[A�3Y"�\?����2;��(���S��U0v���r��`���F��S�:���dA��Ka\���X�:��I��9P�EX3����Ջ�prm>�f�P�3���5R�:K����J&ͯ/�c��d���jX�!M:�[$6bi��5��
z�|��^���.<SFv�/�p�����`��?����%�j#5u�9��\�]7Q��oሩ����8�&t;/!�-�c���w�bh��Z�X�O0xV[uձ�c4�Jn��=k)ST�7�51�<����v��Y������Rq����?;\�\�y�nmw$*��'�/�#�g|O���Q�!ì�����Ҏ��0���i�I�"
��Ah+
z�;1x �Yg�o݌�ڬmoꡘo�i��{Tk}^��)�VR���Rg&�ڃ�����u��.&Z�?os�~jG bP~?_a���I۩L>w���j��O/P��C'�� ?r�����%7��-m�T�1�:�Ac�n;��	�]JG3���u�(Y�#V�`q�9@���fU1\�g:�t�'����E&yb!ۼg�y�����ɡ�����+�����V�ށ?R�ۜ$p�ln�/W�I���}�<�A�*�PR(`���P�uAl8�� g�r<-1��g��h�놈I-u���xX���\c.C|����;�5��{���ф�ӕ���Uy����m�.D����kRr�ܐ���Ǡ���)�F *I��
,0į�>��K�ɦ��\ѷ��d�(��*�������+|̔��.8�Y1N|/���d����UUOEfq�
 A�06��;�E�u�4���"����k��Q�N�����&>�@��9�
���'�1��)���+�B]\��̐7��%��J�^�'<I�<Ղ� �����D�5��}�*R˯]p����TQ���h)'8Ŧ�7��d.����ZB��7��S�����F^�8bn,W����'�w]�� ��[�4OQ4�#�;���,5�:Xy�b~�'򙸵���e��F��U��U	��ob!ц�g֩Y�|��h_��:�DOi��^���9o2���(z��vk���M�_�?{9߭c^=v�f�`��8dKQ���;���H�텄G���(c<���7~HkV�`m��"I�O�:7>
���}�[�KC��K��QH���ݐ$H��O���J������Be����/��k�L�LXn�0rn0q�fr��NU&��YIİ�.�1IF�9�1��Wݖ���HH�h