��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-}�&N��<a�6H�w�#�s~��a�q����w�;�4�ap�Y�By	��k�&IoxYj� #R��°tl��3����2�Yl�<S��':��K�����e8��n���`�=F?�w��	�k	h���d�ue	0�n�{�O0Bm�����ƿ�f#�e^�|�m�5n�w#��G�QuIXJ��� s���Q&�S��?<m�a��Q�!�ș貧�����|mKDt�1T!G�)�W#>��M���:��r��z|t�G�r!7�/�VK�H� �Ұ騴���}�~�!.4���O⍂�|�':-Q�F��@������N�W��Y@�H�+�E|��8$B�-��f|�Aٷ�:�p�`>�c�4�3.ţ���ꇃ�8��>�\��+W2ݜ{���Yit0�Pc;۾Ʊi��獲�j�oD��qa&��T6����^)�
YC��*X�'dC�}�����0�D�﫣�\U�2ͮ�K�z0�LD�$�|�@�֗^������	};ݍ�m�3ɪ�4po����i�2)�^YK���$9�~�S�c���J5W��Q��]�hw�܆�-)=�x���ű�)�[�^���ֹYtk�g2ywz��1����#�b�al�DZ�/{ho_��^b���ǒ�e�]�=Y-��偆Vb������n�@ j�����$ZF�6��(����z�c2U2XHw�v$V!�nڷ���V<m�,+�P!(w���'Z��o�5�]��j�CR������M��eB��X�`��ϼ(�O�̊��6�FW!�	y0�=1��wǖ��)|)*��;M�W��͈�G=}N�ʊ>�t� 0�$$0AݖO���Pē�đi�m�̺�2�{��o wFM��F�]�K�9��
B#{���g�!�G�	='��#E�.�,���B��v���/Q�P�NB6�9d�H����Iʵ�UN#����)H�s�&{b�*wU��YC�4	��qJ�n��� �f�9�3��	�Z'����
�>&�`��f����A8B�]�?��~����2v:L��J	��:5�������$Ot�<^2�jY1�?Z�v;�a5��kYžU�mU�M�a���;�xC�!�E亶Һ0�ecaV�n�*.���U���C���tXw�dZʎ�|�uC�*!�,���*�2դ�룣|_˅fٺ3����-�v��.&�[^�q����@b��6�PoJ҇��E}?�$Uj���9�Nfʦ�y{�Ez��#��f�v�Y��zv�t-��Y������|0	��m�6���;��|��/$*ۋP�S3bi�H��9Y \I�Ћj�Ql������@p��J�b)�
�שoTn�������ȿk`u��s1ݬ�>� r1ܫ��
N�5~�Ȋ�/�:mD2�Ur���5BEy֩I�sCU�޽4��E�`��E����Di���8�"���O-JC��v��LG��Z���q�'�y��0�� ���r��۽wo�գ^~dyB�!�s��t���_2ۣ֬�uL<ѯ*LSŉZ��|of�T�AlG~1���U,NP�Q�5�j^c�Z�(w6#��3�����?�w
���7%���y!U����O�O��|�ּͯ?\�����#2`��6b7���#E���N맔�h �=���d	Q{��6 �o#���fa��2���칑�L�[�컔��f��ޒ��y�,!��d��h���^����K䭊��d2G��Uc��6\�{;O(��SX"��R�^��zt�����i�i����C��1X^
��&�b��X��6��i"�7�ę�U]�[;3��U=K���W�����m<�p�w�\�ύ�������'�`Tt�%H+�H�.ƌ��f��� S=e����"�~���kℷ@���?�0�~#���g��3h�q���Ǝ�yX<-�-�G�fY&�0&����i_�������*7%k��qO�β�| �4",�����͕Q�}��Z��bqh��z���-�i�׿��82w��[p���X�j]ϖh�����C��#� h�