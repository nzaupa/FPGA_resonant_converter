��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l��ӡ;h�>�C�0��-#R�&�`8��2�_E��6�kI�n[�{e傭q�wҴ� u�j;hKb�>�$'���a�t�(�T|�qNW ��J쭓4�[4��V���P��̒�zs��3����������>�ʹCƧ���b64�E�Ӛ���܆���(�K&o4X[�T�@Qh���C�2�hӅh�B��!)�]˃�y�>�E��):2��¨�r_���8�����-��Ĭw�<��=� �r���*�'�JC�#�����KFGui�6��MU�-��ğP�y�/dQ���;�o�dGm�iw%�����7����y���x�ج�j��ĉ����9�������������j�y/�H�tr�(V�=0�[�?A����#��]i� C�-�}?���Q��Bc���y�����cP�������@�E&&�:��'�|�$A6�]`�8�_��nG��w�1+��M���L���E�_�����2�ҥ�w7�9�f�ec���B���PT�]��+�3��ըW�x��^0�	���QXH���������	��c׉���{'.
Q�y��-5R�?Ǽ�hG曝����H��ȽѴ�>4mX�#_{�*n��?(Hȭ��a�����7��ۑ��S�ĕ��&}I���M�%X���9�2dڹ�)/�"H)� ��5K�HH5to�����m���Nb�� �߂ry���Aʝ�n�)�<nUC�(�;��OJ}�@O��oe�l��+��'18�C����3GR9�1�N9��h<�֔��	O��H6��&��3�7x�����%��tT3hզ�c3��V���:�����
�Y~�l�A�P�o��%o՛��We�Wo��lU6�Fx�_�96�j ��D�Z�#Ɵ�q����6��t�P�A\���L�6`��%0�!�-��Z�dv���K�2H�z�P��;�і$Y�ZF��FOǇE�$����k�L�"��]\��'�ڬ�z�u		j=�Hl;��XWr�K�q��ck̢$�����쵈�=v�7�v���[|�6�w�F�	e����\��a�&��:&-��@�� �<�/���\�����'���9և���E���`�֓� ���Mؤt���׬}���~5��=u���*��I��E<%�/������+��Q5ɑ���m������S��hi@WJ-��/���{��Ce3Sf�A!���4�ݷ��M�������y��͛}��bs�\�h�,�ͺ.{��h�a6�q���at�̒�B&�5�z����h���+���C���c��( 0Z|E��6mb��7����k���B�2��� H/DG��, ExР)�8�^��n2�$Ms%�+P�c?�o0op����W�uv�[��h�d6������~������}oqT������"������#"�v�a�U(�5e�����R0Sr
���g��Ê7���E޳����dZ7�h�$N,6�t6!��龦0ƨ���ʘf����?��W,i�,��o�nw��m�TK���|G�J�荏`h9D�y1��lҒ&-U�̊�P+��WJD�jp�� 8A��.(���)d�%5��_�J����V��q�6R30�U��0��fY�P��3k���ӟ\��*Dr�+��y$����ɯV�f8����ȇ��V��E�����O��}$��e�UL���'a���l7�''?T����#��@��+Mv��غF��N֔��Kڍ��,tv�Z���WW=�t���=�ۑ��_ܱLw3K�6]|a�]��jT�EE*$d'V��/��g��w�*�X�J�6�$��,����	
�ay��e��Q�A���=����z�6]�;�&�?�rR�߀�g�L�$6`v/�%��X��,2��eLZ��kA�3`l����r�>uI��	�IC����[��g����=݇��聖+R��M9�	(<���ܪ�+CC�(~��\��7�q
ɋ��A��%3��K�H:�m��{j<͍
��W�?1�&B�9W�[v�)����4���3�+���z+k���<���`%���E�&@�sל2n�'��lF����E�i����<��(��&�Α��/*1�[��������.
������F�X�t�z�!�+���_���@��|5ṕE��<�g�u=MG0�g~�l�kZ:��>YuJ�	�� !C8%�r����E8{���3�Kwn�2�M�*�2p3���]�p��	pL�{AC�`C��=5!�3wQ��;�W9x3;nX �l�8�ǁ��!����2���§���h� ����`�@MF��9Ǭ`�;$wnو��8e'#��"c/��j)�1�H�E"1S�����˾�����iF���5���<������bd{�^ؔy���̗(zǷ���	�>���n��*g9nb��# E}�:f�!�F�G���cs/�#Z��E���G��;������2�$T~�!%j5z�`r�TI^'��cG�W)�M�g������5ǒ�u�g0:&���ȫI`}��f@
ǈ;���ޜ=�h��f׿�V*o�N��ʵ��L����4股�����ѧ"m�_c_��E�mh��C����V��.�|z��R�4bup��}���%����}.y��S�_+�
�ĥ�<2	��h����_�p��EVVl�Ѡ�߭|�Œ�v�Q���Vu~�ɞx�|q��Aw�Q�< �$`���ušK7�d�SB�����d�]6�/����$�H�u�+پ*��k�������*��"���abc1��͕�o�S����p����(��%ZpUJ�\g�L0	�e�HQ��Zt/��h�%2}A����U����t�a��A���2!����z���^v�ܯ��`ekmZ�p@�&��rmP�P���о".�_�x�q�'7$}ۇP����a�h�p�I��XJ��e�󩥎:m������V�|,W^����S:R� �cO�NW�<)�!�B�]@�=K��b*)��	W�D�?�㍖�&�ߋI6�N>�:{|fn]樉7��^!1"�`*Z�)1�A(�y��̞!��<���q=Mx$�ǻlp)���"#�ͣ?�[Ғ?;�w@��~;������9����3�+c�
c�^�����������^���B��br��Fc�s��v#d�{�k')zo��Ӫk�19c!�)d�r��W#����*�h%�U��`
\po���N�FpZ�zF���O�^�=lװ�V�ՉMy�nF�@����@�׷LS�ұ�6��~�n#�*0����D���X�pJtnC�_�tУ��w,��w��(;Z�w�/qj���ǿ���g9w�g=�V
ͧ��x͂
Ut`s�$��{S���������]mv�e���v
���<Y��f�7��4)HS��
���ً�(@�S!��k9cw\�[���j�)���m�t��FO������lzV;x�=��F���� �����S`��+մ2��i'nw<'�|M�xԦ]����L9G��c��3�[UlH��9�>@(�q����A��2(��&��&�FU���+�}�����W�'���i����>�wC�˶&3�c�(��?�!"�Q/e�!��=l,ھD9Z�{�W<C�d����d�?
�4�{N��|��ķ2a)�x�j��Y�6��C�r��WY�wz#��uo����&꩓n�Z��bl#��i�R�$�}x���}wXR��H���kQ�+�a����e�JG�0F�i�m�ok����ҏ�i�z�ק§�}\�'^f�;"�K�ϕq�!A��,��j��\"/Ma��kҤg  �)��Eb�A2([c�ݵ�N2B�=����s�QQL}�"M2���NFq{�seaVGz��"�Ԟ��]��1c��d�.��&j�#��	�O#^٘I`F[�Р����e�p������>��B�6�6�B��O�`��}V��/+�������Q���T]M[,KC�-�V�D�;JD����Ps7R�>
K���u��?β��2T��2�� ��ƘO�vF�b�1-�YX%��n�h��n�1��e��"�K�s���� �3�'ַ��0���^��׻P�A�CT[�c�M��@�����NLԥ��˯fQۖw��ą�Ґ�.�ŀm-Ud$+{�%GZ������V�
�/���4���n-,.M�n�¨T���>�6h/�\��55���)���� �`9��U�U������=͕%|9�z w,v�*�՘��r�!���v��a9�K�B\�76`��ؐ�j��?��g޲?�6KV}9�.ˑ�Fa����;�j'�z�G~bX'�6aR�������ɝ�������$o0�M��#��A7��ן+l-,C��F7f(�ݾB��z�"�yg���ޡ��K5����zd�a�>���(�y ����T6�h��8<��@���G�л7�ZO�}V�Luo���y�	Lj~@�
/tW-����Bg���v��VTB��0�X��aH�z<�vV\.u��˞���Օ�sHC9_B&ˬ���֟���]½�<�|�_F�Q쩅b����7�My,)�f,�ט%6��u&c�Sq��������d^Ek���Ń�ȶ�_��"��d�,�_�i�����f����%َ.��6����p��I���ʇ*�c�YC�$n�g�6�F?��"hҦ��p�'⪫h�e��ҹ"_Cs���P^�I:���nn�Ӿ�=��X�����Ln��
��e#���'��x��G	�qUّydxVo�Oɓ�Bd��/�r�Y�P;Q==������r�>=?sM�3n�J�ZgZ��̋���U��S��n�ߍ�9	>jxQ;r�Cd�������7:��ɸ��q��^�S�;X�+�}Ǭ��VV0�&�61O��9�k�#��u���	Ft�>~*Vk0�[)���?*R��=�+�)szW��ђ�>�SD�a{�L�nC�\AY]̣�ء�4ϐ�#o󤋌��è���'�R%����3�7�}]���
p�T5;ՓNS�/�~DP�gL(e4#+B_0w��t�}ǥ<�D���T�G)�ٴ�|��#$Ӆ���J�fW[q���B��?��x��PG��Ʃ&B	�OI��2���x@X��N�bG�5��/ր'�,�j��1W��p�BtB���Mr����k�.]t|�,v��$��#�u"&ء��^U�)2ٯ��ld�X*J4�d�J�&�T?�2nCp~����7
3k���R��ǜےJ�"a�&�s�c�R�(I!��m�oɒM�s��Jo !�� 4��m�ΩT˞όi��,��=��<��=
.��l
S���)!��0�=���Y1�
Q5�ԑ%�� ��}I�L�'�*���8�_Ӳ� r$%l^1yOX�������@�CsB��;Y�2�u���\^�z4���5�٫� O�35>8�X\��w��3�H* ��B�$=}Z��
)(��
Լ��OeR�Kc<�J���W�Yw��\9��4�8�ɒ�7��=�Q�F���:�W!��g��g,eę��n�5T�i9'��:���v�b��@Sq�զϨn�~����� �:g$3��' FR� Q(��t؀8�������Ў�{�k���0ÐE�X�(s����г�7V�7&�3�&�q�t��y���%�i$e|9�����EX,�?���v�3ׁN�\ޏH'}!�{�g� �vg.�UL�n�{`���=��#i�ׇ��cC���,�d���|Z*qD)	��Ё�'��gi;��3ꨓ:
�B���l��u?�۵�P�VD��J.�
��aW��.Z�]��	�����'-
��ơS���:'X���Ϻ�ػ�-����Dh4v` ���%Ba��k��TimUߺ^�S�� t؉-~]9\��7 K�f�����]�W�����z���i׵pu���f�x����KF�e��X7�\�Zt��S=E^!tR��������QvdB{�^k��"��"��*H,�M'�<4�^J�@�G�ޢV0ӚiO�p�6	P�=tVsyu�"z&�D��U�y�f@����6����d���QL�96\�N7�_�l�sf����x�z�ښ4�a����2�܉p~�n�̂�%�E�8d^/r������|����Վ�% uyS�b���.$Nh���w\+#X��u_�/cg�i��TO�CK�?�?:��Ö��Yc�I�&�N�؈��hx�%�
�P��т���w�?�~A&���B�K| F�$,�&��K��H�K�K�iG�'��p��(����U@�l�(e����	:�4�a��K!�	٘=�楽�4�Y^b���n)(�DEXM��n yp�}���E�O��
(�T��R�o �c�	�%�v��!S،���0�x�4�&eT��򣚠�"�|#�i�nUɭ��jb���-�zx��RE]^����6wj��s���$<��.(p��{
�P���JU�ȧ��Fј�_�����w+���E��f�{;�x���d��3�b�Z�,b,�4ͥ4�������
Z�Xb��������6�Dշ��>���$,��k"�!�D'QkE:}`MX8Q��R��΋y�O����OE]g�DR	A-�wCocyC)�gػB���P��ͬ��U2�{j�	�zp�W� �h���e_�a>��E�;*�	��T�Y+j_q�sN����s��-����?()Bo�0�[�����\���a��$ad���xj=8�rΣ2�'�^��\��i����)B�=�o�_��z4�w�;q��_7��C�iD�%�p�,�*1�{��Ék+�.�&
煆OT�6��c]��i:S'��"���T*�1h�!��['���E�Q9�~��ŗ���'[�~�$Y��T]4�4����%(�	�$�V/��л-�j��\ `Y�Q���I�ljȰ0Y� �����|"_VU.�^O��歾�ER&E�P�ePw�`>��q/R	* 5�b���+�F����Ԍ����Xe��[t�G�f�6��U_���u~ѵ�g�� [�"60����[9�R����ӏ���C�
u�0�f�Jd!��=(�~Ko�U|���E�`�t�IlH�n���vT�H1��١�����{.ˈ'����{ݬ4�0�h7*ٵ,�����H�PoQxjI��h0&�����Gd${]��j
j�Cڗ�,d4_�V�v]��0J�2�h�tX˻��VZ�F�����l^��P�~�:��u~Mt��AKW��'�9�e��8_���lF�KC� ���t��iJ �,{�)��lM�%S*���'��Uֳ�v2�?����Z�i*�Y:sbm.Y���wf��q���*`��`XțB1