��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_���x�Ay��[=i�,E�aiF6
��>g��,��ψ�~	�l)����V
�jh�F{�iOI�:+=���l�P�2h��+Zﱻ������L�����K?�ct�����Gέ
��.T�|\*`��V��"�+ZP����7�"ʜ1_� �,��Rz��5V�N	�(6l5���7'�y�(g�d����}����W}�3�vz/��-�YUEBƌ�R��}MV�N`Ӫ^V��e]�>���E�R��:�Vw��Y�$�zv��f��u�_p�1�xc��4z�fw�{-��.cf�%�\��j���@�����*o N��a�b�$z������eT�����S��wǆ�9�!;����.����RV�o����;�C㗊��b"Of��He���[p\��kc� �g7g&2�+���&Kܚ�U���Na�ց���y��~��_��Qs��e���Q����(����\A�C���@�xq�����[+ W@ph@�"��͙�5DY�D$�i���U����� ��ߟ6ZC��s����� ���
h)�zw��Q9'ޓ���%�!M�o�F��#~Qo�{�Y�4���&��`��r�c�y_gܚ)��R}3�<�	O�� �#����q���ӷA[�B�&�1���<��ㆅ�BC��λM��9���8�*c����\��[:�K8�of�19p2S\?�[B���
q�r]gY��Y%�wV�����+���&]���t$3��Ͳi����Zn$^��sq>ɧcc{-73���[��q��v��JZ���r�荿�J�j ˍ�ɼ�kH�s(K�o��j֔���x�Qhz�d60@�@�C�UZME�g
4b���o��,��K��L�H��aZ��H�E�d�/�c��&������P��Mԣ޶W���6h���.vf�$u	tA}���A��,	�F1�ֶ5w)��KK���Ry ��eɄ^��²��/�&�#��$i�@�F8���w�v���),�,�|̈́
���%�5�E٠gG�����01{�����\��_A�-�-��)�C[�nĝj�$e�_6r%mvT|P�J��(����y��U���&�eaD������f�3���~�����vÂ�5e$;�n�K�FOEqT��Wf�m���Kk��4T���sR�����d��A+ ��|Ӯ���Ӭ���*A���uu���鿑�E�])7Z���ǥf�8q�9虥4��U��.�{�E�9,}�,�Y�1�B�d�ټ�����l�Y�����ؽ���B��6���̾�B��[um� p[�]'�}r�̰QH��i�l �*���J����v�[��L�y��S̱C:H(�����,�w�z8Y��Q�Tj��[�b�f�/�̙����G�
o�`���$�Lġ.���,�i�N|?��9, �;��V��s�]�Ӭ��G-N�櫈8���&ڥ�5�`�+����Li�Q�a��]�:A�d�n%Ŕz
�����G���r͸�Q:��^�ʧ[�z`1(��ek�;�w^��]�,�I�O���a��Ƿ��6sD�� �a�^��13���E�T>�;��òװs6?�.?�ӚZuw�%�;S��{����R�.6z���gHӿW������f��ZPx��(g���f�BLn�2�S{ki4{�V���=lP��
ש��-R���V��b�⎮>�x�]��v����$��(&��c;�/R�A��s��crM�B��$@a���6�s�5�l{�|��9;L!~�W�|�u���/To�_-Ch�s�Nh�h�H�Q����8����'����n�N�z_x�gO��d���"�c��)����,ěc���{$� Qzn�j;\+\6��15�:�G���\d,%s�*s���2H�y�fxĒ��ͨ��'Y�Xn():A�h�8�g�P �c/d�t	�0�ήձ�\�"ԩ��L�/��%��t����wT��K,,7�z8$� �dPe}л4�%�RI���+q�}�n�Q����	hQ��tsլ�R_�|{�»��݃��|��"�ĥӤ��Xx��g��	^��~��i�j����|W�|��9��ϵ5�41]8��5�kS
*4��<��d�>�����D�%�F�x:�r��n	҉�A��[-����B� ��Y�MA��:(5�Q�/�C��;�^��=�dy
P�[�h��vJę��(���d��C(����aJ"�L�<.?l����WG��u0b�]! Y�H�p8����0p$#��A�2�)�\�3��f�HaT�`
����(�5�E"�X�C!�r��eK�G��J��Y��~����x�O�|k�a�@�q$kչ]/�>����#�U�rM���ĥ�_5����u���s�~��F��tq��6%(# ����w���-�v����F��o�-B����Cr�F���痙�[8�q�k��sf�~q�A֦"�-i�>&�>w �E�I�(�ݏ�ީ�<���N����O��k}�bo8��P�Sl^a8���o=��aj8���"��>���b�ʑՂ2E��a��r|���8��J��fΦ���`\ӈl5�\��Qo��L�1)���dǄ�v���[D=)A�z�qO&C�k�?k�'�� p�lͷWF���V�uͶmC��FKL	\x��n��R�ѳb�K�i&`���)��.n�"}<���x�"J����qN��x�;�+)`[���m�:˭��,E]�A�zҜþ\�|�ס���v�PAp�%0�[:]��D��=fة3�����l�P��\�pOG3H<5b��MV��q-��&i/�%�H���.(c�~�_�ȻB�3G!>�$�4�I�F�!�[<CX��_n��T�d�W��}��h�$g	��:B��q:K�O��\w����޸�ۄC�������gv��k����ܺ�?A���Y�9�*��_�XX�ȕU��9���Xn��GQ �J��0�����>����:l��PaX2^	z�1*h0�B�u�u8�*F�h�9��`����B�i����'���Z�Q��z������91�AoJ5,�颕�Mk���q��[��ٺ��맓 	��@{1nm:��B�E�u_:;Up�w�~���}Vvq�HK%3�:RL�{	JCp��)���a�iP�*�x��=D�M�!�Af�~�R?T��"(��Ѐl�%���A�㫔@%k�Y�;�#�j�O�j�t��"^���-Y<jݳ~��锅��7��z_p$3A��B�sڊ��``tt=1�-�ijK�V���ߧ.&~�9��aWC�,�o[ U6�-�o:��ZP� ȣ��I}\��w���FKBx�zF�oj�S(������� ��
Z����*{�K�@�m�	���k��}ZS�4��v4�q"j�*Y�Ќc+,q� ����A�����=:�W�q��G�DZ���c�{W$�;߼�w�kn�lf�	�_w���duf�n��֓F��;�r�^6ߥ�W)1!�h|��G��y�/=���v�����ћPro�d�#Q�� n􁕠�� ����3��������wZ���w��Q�9Q�&])^;�sB`�C{��	�N��jӦ�P4��c��@0�)����pY�&��=E:Q���0���KAR���-�[q�)�#�*i��.V�N'����!�B�
�*����xN��\J�h!�"ۯ�^yu�]IzE0�b~%�/L����rUG�����=���qDdw%!�S'��� �i�U\4]-��!� ��i1�`�����	Eo������lc�R��:U���`]#�9����D���Q�}����t�/c$F���F�7D.�tArk�Q��HxX��+6}C}��b$��,{0,��~8�79@����
�����D �=j6�t����/�I0H�I�������A9t6A��Л�QG3�`٬��w�A���3;A�|_z)�<�]�$��b�A�s�G<�~��إ����E!|I� eը� :�-c�~��N$1%0��^�Rf�v|�P�1�=�R���~��vtbwYA<��l�������zJ���N�.����%$��T`Q�P-肱���jܴ��4��G�*(��[29w�</[�1�殫y�AH���#�L<�X �Ly^GUʆ��F��N�x��
�$+����5�zoҊ��b~�(�7}�S4�cO���1��MF�%a9m���$X�g����M��h�Ԇ1KcK܂tD��a��=���G[U�n�������5FC+t?\dڊ��I����΢�p�
��'äsaw4Ѫ���8	����[�y�%���3μ5�K�ù����s��?Ӫ�.����(�~>;�R��co�<�S=�B�H&��Z�X�Z���a��)�:s&���It���[퇘-#��b���>��|cT8T�e_�>Ѿl���-��`��ld�9�W�D�9b<[�5fя�n<>*��/\���/wA�{ 젠�Fcf�������z�<`���
�Bjņ��Ҩ� f���M�e�\!��B~�K���}�/>�p��;?
���7�[Ko?
���҄������	�S���I'bɥ�3���~P�H��!X/��Vؤ	������@��DN�H&%���_<�Je�7�8QK#�m ��D�As�������̭�
����Azu�B�ӡr�.b ���%d�Kʜu)����W`�������;���1X�XJ�M��2��7���d��"��_ͯ^c�Ft�i��tVQ.|;��n��'�ҿn-{��q�g/�P���.�go�<� ]_����������6��&����M2&���_?�����)%i�1��F^�I '�Y�01M5-�~�(ٳ`K�E+�l�p�H鳮7�!̴����滹3p�h��)�����р�
 C�e:7ݢ��󯴖Fp��.�p�0��j5� ��K'����EяO"�����i-�֙��X�>d���'"��D���Ϟtk�����S���72"�6mO�C�K�{���s��W���f���4
yO�S;v�
�Udf�lΘ�3Z���Ku}�}�3���RN
_Ȟ3�.1�]��v�& ��)������#�5q�B٤Y�:9�F���P.��{x��Ty�鋹�| ����m�g����v��!nI2l�>a�i�;�zw�Sj��,�,<z��l>����-b�I��;�g�׫�#��Ƿy.M����~�cj1��5�E���V�[��b������mK;T��nDt����3����&2~G�5|�q�Hu|Q1�ƪ"gr�3�Oܹ���c4�j[�\�a����^�j�&}�Z�p�����y��VA#����j�iB��a1��ف6�2u�M��`_����ᨃq� ��v�GB6�3˧T�� �{o����5QoR�ϼ�5�L���י�r4�Р��͠��I�!Ud���8��rY� lTI�^�(D�A#9?�g{#�[Ԭw�.g_�$���fd$lW��%Q����P��
_è�x���� ?�	�1������22H��U]*"�>]�Qڵ���y;-Ui�%&jq�U�v��n��"���x�Gy��'H/�p��%�@���0���J��Vm��g�~��� ,��chM��Z��Ӫ1�G�E���A��Ϊ���������-
���}φ�z���T�f�\p��<�P\�P|�G�d��Ѧ0,Q���Y\��Z�6�Z7m����9��X�N�緙M�x��]�^L#��Y;�k꩜�x[g�c�~*�����IY���q�Z�I�Ki�[@���IM��<�K|�iV�@�5K�KX�84}�T;���zWe�k���vI��$�B"|Px��X�8���h��}�b)aI��"3O�2��^#~��b�(�I�b\w}����n�.r	��C�N��M�;6,�9����Aw��|��b8���@*����(��}����a�mR�r7o�qH��
<�����&�s�.�Cl4���9�W��:N��T+�(��	9�n5R��c!q^�f4)ƠJ$c��ј����?�v2����u��&]?p�u���ewa�ӳ�d���-2'kHX�h"o��<G���lpBL�v��������r��8�V1gWх$�Ǉ愍 �|-A��H��	�(��`��4 �b9I�<[�Y��V������	�aR�
$ڝ������#�@aB��r����)�w���)��a5c4}�Kat.I�NؙX(sz+���e���n�u�|:��^����D��Ju����3�3kt�fi���D8�����3��M�N��n6Լo�@�洂(m�����!t�~�dCS�ck=uco�:z�'�CV:��h��U�t�ikk�K5G~2\ �bk�-�CG�Պ�g����I�΢ ��|��u����5y7Y�cഈ~k�� ��\�fܕ�D��Qv@b�u�3Te(�RM}DF"�G+�y[U������C0�Ow�O�N(Ha�*_��	]�Q��tԺ�4�ֺ#�$ ��֩�ni�6��4����9��k�k�6��ʍ��{��G0E��߫�iHy��I��S���:Ȳ&�E��t�y���O.���r��x�8�P�=��8K���P+�?/)X���F�A�;�d�U)��L���0+�c�C���~:[�W�R���<����>��?%(��?��.ld0��Y�����}���}@X8A�vA�O�@.Gv&6�M�4�N��UަTy"=�R�4���)�=M� sp���zx��k/H~O��$�A��E=�U>F'S��t���gM)C�V�1�_��Ѫ\@��M������%��UX���B�.�7B��0�'��p�o쏀�lU�}�ƺ����K�=�h�2�N�� :��-H� sW�'^����8g�,��R8�$^v��b��?n���&�C�=m]E�I�9#��q>b3?��Q2��e"��ə��-wF��حw� *�s)C �Cӕ��-�9� �����	flg=��L���Ae�[4�Ƚ�N�n\؏J���Aܪ #�}v�P�����W,���F{�2�����9Qԡ��SD��ջ�~�'(�R>�ljM@,?*?4a�m�e�2���+^�؀��~䗱�{�%`0��+k�����,��� ����A$>j}�e�	O�/�~i���ĭ��S����9�߯�#�GO��Z���:��9��W!���)�	��f0��Q�#N�c��7��~y���L���	-�Jy���7x��ۈ��!�8�f�N��.�q��exR�r~&\/}ȹ�����EL�{e��D�[�r��ny�>�)Rv]�S����L���v-�Х�����Q��9���0!_��&i���)�Y��64�e�">�VP�m��l�#�o��E?�����aA��{���[���傣�NTeg��ji���(���ʐ��y�(Dj��I�Ca6��*��nu�)uj�j8�\�]ý Da
[���<�>�w8s�o7N�0���\x
�מ7��fI��ϠY�P��#-DF�t{a�j��]d?��A����e�b\���n�@!�S`����U�f�GK�3�6�N����Oy��U�o�����5�8ƓOz���v��~��=���c:c�e�{@��ڼ��>�nƢ��.��gS�-�2.�0��,�F�>�nɾ��ӻ �TaB�&���
ʊz�|�jl�����ݤ�^D^Tk�Za�e�˭�W� `5�磏�IW�N5�� /H#�@:Y�~�YL�����ý���Ns����?����JZvڥE���B�L��?�w��%w.��O�����yE4���I��7�Oi�j�#���!av=E�$���{N��i�{��Vks�M����̈́�<ܪ���$���D=��󌃷V��#��N�VB0zq"3��!��L'�"e��-��ce���7��kt����<b��yek��5�Zb�v��ǣ�*��I�xπ��6:4L+��y�{c#t�@� �,�Iո�s%m�K98(�R����b����t?�G�Rlj$�����:;��C�o.��X���L~w�O����Eu�Ο	$QR(���y���p��@?�c���;��ᳩn�O���C�Y��U�	
j���h�@�2Xu���Q�}ח�̅N�=ųg��dٖ�;T �_)��uiy	+G�<� �u�ߌ�M�q��*���|����'��d��D0�R��m��l�*y���r~� ���	W}"�i#��vU���*����YjX��H%��R��}>���
����-�j���i�y
*ȅ��^��i����y=�'��K5���!��A�p�gy��#>��,�L��qX�O��t;��Q�����n3�`�A�*i�r��W��i�^_��2���
�ogc���e�3�a4(���s�t���_�C����t�Ὦ�?��p�����;@h&�#������������ˆ��-_L ���"���n�y�Zwa������g�A�U�A��(+�k��=@Ph9Ć����Nc$�,��"�/�[^�d�M���S/���<}URf8�+�ec�vj���7�驩�v?�Szt���
R�[�r���.�!�I��XF���)�Q�,��%E�ߴ%�#�ɚH$������14���n�ېa=�����䮕�T�8|�k\?�x�K�P��Vn�F���a�(�1���-��e�vf=36 wj�K Ko?��hR�`1�z��X���m�
���A��=Π���B��� �3j�:���4��YӋ�NqO ��BI�]��L���%>����^F�(f�:E��	�!���&���<�;�Ƿ�'�Y�P��Յ�0���7����6H��1]Y�DV�����ȵ79­W0��+����{=��sKu�����o%��s���}s]a+U�����l��5e��'��������[�U�DX��3nW{,YI�(�:�\+�hM!d_w��O�8�AOr�&�epd)��h3�㢩v�]����hW�o��q,�����v�M�|��yx��V}�$f�΁� �D`�lFE�K�l��h����;ᦦ���,t�g�y�Dd��h�m��}qa��ƅ;>k�9���uU�f��>�r�Ea�x4����1���0+g|XՇ�k_�ќ��j>	����i��rb��ao�	�B�Q1��֍H�D�;�mQ rU���1���2�e4�˥toK��w�慝7��i�0_r麺L�h[^���3OXf��ͅ���m�g�ZWYOãH�
(��$'L��
#�=��7��Y'h��1�6	�T�����m���M,J���M�DI��K/XJ��=�i� ���T�j��j�{ӎ�s>_R�4���c)��7�}�OG�jf����ɐU����e`U��O���ԍ��s8��_����0�������gL��b|p,is�"�"<%M6��3*���}D��6ub�����V�^-Y�D��E�{
���Ã����Ssi]
%D��H.�#1%�<*C�M��y���X����I���:�[7�y�%�y��i�����eC�RY`.o�Tg�T&�p����W�F(o`9d�K/e��S0&����Ã�=4����N窆j��-�G�������T�f^�����P&���m9����e����D�<�j���Aٔ�=��%#��r���H��/IPg�(��8qk�W�e<w�q#"�Ҹ�h����J�<;�g	��R��^��&��o��Euk�Q����,�2)*BO����A�%��=��o�JXc�ouS�L"-!�.*�1[b�8�!A&׍/}��ɎT.O%��=��g�eM�+,$}���	�M�z�H�ǣ!��K��O�y�D['3�-�ꊋ����2}5���Pn<j��
��ĸ�U�d��K��s=.ȼ(���N��N������^ߋR�%{�$x=Lv�P2	�f��5.=�!e�l�J�ª��w��\��;�./��S���)���]�ø'V*�f;��	���r�5:i ؙ'j�x���s�:m�Ϧi�z�3M	�5�b���	E����;w��c>F���Ð��<i��x0�g��sU�][2�U����2n��
���A#[�5���l*u�=Q���]����J��h��+-�l�S�"��yNS���r��g	$(���)�4��=��O�u7s0@�W��\�m��V�r�O�u$�{pĚ��������ˋr�#�E���o�FY�<价�_����@�>��-��=��)2	�$��.��X�\U��A/�������X�C,s][I$�(�Ӝ��C���l0�!؍9��uO ��q1\c �r�ஐ\�*���Q���
$4ON���gu�F�]E�I�~�b�� �k�Qy��u�3#&*�܁��������(�0��hѿ6��"c����Ou6�s���vj2.}P2?�e)�hΜ���J�*�-j�c�)~�Re=�as������k�)T��t�s	����6��b
̳�&�+�Y�3`w�~��Dܹџ��>�4��Lj��-:���\ ���i��`JA+���2�����΋��Ik�`S�h��7�H�k$t��nr�M@�`�"��PxY*��I�����N��������l9�k�!
���6���s�i_u#xD���vD�V\���(�T�(��A*pa;��C|ʇ�8����� Ҋ���O��R2^��=_uQ*�i#h���r1�U�����)�]����j�-蘻O!���Ԁ�Z�\%6J�[��d��vB1z{��]�����p-4�]�a.ߤ�DL yZl�G p>��d�����E:\1h���G.�-�s'��I���]��t�i~�[!Ï�WD�c[�*2�x���H����p�^�|��H8C}���,?q��#�<}Ѱ/������W�l�naS&Q���E�%�kh*��K�Pr�P�!���VƘ�9�O�A��X��z�{G����$#�\/ ∩Q��6U�'i�s���U����A3� �o9��X��+�C���	���M�Оv$��Ǻ;L�nbH�t�@�՝m{|[�2�őC���g吩>1��K^�����K��cY���y s�eK@��B��E�)��c�X뚣�������2XV��>_t�o���t�n|�.No0�(���� X׀E���{�/�����
>YK�杜��
A-l����K࿭y-lq8q��`���q�a�������i���E*�Za�P���d����h����೯��=�����»=G����|�=|�fM�^k��X�@���WB����o	a�!�-��dg��/��p����@}������R,&	D��BiY��Zغn�d�ʫ.��A�D樒м%T��6��0����R	T`��`wz�K��x5D�J��hjԌX3����%��i�*�v�N�FG'�6���8&�@�qC
�߹6v!ie�lw�R��F��2i��1��J2����:�@"I�,ƥd��1�Do�I��T�\VoLZmz��~�6vs�T���3��Ǚ�/�&W�<q|}�V&=��x8Ζ��4�����_�6�WT�,�e�j�������I��=Pn�A��WamY"VԊ���Dۃ<;N�#������\B��@��(&�|�6�4��QA�=����\?�rs1� g�4]LD������(�4k��U}���]F��jI��^�N�*Q�F��$h�%i�0c`�Q�)�g��W���]I�=j�Em����(D����o������ҹXu/���FZU85:�W�D3XF���G�?-aþ�M�R����}Id(t�A&v]�h�2{�a{���[ h͐��`�p�1���@z�}5/i�����b�)h7��L%���OSS�RM���ɮV꿀�̧����m�n�B0it� � �� ��1�K4�/Q=�s�y�m<����D84�ZJp߸���v����P}�Ҙ[���]�������3�G�xq��;��ɩ�nwB�T6�r����%�G�S��S��˴�6/���:�FG�����#ݙC7&�2	�T���Ƒ�¼�P	Pڰ�3��,Ԛ�җ�T�M����5=T�[�ʆ�;�z�rB$�=�&IQw�5[_2٥��`�½'��G��p��+���jw�0w�^0,����֓K�U�������q�#N�-�M��s �zl�cJܥ��ERY�Wy)���F�o����	�Gf���(�#Ƕ¹#�=�ݙW�:�w�#�WŔ�������RH;�kȁ4� � �Fo���"�L׿�|z:�|�n��G�x:|�X��0�2��So�c���L`^��w�r�XIڳ�����1�{����Oiy9���#����0?��W�+4/L*9~JRK�R>"�(�}�낙�ݗ�yB������[��"�74<c��(cL����8g�