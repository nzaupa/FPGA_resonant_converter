��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`wR4Nx�8g�aB��=�@pfp5�I�ߍ ��;� 2_�Y�~�o*�n�o����C/ �ڹ@���xg���rHU�<�R�����k[��8�M��k$ 	�,:�Z�`:�t��%i3���s�8�x&M����^\��.����1I3020�M��K�����xL]���<C����
H�?n��P��S�aM:�)D��� �YZv5��q�E|����N_|��B�q'7c��&t�73 i�}^�N���8%	K#R���@gP�eQ�<Y��7�)��r
�e�0�����YE훓�G���>YV��I�*�����/�D�M��(^o�-ܣ��!qAO�p�̂ՅrIK�c<ɈgG��R�����a�f�F�J0@?��F��/٬ns��f��,\�럷�m}#3��V�����S"��iõ��"�g;��4M��r~uEiƋ,�m��J����}[U�.�B������`8X���:�x#b�̧S��3��N���)���n3�D�\X�����@�?>iأ~)��@�-"\���w�mZ�ۚLj�z�p�B��~�(/�+7Z0����f�tZe!��l��r�{��'�[,r0�ޝcԻŮ�&�<�<�x'�k���N���5	�[A��W��+�A-a.4�x���h�iÛ�%t��������n^�W�_٭��� /) z����-$F2�g,L	���*�[�p���퉆��2 @1B��:��C�zCJ8�C�T�J�����'=Ѭ��6�/c��C�N�%	w�T:�<hboS��i���\�������r����Ko�Byf�;'��opy; �O���_���$��3]�����N����~MR��J�Oer�:�c�m��0jX�Y���%J=�d�b`�l �:�z')1�#w^�lη�M������i����G��b�Jn���nAdU�+�\ŊNp�ڹX�?�D̮!�!G���W8bw�*H�8x��P���yҀ$k�_9G�C�!�]bu鱣C�����^��ۍP�<�:�b��!~+�Q/��`�����X�uF��x���8Y��ٻXv8�i�`_���:�u��k���������e��횆FG�1A��ai�6b�z�7h���9��l���D�f���`��=�WB�g�V;Ӕ���I��7&
h�p�N�P�����5��/Q�9n�T�ȥ�kwj�r��|�q2��)Ll�M
.&d4���<9��ނ�t��hS ;b��&|_���G0���NZ�ȕ���Ó��>�3��KQ(����f�����&���s��Ѿ����O(��S
��=�v5x��<����@������
� j��Y}s��Cnqp%\kcs?˂
m��-C��ws����ۜQz�=��-|y1�������������7�� ̨zs����Sl=z�=r%��¹&h��.�aؼ1�z�\`p��j |��Ys�n/������j⮷�{��o�P+h��9��v�Sqe����	.e�z�����R´��h=���vY.r��cHHI�k5��!>�-2��{y�y�D�0����礐n�:�a��(�� �J
Hڕ�JӁ�c_����X�#�ꊿG5r!�Ǯ �qZO�rLn�-�o�5Yd9
������aAO�;��W����<΢�;��Ǚ�_ƅ�1&��]D����H
�E�X �JE���-�B���Mύ��c$��3��<2����jǊ�.��m�9��u��L%x���F��Ĥu=bĠ{Z,|h0-�T��:�i���'pu��$�{���b�6�͵� ��5�(�t�2�դ��R70oǨۤ�$�:FJ����P��ś3�]�n!L����.��BK�����S��C�p��H���
1\�_�{YGB<T͋~��2���m-�aQ���AO�s�e\h��o��f�`��_^��?��W'[�R���(����;�V%[�u�Ɋ쎋���z6�%Z`úN̺ԪY��z�����x�5fz�Lf`�qf�FRh�%ex�G���l_�B�����%kh�܁����z�o�M��#"�����1�%�?�b����0���ݑ6��gw�]��o�N���@��G���P��4~ر\�m��m?	*��[w Q4�Nւ26-w;^�ѐ`/�b���R�D>�<S󿚄j
��&�4�Tu"��E����X����VX�:4v��
`f���2�	|��1�"�V����J!� �|�IR#���v�Kщ�Q�}�.����ї�&��(�߷�X���AꖐY�apѩ4.$R���S&xq{|��jzⴆ�e۫��@윕������*�.�E��ޖ���D�*���2�J�w��l;��d	�!*Ϲ�.9W���j@@���ɉf�aTޏaq4�|�����%���KKKV�z}���ۙo��"�z��Z�gc�J2�A�0�M�H�o�پȞ2��O��E2 �Љ.�ϼ�1�CN�J&UԩDU�]۞Ȅ��Ĺ�=�<���#��۟�p��!��؉U�Ŏښ�f��0��J�f�Q�^�27;�3Sǒ���2�	��\����&֦��4��b2��o�8�C�Su:��Z�k�j��3Ѹ��C�<[���'�R4ɣ�����v���)�d�ۍ$�4H��b�	�����X����_�45���%�v1��::J|b
ӈ?����P����~HG�����NdI[@����Q$vj��h�.X�|���M��r&K����=�̓������{�h^��Ѽ�{+���|��v���R��6췏�x!,�! wIۖ���Ep��� @��҇�ے�U�'J ƞ�j8nP��[b�0ͦn��w1���,T`}�(��+z{W-as[� �cS��X��j��ׁ4�p��`����q��Ӈ�6h���Nl����d0��!N7��X�A9���D�-�YY�������h1>�$��&�� �L�1��%�F�<���oXu� <���.iBj$li=~�Z@��1	� HP;z��I�1d]�Bz&�}��[��i�G/U�w��/B֥.��nb�jB��nD�C��˼�:��g>�׀L&�\p o3$�!�q����dI�����'��GM�ǌ�^�e�U���ᙾ��z�F���Xe˼��j&�"�x�� �R�N�qiI�͏:G�4Z_�K4G��W�	���9��w�7(���d(����ȝ%ݱ�7j��o˃���˕�4E��~���J�A����G�(a�Xȑ���C�#���y�$/�Σ��a�� -f�
����/�8����.(c���q@r�����f�����e7k�8���^@�`
D|�6[od�T%P�PW������tT�7�x�P����ѽ�n*d'I/���4r2	N��<v%4^{�}� ������{n�e���{'���i;?ɎO�:0ňBU���N�Z�;�6w��ӹH�3���QX~���h\6��Ő� �?=4�k�)�?�:V�-���F*����7ͬ�mQ13�7������O��|_w^��7�(�`��w�LQTt��A�p�����cd��~M�����hBP_�i�zIR�=�����[����}���A:�/~�w�� ^-j�mEkt~ڼX�f^�4����7��.���ަ��I��u�W7��㍒�G}9�*A8+�h��6��>�N����㸛T?nY.���$Z�V��}���#�D6
�Bn�
�xmB�|`�xֆ�Wt?�@�ϳf�>�Gm I�q�M�68	����.��m�h��v�=>g���ˍ>�PV�Z}0f;wz�+.��Q�l�a�,��9ֈ�@�`��?ݤ΢.�@$�}q�$�:���� Cd􈰓����7vwu��_�?t�;�����q/����d��@��Oi�[�gE }�)�<G�E���}�*!���MO?�
�f�ݚ؞Jz���*��GOP���<@ې�ط�ɋXC��S�����Ii���ڌ�+8E .�1��J!B��w¹��^T��=��T����.Fg��A��NA����:l��R��KPl=��FC���q�x��v�pw��v5>f�� {�wT/ap��A�O�:�!��P\���(�A��Ȅw|l5c��8�"�_f���vȞ(��{�t�g��`�l����nO�س��]��}qts!�����57���e�{z���"TW��ri�i�n��i��֣���l��X)Y$��&
���G��yS�"AH|����x_���r�I(�HV�ԗ���ό!C��Jzt|�>%����j���O�AW��_����~[�Z�"��T�:���1q�"�)������ �r,��sI̴�|G�Вe.3KQ���;�E-� ]�&;�3/�_`ά|,�����DE����,z#$M'�kA���%ɻ`a� H�������b�1��Q% g�r�
��wj-_`�w�wn�$�z�
�����b�Pʴq��T���.VZd��&�`-�xN��a�h�☈���X��ȵm�׀9C�EW�P�Hu2��ʗ�͕����|�Ę'oѮL�k��ҋ�b�n� ���*�wL݂Q�41���-[�K�>	�:�Xr���I�5�n�AΈ���5�@���.-aW��-��ժQ��FwS<���g������^9o[�h��p{ܞ+x�lW��V�����Kv��/������̓�M�U�WX�H�M�jY|/��.�1� �s���Bl]ҩ���$��'%�@�+M-ΔQSp�|0/Iz�uYc4z��M��"7��r�O��o�"[,�d��tX�T�I��%�)��'�� O��N�����E26�o�2j���1?qej,��I�`�@ȕ-�AmBm��]�<�����P|���z1x�@*_��nM�����	� �@s��K�,I���t]��`qSո�A���
����`�]0�'�[\����J��RJ\�8�A���v�{���LB!?�	!f('^��: ���ؕ��xա>�m3:�I	�~��%����!Q)�.�˚� �{��"�]Xs�3��R��_M�AmF�c����@]t����<�����P�T���!=�i��~� XP��%�'�S%.^aL�+�����FQ����z�Z����Z
S��9HB��G.9琮F\';���@>�{�H�&ۏ>r�F�;�l�w�7W��@���Г�t՚�!������J�I���Y&��F��܂��%��s���h3�N6{�!�Ap��J�H>�\짉&G��$�3*="���aР�������y
%�1���X	���s���wU�낙��P��>�ǆӝ߀�E8ծᅱ@R�v���%o�uՑ ��"��9^��jї [gP�6�n��J����`�VD���XOH}y�b�:
��^�m��u��{�M:�ﭠ�}
�Ё�c[}kx<|�-53gl����B	�Z��@T�%UO���LgNc�2�>˾WA��#�
%HN�{����e��?�e��~�m� ��$g����6���϶y����������|�����v_�}; 5�����>�u�!+�Jg�*E��:A�@��{[�Y�|�Pg3����r& ��������
	j�A6�M}�*�g��w|��:,IA��P����'��:s��3<*�y�)��:�����i��.���Փ����)�S��óD�D��V4c�(�ks�f}�@�[~m,�`�?gk!3G�_��]��`�&�`2���Q�L�.��@6	Ҁa"sq ��	 >�%��WzQ��	ޟ60N�PM����Ɲ�\J���<�B$QҒ7l�+t�̧~�i)}�࣫���D�\J#כ8���X��K�l'��e�N=/Vt��8�f�E�V�+��AT#w��w�w�����vUmܰ�}�H��S�]5��`�1W%�V���d�TX��.fF93J.)7��@	^Lz-�X�u�e	�W����x0}"SDM0{������K��ʰ�Rst��O���Lz���O��lF�uN����"�rYhh�$��:�u�ҧ<{���
U�%֑��$�M߸�z�%V��^��*>��Rq����>���6���E�f(O�������\ s�c���A0��=�%���m�צl�� d�#��b��W""����5p�ͧ��P\�q]��N�C.�X$�P!e$�5���G�P��;���D����%,?#�[�ULMVJ�q�v�,��M��"�:l=�vl���'��&Kr�����
��ܔ@�Y!�g}�h�$.g��U^����C
�{`��C�Եo-?ܹ���P���&"���+��:G�������l7����?2��3�J�6�
�C4�cgr������Ke����m�Yr��	W��;��a�1��,7�I�|&�ء�-m�6���l�7�fDqh�<��v���0��O�q#�L���3Z9gv]����߱*�=�\>yr�����2u�!9 ���������lx[���߯�P�J�������ɏ	��;d)
��ˁ�a�kp+6:S���O���A��M�g���}��"����]7�B	���/E^�U\�טI?	�̻sy�(t��>ߟVP�7>W"�zC'�5V�[�\�#�)d���gd� �3����%������Ǻ�_[8�nb�Ȝ����ɣ��