// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 15:05:47 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Kud1RDYTDXUneivDgMBZWZ00o3Z3eAAgObvNmI73kF+q7aylPx7Vmrdbkav6rpcC
Lg1+ngX+4eyNCwfq3yYVMv8pAOIXYwApkvRVbypyV9pg8RYPzqLrUUnJyWyLNUwl
teEp3LS7fWpGShocv5n+/YrZKmW2LO3KgH550UtHVt8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2064)
Ok9kvX81FD4XPrQPLgvQ0uv7q06OZlvu0awbSLfys9wNyewx38Z5cJFCxHwoXM2t
F8NI+a4G9GyXegQEDNMMjL3+qiJfX5iMrCWVKvFrn4sEBLEshih+n/NfcJiUgjEm
q+N4kCbVljUxYVdbt6sKPHjL4cVk/OGinCw+ScexkxpnvTBOtaOth9s/BuwRbtSH
Wm6VkM/zDhNBHqo1dVUbc/bV/I2A0SI54cm9Sy4lxTGapGvkPBuhUjPRYZQDzmE3
gxrUNGWpejU/apvziOa5/iOPZTzM9VIa5j756NZBQ/O4clca9C9+iX6EaaMr+H/G
2hGrLhLaMFMVXdL5urSg4CfNxVn+dkwATH6xy/5OUbz4mCY5NMujuj8kIJfwF0Xs
+OC/iv4YglKiNQo8iWQD+sB5S8nCQSvVbqffUnhVMYVJGto1KCkcAHurH50VRWAp
i4uTcyUM6cPhiK+SM06l53b5mWEuC84C/ZSwG8pP5nDCGpQD04qVCZiUVp/1mjTE
4qAa/E63sfAPR2NSO35ZEu6zSjv3F/XFGuecUyNPiMCoDGpLL2CbiyEkpFR8c/UI
D1+TIHIYvw9kas6q/xsAqmug+pqyVJCuazvOWm62F8pP5EUTiHGQfLPJEvlHwWAh
IeegxN4g+4uBnTwJgioJRAddcPZN2/MQZeg925c9D/0dGRQI/L9wXSy4bF8/BnhJ
bt2bh4dAPk5mryd4d9GT+CmXangjtdKr9B8YfOHxw6IhFo74Wtg+mZkc5xx6XBrs
cOMab7N6rJDuIuS4RtIY2btnYen0WU26ZVXxj8TkAhFWCxqjP9LumqKAkccBpTdI
UbPWNhpQAHLG7XZkXG8VBWib52xbvgSH/f8GiK2wEO/DUC7pCgIxBYXwb6yz3AH6
7T4/Uk41KT4jL3O1uNYURxCOgMUxaAiYNZiWWC4Vm3a9uysQdoDzL50yOCmZi9KA
f70DP8Q0z/WLmBrNrnvkimxhuzkHbYzLnGW64Z4WPLNSKgjbfi8vIDjRqgHCOd7W
DaYCaBihxQpZfJXtgGPlrEorEA4ef0B4nInq8E8xmw2txA0NpFCcG3xF8nuLpZpZ
Nu05QyIPlbhtijWFydqWvyk2ndWyRmhJ+cxmCrZdkkZG8AA+maWD10LLOM9yNcrz
AEViREnFhz9HuwtP6KcpdGxtyuBe21LJ4hf0q3RCZNMu78t5+lARWkTT7KGFLuGk
APYIi4LKxSW1XxuhOp5yySH2Tj+4Ws6mtuojs5jPZIONdro/KJbV03dpd6tvUx98
DQn/t94U2W68VzCQ0nHg/s4SHqBnzkZA5vZsT9cxFhCAOdLaoVHlMkTpSSQbtLDV
51scn+la937cEWSFARF1KpoKwy52zvpLkG11305CrdP+5if+qAelkgM1ZtjeQmh7
45c+onIDlJYRVfP7V0PDEdXGrEgMrebm0iU7T0MdoTPIidmBe/1lIa/iSxF+Z1u0
TQA8li6u0uPaeGhRyKD+5mfLrDOGGe8Bb6K8kOv+LSReleN3i20LenNi/isuNeXR
97jYh5XRajluiGlXizHk+vqMkCmdnKE8bk5sjBamcp0g10IqHbwP3e5JYb13jeAl
d+q9d0Qggj682H/gWeoc9GAEbXYr5W+KvKZ43FYBYaitkb4Vs14OV7zWcLbeifz8
x52UOw4jN9oLWLPyOuXz8nyrqXWxfjtNSH7KyKHWfYhefW4Z24DdukmMMI6OawGw
MgooAvs5TZkOgUHQ8sE8sgbGZtyB16faEmVfQD7iOxpIk9qV0OoZM1j6mZKs75ze
7o1kFcRh0cMeTOLibVmllf/47lUDuXK9M9wuP0NxSSYc6ZLq4MT39JEnNDX0NugZ
WSVLLSyXV2I/BL0/IiLgPgEXF7/K12E180IHvGU5NZwQGZGTksulc1EW75RZ5mxd
jsODiUuyU2oO6bMTyf9/TX4YvO20BTWIDA3lA87tlRqGhBu277395ox5+DHoQIBX
ztKTewXemu+8/3TOlFeeGgAoikoIwIvtxM3eyI2YlzNKbuvtNcn/YCn91x1tXCrg
X3fmkHF1eURoJtclO9QanurQ37+hwovd3f57kgsoOu6QUmqAfV/97harLslJ4Cn9
+tc9lKe+I1gvdRrkBOGW+dDPSEakORwvhFpRRdy0RanLiuaWF/k+lK9hZdCoT1lT
uKFwHO0W79fZMzdXfr7Mc2q87WJqnlh757RIUyU0492Q9CfTQM+j/3N45tOr8CX3
PZtl8z0AXbMGsIxEhgTTxX21xaVqWf1oevRkq2mj/8vogy8u8EGQ5P3sVvj6Bjhf
uIqyM6rp0fUC673IdE/6Q/pgbZfxkQNKcr+6RmGBj3xZtdGYbN39tWMHKEpMUsYB
su6BEkWWJYTC5tfYjQN+dTpI0ucF/WejvDhA9t4nsXJyygOmWoS7N8cYVpDoPm2o
F4lK03KviclrweRVpBnx0xtmzVy0oepdrI0g8FSc92BE0w1fOa00fVFCK+Wj1ri3
2SDdLHlsmDfCrG5IqjYh9A9TTzYW+zQkPcyVh1AUbvBBOjKJAhVODZ7jpD9vW62q
RnNo9JiTIeuk6jDS/1vc/2DvhGkFes+OfB9jt9blh2bKiUwtbDuRslTSNOAvn7+n
FFe+pGLCBINxgTnzbcWQmid9LSTH+LxXg/3D542tJVU0hoXdXYG9kWL1N32hClWU
2qGErQHo9My4psr2xwYio51Gd8n3+wmdkXrVd4sb5sLFp0ywd/9L3aemr3X4w6UC
`pragma protect end_protected
