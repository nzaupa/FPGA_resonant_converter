��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-}�&N��<a�6H�w�#e�S!=T�c�+~�
e�� b^��>y��Z׀vi����m�?3�QEx�~��/ҝ��E¦���Tc.ǟ�k�5�39��D�v'�(�ɍ���_��{:Ow��fAdi�lu�xY�8g*I�.��x�Ǌ}]Gy�!u�N�.�P�"!ܒc�0��ЍՔkD���Ҍ�ǃz�@L��h���lf�!��6~|+ޕp�=8�U|?ѻ?#�����jX��H�A���Hj��묅%��;ol�$gM��r
��;�vy���Vop"���|����݋E���4�s�ʪ.I��t^9�w�#\���n���T5�{���X��.ὑQM�=Ćb��%�E�5�U����W;�'���7���Q
��ӂ������!�����5���3p��l�6yx��� �;.��M9��V�/��kv���qk��:�U�X�3���שĖ��b	I } ����o�$�op��s�}`;�;m�&}aA����� 9�DX�%����Ru�������F?��WhW,݊�}�8���}��$���c_�m���P�b�3�DH��|[�������{7	�a
��&Ɠ�p�}�.�$y�+0�6il���`�.���;�8)�c�Y1ox���9�����$��]�WA_Q8u^6�T;�#�cEo��n]D9��wm�<.���9���N*<�L��x���]����YD��#9؜u��M�ȁ,�m4���@aY��
�|;�Py����=��5�[?m��R���R��}���O;��c�rK���)*�Ca QJ�N"K�ɻ_�[���3�(h�oX������~�L#��!�A�:��$�{K�!ޘ�V�2l�IЪ�]�t��W�E
��n����7 �Ь�M~�cC�
��ؓ�,�q|惞1�(Q��W�Y|��M ��MK���R_T��@�3j5��^j!�C@E��#B(�ŬΏh���#��+j�O_0w�k�楲0h����:6��^u볭��{��@���`���Rȉ��hTF�A0�v��v�5M2�Œ�5�#v3��.qO�^}��B�����,���m_0� [_�'ޭ������*�]n�o�f�!�/=RT@�js��>v[���%�G��A+�fM]@5-�H���́ݧM̤��Vr���R,�U��<?���ϙ����"���\e��e�UjV����U�e)2
�ۈ��SM$�۲2���q�wl|��k:�Y]y��nZ�����w�����T��U#��w�����F�(����n�x9���Cr8P�ʊ7]�M~sh�M]p#e)/�����Y�9yP︧~J���X�<����Ewg�Z���2�9��K��{T��k�H�Ȗ�0Z(���km�%$��%���f�[T3#�u�i"-ş6n\Ѳ��%�V��)��}�G]�\zȒ!^b��^�(�$U5�0��p���f��;���Я���Gl\�*E$�5����!�Z3S�Wl����}��/}"/�ʽ���Zg%:�
��\�\�a*4��Y�����J�ի��8�ʒ�5S�t�}��S}K��zP��9ήt/I�jJC�E���@��yN����E��Ii�!��A����h"���-�a�Uz,��"v<���EaJ��B�Cr�v�DJ^Q�߷eD>��T��x������ �BNOu��"�U�>t���.��:���gL˸��.�M�[�N�=g$��_��m���_�A�g!�!ɝ�5�E���c2��}_`�ެ���O-��+Q�A1�PyLHаZ&�a����0Ｌ.��$}��	�&�'�d(�w[\��4���~Y�k��[_�A�9'�/<�d�&jbv�3:��+~sb=�\��a@~�3�T�,g�Ĕ.��f@ '�՗FwꙔ��q[��ARb`� e�����i���S%����^
�6��vYƅi8	W,Mƭ*d� u���(|m�0́�5���n�%���S |�06w� 8���63Tܤ)�݈ڽ�p�:�Y���E����gZji�@b[� ��K��