//------------------------------------------------------------
// Project: HYBRID_CONTROL
// Author: Nicola Zaupa
// Date: (2022/02/14) (10:37:59)
// File: trigonometry.v
//------------------------------------------------------------
// Description:
//
// Compuation of sine and cosine of an angle [-pi,2*pi]
// angle  x 100
// output x 1000
//------------------------------------------------------------


`timescale 1 ns / 1 ps
//`default_nettype none


module trigonometry (
   o_cos,    // cosine of the input
   o_sin,    // sine of the input
   i_theta   // input angle
);

output [31:0] o_sin;
output [31:0] o_cos;
input  [31:0] i_theta;

// output  signed [31:0] o_sin;
// output  signed [31:0] o_cos;
// input   signed [31:0] i_theta;

// wire [31:0] o_sin;
// wire [31:0] o_cos;
// wire [31:0] i_theta;

reg [31:0] r_sin;
reg [31:0] r_cos;

assign o_sin = r_sin;
assign o_cos = r_cos;


always @ ( i_theta )
begin

// computation of sine and cosine using integers
// taking advanatges of look-up-table
// input angle is multiplied by x100
// trigonometric output is multiplied by x1000

case(i_theta)
      32'hFFFFFEC6: r_sin = 32'hFFFFFFFE;
      32'hFFFFFEC7: r_sin = 32'hFFFFFFF4;
      32'hFFFFFEC8: r_sin = 32'hFFFFFFEA;
      32'hFFFFFEC9: r_sin = 32'hFFFFFFE0;
      32'hFFFFFECA: r_sin = 32'hFFFFFFD6;
      32'hFFFFFECB: r_sin = 32'hFFFFFFCC;
      32'hFFFFFECC: r_sin = 32'hFFFFFFC2;
      32'hFFFFFECD: r_sin = 32'hFFFFFFB8;
      32'hFFFFFECE: r_sin = 32'hFFFFFFAE;
      32'hFFFFFECF: r_sin = 32'hFFFFFFA5;
      32'hFFFFFED0: r_sin = 32'hFFFFFF9B;
      32'hFFFFFED1: r_sin = 32'hFFFFFF91;
      32'hFFFFFED2: r_sin = 32'hFFFFFF87;
      32'hFFFFFED3: r_sin = 32'hFFFFFF7D;
      32'hFFFFFED4: r_sin = 32'hFFFFFF73;
      32'hFFFFFED5: r_sin = 32'hFFFFFF69;
      32'hFFFFFED6: r_sin = 32'hFFFFFF5F;
      32'hFFFFFED7: r_sin = 32'hFFFFFF55;
      32'hFFFFFED8: r_sin = 32'hFFFFFF4B;
      32'hFFFFFED9: r_sin = 32'hFFFFFF42;
      32'hFFFFFEDA: r_sin = 32'hFFFFFF38;
      32'hFFFFFEDB: r_sin = 32'hFFFFFF2E;
      32'hFFFFFEDC: r_sin = 32'hFFFFFF24;
      32'hFFFFFEDD: r_sin = 32'hFFFFFF1A;
      32'hFFFFFEDE: r_sin = 32'hFFFFFF11;
      32'hFFFFFEDF: r_sin = 32'hFFFFFF07;
      32'hFFFFFEE0: r_sin = 32'hFFFFFEFD;
      32'hFFFFFEE1: r_sin = 32'hFFFFFEF4;
      32'hFFFFFEE2: r_sin = 32'hFFFFFEEA;
      32'hFFFFFEE3: r_sin = 32'hFFFFFEE1;
      32'hFFFFFEE4: r_sin = 32'hFFFFFED7;
      32'hFFFFFEE5: r_sin = 32'hFFFFFECD;
      32'hFFFFFEE6: r_sin = 32'hFFFFFEC4;
      32'hFFFFFEE7: r_sin = 32'hFFFFFEBA;
      32'hFFFFFEE8: r_sin = 32'hFFFFFEB1;
      32'hFFFFFEE9: r_sin = 32'hFFFFFEA8;
      32'hFFFFFEEA: r_sin = 32'hFFFFFE9E;
      32'hFFFFFEEB: r_sin = 32'hFFFFFE95;
      32'hFFFFFEEC: r_sin = 32'hFFFFFE8C;
      32'hFFFFFEED: r_sin = 32'hFFFFFE82;
      32'hFFFFFEEE: r_sin = 32'hFFFFFE79;
      32'hFFFFFEEF: r_sin = 32'hFFFFFE70;
      32'hFFFFFEF0: r_sin = 32'hFFFFFE67;
      32'hFFFFFEF1: r_sin = 32'hFFFFFE5E;
      32'hFFFFFEF2: r_sin = 32'hFFFFFE55;
      32'hFFFFFEF3: r_sin = 32'hFFFFFE4C;
      32'hFFFFFEF4: r_sin = 32'hFFFFFE43;
      32'hFFFFFEF5: r_sin = 32'hFFFFFE3A;
      32'hFFFFFEF6: r_sin = 32'hFFFFFE31;
      32'hFFFFFEF7: r_sin = 32'hFFFFFE28;
      32'hFFFFFEF8: r_sin = 32'hFFFFFE1F;
      32'hFFFFFEF9: r_sin = 32'hFFFFFE16;
      32'hFFFFFEFA: r_sin = 32'hFFFFFE0E;
      32'hFFFFFEFB: r_sin = 32'hFFFFFE05;
      32'hFFFFFEFC: r_sin = 32'hFFFFFDFC;
      32'hFFFFFEFD: r_sin = 32'hFFFFFDF4;
      32'hFFFFFEFE: r_sin = 32'hFFFFFDEB;
      32'hFFFFFEFF: r_sin = 32'hFFFFFDE3;
      32'hFFFFFF00: r_sin = 32'hFFFFFDDB;
      32'hFFFFFF01: r_sin = 32'hFFFFFDD2;
      32'hFFFFFF02: r_sin = 32'hFFFFFDCA;
      32'hFFFFFF03: r_sin = 32'hFFFFFDC2;
      32'hFFFFFF04: r_sin = 32'hFFFFFDBA;
      32'hFFFFFF05: r_sin = 32'hFFFFFDB2;
      32'hFFFFFF06: r_sin = 32'hFFFFFDAA;
      32'hFFFFFF07: r_sin = 32'hFFFFFDA2;
      32'hFFFFFF08: r_sin = 32'hFFFFFD9A;
      32'hFFFFFF09: r_sin = 32'hFFFFFD92;
      32'hFFFFFF0A: r_sin = 32'hFFFFFD8A;
      32'hFFFFFF0B: r_sin = 32'hFFFFFD82;
      32'hFFFFFF0C: r_sin = 32'hFFFFFD7B;
      32'hFFFFFF0D: r_sin = 32'hFFFFFD73;
      32'hFFFFFF0E: r_sin = 32'hFFFFFD6B;
      32'hFFFFFF0F: r_sin = 32'hFFFFFD64;
      32'hFFFFFF10: r_sin = 32'hFFFFFD5D;
      32'hFFFFFF11: r_sin = 32'hFFFFFD55;
      32'hFFFFFF12: r_sin = 32'hFFFFFD4E;
      32'hFFFFFF13: r_sin = 32'hFFFFFD47;
      32'hFFFFFF14: r_sin = 32'hFFFFFD40;
      32'hFFFFFF15: r_sin = 32'hFFFFFD39;
      32'hFFFFFF16: r_sin = 32'hFFFFFD32;
      32'hFFFFFF17: r_sin = 32'hFFFFFD2B;
      32'hFFFFFF18: r_sin = 32'hFFFFFD24;
      32'hFFFFFF19: r_sin = 32'hFFFFFD1D;
      32'hFFFFFF1A: r_sin = 32'hFFFFFD16;
      32'hFFFFFF1B: r_sin = 32'hFFFFFD10;
      32'hFFFFFF1C: r_sin = 32'hFFFFFD09;
      32'hFFFFFF1D: r_sin = 32'hFFFFFD03;
      32'hFFFFFF1E: r_sin = 32'hFFFFFCFC;
      32'hFFFFFF1F: r_sin = 32'hFFFFFCF6;
      32'hFFFFFF20: r_sin = 32'hFFFFFCF0;
      32'hFFFFFF21: r_sin = 32'hFFFFFCEA;
      32'hFFFFFF22: r_sin = 32'hFFFFFCE3;
      32'hFFFFFF23: r_sin = 32'hFFFFFCDD;
      32'hFFFFFF24: r_sin = 32'hFFFFFCD8;
      32'hFFFFFF25: r_sin = 32'hFFFFFCD2;
      32'hFFFFFF26: r_sin = 32'hFFFFFCCC;
      32'hFFFFFF27: r_sin = 32'hFFFFFCC6;
      32'hFFFFFF28: r_sin = 32'hFFFFFCC1;
      32'hFFFFFF29: r_sin = 32'hFFFFFCBB;
      32'hFFFFFF2A: r_sin = 32'hFFFFFCB6;
      32'hFFFFFF2B: r_sin = 32'hFFFFFCB0;
      32'hFFFFFF2C: r_sin = 32'hFFFFFCAB;
      32'hFFFFFF2D: r_sin = 32'hFFFFFCA6;
      32'hFFFFFF2E: r_sin = 32'hFFFFFCA1;
      32'hFFFFFF2F: r_sin = 32'hFFFFFC9C;
      32'hFFFFFF30: r_sin = 32'hFFFFFC97;
      32'hFFFFFF31: r_sin = 32'hFFFFFC92;
      32'hFFFFFF32: r_sin = 32'hFFFFFC8D;
      32'hFFFFFF33: r_sin = 32'hFFFFFC89;
      32'hFFFFFF34: r_sin = 32'hFFFFFC84;
      32'hFFFFFF35: r_sin = 32'hFFFFFC80;
      32'hFFFFFF36: r_sin = 32'hFFFFFC7B;
      32'hFFFFFF37: r_sin = 32'hFFFFFC77;
      32'hFFFFFF38: r_sin = 32'hFFFFFC73;
      32'hFFFFFF39: r_sin = 32'hFFFFFC6F;
      32'hFFFFFF3A: r_sin = 32'hFFFFFC6B;
      32'hFFFFFF3B: r_sin = 32'hFFFFFC67;
      32'hFFFFFF3C: r_sin = 32'hFFFFFC63;
      32'hFFFFFF3D: r_sin = 32'hFFFFFC5F;
      32'hFFFFFF3E: r_sin = 32'hFFFFFC5B;
      32'hFFFFFF3F: r_sin = 32'hFFFFFC58;
      32'hFFFFFF40: r_sin = 32'hFFFFFC54;
      32'hFFFFFF41: r_sin = 32'hFFFFFC51;
      32'hFFFFFF42: r_sin = 32'hFFFFFC4E;
      32'hFFFFFF43: r_sin = 32'hFFFFFC4B;
      32'hFFFFFF44: r_sin = 32'hFFFFFC47;
      32'hFFFFFF45: r_sin = 32'hFFFFFC44;
      32'hFFFFFF46: r_sin = 32'hFFFFFC42;
      32'hFFFFFF47: r_sin = 32'hFFFFFC3F;
      32'hFFFFFF48: r_sin = 32'hFFFFFC3C;
      32'hFFFFFF49: r_sin = 32'hFFFFFC39;
      32'hFFFFFF4A: r_sin = 32'hFFFFFC37;
      32'hFFFFFF4B: r_sin = 32'hFFFFFC34;
      32'hFFFFFF4C: r_sin = 32'hFFFFFC32;
      32'hFFFFFF4D: r_sin = 32'hFFFFFC30;
      32'hFFFFFF4E: r_sin = 32'hFFFFFC2E;
      32'hFFFFFF4F: r_sin = 32'hFFFFFC2C;
      32'hFFFFFF50: r_sin = 32'hFFFFFC2A;
      32'hFFFFFF51: r_sin = 32'hFFFFFC28;
      32'hFFFFFF52: r_sin = 32'hFFFFFC26;
      32'hFFFFFF53: r_sin = 32'hFFFFFC25;
      32'hFFFFFF54: r_sin = 32'hFFFFFC23;
      32'hFFFFFF55: r_sin = 32'hFFFFFC22;
      32'hFFFFFF56: r_sin = 32'hFFFFFC20;
      32'hFFFFFF57: r_sin = 32'hFFFFFC1F;
      32'hFFFFFF58: r_sin = 32'hFFFFFC1E;
      32'hFFFFFF59: r_sin = 32'hFFFFFC1D;
      32'hFFFFFF5A: r_sin = 32'hFFFFFC1C;
      32'hFFFFFF5B: r_sin = 32'hFFFFFC1B;
      32'hFFFFFF5C: r_sin = 32'hFFFFFC1A;
      32'hFFFFFF5D: r_sin = 32'hFFFFFC1A;
      32'hFFFFFF5E: r_sin = 32'hFFFFFC19;
      32'hFFFFFF5F: r_sin = 32'hFFFFFC19;
      32'hFFFFFF60: r_sin = 32'hFFFFFC18;
      32'hFFFFFF61: r_sin = 32'hFFFFFC18;
      32'hFFFFFF62: r_sin = 32'hFFFFFC18;
      32'hFFFFFF63: r_sin = 32'hFFFFFC18;
      32'hFFFFFF64: r_sin = 32'hFFFFFC18;
      32'hFFFFFF65: r_sin = 32'hFFFFFC18;
      32'hFFFFFF66: r_sin = 32'hFFFFFC18;
      32'hFFFFFF67: r_sin = 32'hFFFFFC19;
      32'hFFFFFF68: r_sin = 32'hFFFFFC19;
      32'hFFFFFF69: r_sin = 32'hFFFFFC1A;
      32'hFFFFFF6A: r_sin = 32'hFFFFFC1B;
      32'hFFFFFF6B: r_sin = 32'hFFFFFC1B;
      32'hFFFFFF6C: r_sin = 32'hFFFFFC1C;
      32'hFFFFFF6D: r_sin = 32'hFFFFFC1D;
      32'hFFFFFF6E: r_sin = 32'hFFFFFC1E;
      32'hFFFFFF6F: r_sin = 32'hFFFFFC1F;
      32'hFFFFFF70: r_sin = 32'hFFFFFC21;
      32'hFFFFFF71: r_sin = 32'hFFFFFC22;
      32'hFFFFFF72: r_sin = 32'hFFFFFC23;
      32'hFFFFFF73: r_sin = 32'hFFFFFC25;
      32'hFFFFFF74: r_sin = 32'hFFFFFC27;
      32'hFFFFFF75: r_sin = 32'hFFFFFC28;
      32'hFFFFFF76: r_sin = 32'hFFFFFC2A;
      32'hFFFFFF77: r_sin = 32'hFFFFFC2C;
      32'hFFFFFF78: r_sin = 32'hFFFFFC2E;
      32'hFFFFFF79: r_sin = 32'hFFFFFC30;
      32'hFFFFFF7A: r_sin = 32'hFFFFFC33;
      32'hFFFFFF7B: r_sin = 32'hFFFFFC35;
      32'hFFFFFF7C: r_sin = 32'hFFFFFC37;
      32'hFFFFFF7D: r_sin = 32'hFFFFFC3A;
      32'hFFFFFF7E: r_sin = 32'hFFFFFC3C;
      32'hFFFFFF7F: r_sin = 32'hFFFFFC3F;
      32'hFFFFFF80: r_sin = 32'hFFFFFC42;
      32'hFFFFFF81: r_sin = 32'hFFFFFC45;
      32'hFFFFFF82: r_sin = 32'hFFFFFC48;
      32'hFFFFFF83: r_sin = 32'hFFFFFC4B;
      32'hFFFFFF84: r_sin = 32'hFFFFFC4E;
      32'hFFFFFF85: r_sin = 32'hFFFFFC52;
      32'hFFFFFF86: r_sin = 32'hFFFFFC55;
      32'hFFFFFF87: r_sin = 32'hFFFFFC58;
      32'hFFFFFF88: r_sin = 32'hFFFFFC5C;
      32'hFFFFFF89: r_sin = 32'hFFFFFC60;
      32'hFFFFFF8A: r_sin = 32'hFFFFFC63;
      32'hFFFFFF8B: r_sin = 32'hFFFFFC67;
      32'hFFFFFF8C: r_sin = 32'hFFFFFC6B;
      32'hFFFFFF8D: r_sin = 32'hFFFFFC6F;
      32'hFFFFFF8E: r_sin = 32'hFFFFFC73;
      32'hFFFFFF8F: r_sin = 32'hFFFFFC78;
      32'hFFFFFF90: r_sin = 32'hFFFFFC7C;
      32'hFFFFFF91: r_sin = 32'hFFFFFC80;
      32'hFFFFFF92: r_sin = 32'hFFFFFC85;
      32'hFFFFFF93: r_sin = 32'hFFFFFC89;
      32'hFFFFFF94: r_sin = 32'hFFFFFC8E;
      32'hFFFFFF95: r_sin = 32'hFFFFFC93;
      32'hFFFFFF96: r_sin = 32'hFFFFFC98;
      32'hFFFFFF97: r_sin = 32'hFFFFFC9D;
      32'hFFFFFF98: r_sin = 32'hFFFFFCA2;
      32'hFFFFFF99: r_sin = 32'hFFFFFCA7;
      32'hFFFFFF9A: r_sin = 32'hFFFFFCAC;
      32'hFFFFFF9B: r_sin = 32'hFFFFFCB1;
      32'hFFFFFF9C: r_sin = 32'hFFFFFCB7;
      32'hFFFFFF9D: r_sin = 32'hFFFFFCBC;
      32'hFFFFFF9E: r_sin = 32'hFFFFFCC2;
      32'hFFFFFF9F: r_sin = 32'hFFFFFCC7;
      32'hFFFFFFA0: r_sin = 32'hFFFFFCCD;
      32'hFFFFFFA1: r_sin = 32'hFFFFFCD3;
      32'hFFFFFFA2: r_sin = 32'hFFFFFCD8;
      32'hFFFFFFA3: r_sin = 32'hFFFFFCDE;
      32'hFFFFFFA4: r_sin = 32'hFFFFFCE4;
      32'hFFFFFFA5: r_sin = 32'hFFFFFCEA;
      32'hFFFFFFA6: r_sin = 32'hFFFFFCF1;
      32'hFFFFFFA7: r_sin = 32'hFFFFFCF7;
      32'hFFFFFFA8: r_sin = 32'hFFFFFCFD;
      32'hFFFFFFA9: r_sin = 32'hFFFFFD04;
      32'hFFFFFFAA: r_sin = 32'hFFFFFD0A;
      32'hFFFFFFAB: r_sin = 32'hFFFFFD11;
      32'hFFFFFFAC: r_sin = 32'hFFFFFD17;
      32'hFFFFFFAD: r_sin = 32'hFFFFFD1E;
      32'hFFFFFFAE: r_sin = 32'hFFFFFD25;
      32'hFFFFFFAF: r_sin = 32'hFFFFFD2C;
      32'hFFFFFFB0: r_sin = 32'hFFFFFD33;
      32'hFFFFFFB1: r_sin = 32'hFFFFFD3A;
      32'hFFFFFFB2: r_sin = 32'hFFFFFD41;
      32'hFFFFFFB3: r_sin = 32'hFFFFFD48;
      32'hFFFFFFB4: r_sin = 32'hFFFFFD4F;
      32'hFFFFFFB5: r_sin = 32'hFFFFFD56;
      32'hFFFFFFB6: r_sin = 32'hFFFFFD5E;
      32'hFFFFFFB7: r_sin = 32'hFFFFFD65;
      32'hFFFFFFB8: r_sin = 32'hFFFFFD6D;
      32'hFFFFFFB9: r_sin = 32'hFFFFFD74;
      32'hFFFFFFBA: r_sin = 32'hFFFFFD7C;
      32'hFFFFFFBB: r_sin = 32'hFFFFFD83;
      32'hFFFFFFBC: r_sin = 32'hFFFFFD8B;
      32'hFFFFFFBD: r_sin = 32'hFFFFFD93;
      32'hFFFFFFBE: r_sin = 32'hFFFFFD9B;
      32'hFFFFFFBF: r_sin = 32'hFFFFFDA3;
      32'hFFFFFFC0: r_sin = 32'hFFFFFDAB;
      32'hFFFFFFC1: r_sin = 32'hFFFFFDB3;
      32'hFFFFFFC2: r_sin = 32'hFFFFFDBB;
      32'hFFFFFFC3: r_sin = 32'hFFFFFDC3;
      32'hFFFFFFC4: r_sin = 32'hFFFFFDCB;
      32'hFFFFFFC5: r_sin = 32'hFFFFFDD4;
      32'hFFFFFFC6: r_sin = 32'hFFFFFDDC;
      32'hFFFFFFC7: r_sin = 32'hFFFFFDE4;
      32'hFFFFFFC8: r_sin = 32'hFFFFFDED;
      32'hFFFFFFC9: r_sin = 32'hFFFFFDF5;
      32'hFFFFFFCA: r_sin = 32'hFFFFFDFE;
      32'hFFFFFFCB: r_sin = 32'hFFFFFE06;
      32'hFFFFFFCC: r_sin = 32'hFFFFFE0F;
      32'hFFFFFFCD: r_sin = 32'hFFFFFE18;
      32'hFFFFFFCE: r_sin = 32'hFFFFFE21;
      32'hFFFFFFCF: r_sin = 32'hFFFFFE29;
      32'hFFFFFFD0: r_sin = 32'hFFFFFE32;
      32'hFFFFFFD1: r_sin = 32'hFFFFFE3B;
      32'hFFFFFFD2: r_sin = 32'hFFFFFE44;
      32'hFFFFFFD3: r_sin = 32'hFFFFFE4D;
      32'hFFFFFFD4: r_sin = 32'hFFFFFE56;
      32'hFFFFFFD5: r_sin = 32'hFFFFFE5F;
      32'hFFFFFFD6: r_sin = 32'hFFFFFE68;
      32'hFFFFFFD7: r_sin = 32'hFFFFFE71;
      32'hFFFFFFD8: r_sin = 32'hFFFFFE7B;
      32'hFFFFFFD9: r_sin = 32'hFFFFFE84;
      32'hFFFFFFDA: r_sin = 32'hFFFFFE8D;
      32'hFFFFFFDB: r_sin = 32'hFFFFFE96;
      32'hFFFFFFDC: r_sin = 32'hFFFFFEA0;
      32'hFFFFFFDD: r_sin = 32'hFFFFFEA9;
      32'hFFFFFFDE: r_sin = 32'hFFFFFEB3;
      32'hFFFFFFDF: r_sin = 32'hFFFFFEBC;
      32'hFFFFFFE0: r_sin = 32'hFFFFFEC5;
      32'hFFFFFFE1: r_sin = 32'hFFFFFECF;
      32'hFFFFFFE2: r_sin = 32'hFFFFFED8;
      32'hFFFFFFE3: r_sin = 32'hFFFFFEE2;
      32'hFFFFFFE4: r_sin = 32'hFFFFFEEC;
      32'hFFFFFFE5: r_sin = 32'hFFFFFEF5;
      32'hFFFFFFE6: r_sin = 32'hFFFFFEFF;
      32'hFFFFFFE7: r_sin = 32'hFFFFFF09;
      32'hFFFFFFE8: r_sin = 32'hFFFFFF12;
      32'hFFFFFFE9: r_sin = 32'hFFFFFF1C;
      32'hFFFFFFEA: r_sin = 32'hFFFFFF26;
      32'hFFFFFFEB: r_sin = 32'hFFFFFF30;
      32'hFFFFFFEC: r_sin = 32'hFFFFFF39;
      32'hFFFFFFED: r_sin = 32'hFFFFFF43;
      32'hFFFFFFEE: r_sin = 32'hFFFFFF4D;
      32'hFFFFFFEF: r_sin = 32'hFFFFFF57;
      32'hFFFFFFF0: r_sin = 32'hFFFFFF61;
      32'hFFFFFFF1: r_sin = 32'hFFFFFF6B;
      32'hFFFFFFF2: r_sin = 32'hFFFFFF74;
      32'hFFFFFFF3: r_sin = 32'hFFFFFF7E;
      32'hFFFFFFF4: r_sin = 32'hFFFFFF88;
      32'hFFFFFFF5: r_sin = 32'hFFFFFF92;
      32'hFFFFFFF6: r_sin = 32'hFFFFFF9C;
      32'hFFFFFFF7: r_sin = 32'hFFFFFFA6;
      32'hFFFFFFF8: r_sin = 32'hFFFFFFB0;
      32'hFFFFFFF9: r_sin = 32'hFFFFFFBA;
      32'hFFFFFFFA: r_sin = 32'hFFFFFFC4;
      32'hFFFFFFFB: r_sin = 32'hFFFFFFCE;
      32'hFFFFFFFC: r_sin = 32'hFFFFFFD8;
      32'hFFFFFFFD: r_sin = 32'hFFFFFFE2;
      32'hFFFFFFFE: r_sin = 32'hFFFFFFEC;
      32'hFFFFFFFF: r_sin = 32'hFFFFFFF6;
      32'h00000000: r_sin = 32'h00000000;
      32'h00000001: r_sin = 32'h0000000A;
      32'h00000002: r_sin = 32'h00000014;
      32'h00000003: r_sin = 32'h0000001E;
      32'h00000004: r_sin = 32'h00000028;
      32'h00000005: r_sin = 32'h00000032;
      32'h00000006: r_sin = 32'h0000003C;
      32'h00000007: r_sin = 32'h00000046;
      32'h00000008: r_sin = 32'h00000050;
      32'h00000009: r_sin = 32'h0000005A;
      32'h0000000A: r_sin = 32'h00000064;
      32'h0000000B: r_sin = 32'h0000006E;
      32'h0000000C: r_sin = 32'h00000078;
      32'h0000000D: r_sin = 32'h00000082;
      32'h0000000E: r_sin = 32'h0000008C;
      32'h0000000F: r_sin = 32'h00000095;
      32'h00000010: r_sin = 32'h0000009F;
      32'h00000011: r_sin = 32'h000000A9;
      32'h00000012: r_sin = 32'h000000B3;
      32'h00000013: r_sin = 32'h000000BD;
      32'h00000014: r_sin = 32'h000000C7;
      32'h00000015: r_sin = 32'h000000D0;
      32'h00000016: r_sin = 32'h000000DA;
      32'h00000017: r_sin = 32'h000000E4;
      32'h00000018: r_sin = 32'h000000EE;
      32'h00000019: r_sin = 32'h000000F7;
      32'h0000001A: r_sin = 32'h00000101;
      32'h0000001B: r_sin = 32'h0000010B;
      32'h0000001C: r_sin = 32'h00000114;
      32'h0000001D: r_sin = 32'h0000011E;
      32'h0000001E: r_sin = 32'h00000128;
      32'h0000001F: r_sin = 32'h00000131;
      32'h00000020: r_sin = 32'h0000013B;
      32'h00000021: r_sin = 32'h00000144;
      32'h00000022: r_sin = 32'h0000014D;
      32'h00000023: r_sin = 32'h00000157;
      32'h00000024: r_sin = 32'h00000160;
      32'h00000025: r_sin = 32'h0000016A;
      32'h00000026: r_sin = 32'h00000173;
      32'h00000027: r_sin = 32'h0000017C;
      32'h00000028: r_sin = 32'h00000185;
      32'h00000029: r_sin = 32'h0000018F;
      32'h0000002A: r_sin = 32'h00000198;
      32'h0000002B: r_sin = 32'h000001A1;
      32'h0000002C: r_sin = 32'h000001AA;
      32'h0000002D: r_sin = 32'h000001B3;
      32'h0000002E: r_sin = 32'h000001BC;
      32'h0000002F: r_sin = 32'h000001C5;
      32'h00000030: r_sin = 32'h000001CE;
      32'h00000031: r_sin = 32'h000001D7;
      32'h00000032: r_sin = 32'h000001DF;
      32'h00000033: r_sin = 32'h000001E8;
      32'h00000034: r_sin = 32'h000001F1;
      32'h00000035: r_sin = 32'h000001FA;
      32'h00000036: r_sin = 32'h00000202;
      32'h00000037: r_sin = 32'h0000020B;
      32'h00000038: r_sin = 32'h00000213;
      32'h00000039: r_sin = 32'h0000021C;
      32'h0000003A: r_sin = 32'h00000224;
      32'h0000003B: r_sin = 32'h0000022C;
      32'h0000003C: r_sin = 32'h00000235;
      32'h0000003D: r_sin = 32'h0000023D;
      32'h0000003E: r_sin = 32'h00000245;
      32'h0000003F: r_sin = 32'h0000024D;
      32'h00000040: r_sin = 32'h00000255;
      32'h00000041: r_sin = 32'h0000025D;
      32'h00000042: r_sin = 32'h00000265;
      32'h00000043: r_sin = 32'h0000026D;
      32'h00000044: r_sin = 32'h00000275;
      32'h00000045: r_sin = 32'h0000027D;
      32'h00000046: r_sin = 32'h00000284;
      32'h00000047: r_sin = 32'h0000028C;
      32'h00000048: r_sin = 32'h00000293;
      32'h00000049: r_sin = 32'h0000029B;
      32'h0000004A: r_sin = 32'h000002A2;
      32'h0000004B: r_sin = 32'h000002AA;
      32'h0000004C: r_sin = 32'h000002B1;
      32'h0000004D: r_sin = 32'h000002B8;
      32'h0000004E: r_sin = 32'h000002BF;
      32'h0000004F: r_sin = 32'h000002C6;
      32'h00000050: r_sin = 32'h000002CD;
      32'h00000051: r_sin = 32'h000002D4;
      32'h00000052: r_sin = 32'h000002DB;
      32'h00000053: r_sin = 32'h000002E2;
      32'h00000054: r_sin = 32'h000002E9;
      32'h00000055: r_sin = 32'h000002EF;
      32'h00000056: r_sin = 32'h000002F6;
      32'h00000057: r_sin = 32'h000002FC;
      32'h00000058: r_sin = 32'h00000303;
      32'h00000059: r_sin = 32'h00000309;
      32'h0000005A: r_sin = 32'h0000030F;
      32'h0000005B: r_sin = 32'h00000316;
      32'h0000005C: r_sin = 32'h0000031C;
      32'h0000005D: r_sin = 32'h00000322;
      32'h0000005E: r_sin = 32'h00000328;
      32'h0000005F: r_sin = 32'h0000032D;
      32'h00000060: r_sin = 32'h00000333;
      32'h00000061: r_sin = 32'h00000339;
      32'h00000062: r_sin = 32'h0000033E;
      32'h00000063: r_sin = 32'h00000344;
      32'h00000064: r_sin = 32'h00000349;
      32'h00000065: r_sin = 32'h0000034F;
      32'h00000066: r_sin = 32'h00000354;
      32'h00000067: r_sin = 32'h00000359;
      32'h00000068: r_sin = 32'h0000035E;
      32'h00000069: r_sin = 32'h00000363;
      32'h0000006A: r_sin = 32'h00000368;
      32'h0000006B: r_sin = 32'h0000036D;
      32'h0000006C: r_sin = 32'h00000372;
      32'h0000006D: r_sin = 32'h00000377;
      32'h0000006E: r_sin = 32'h0000037B;
      32'h0000006F: r_sin = 32'h00000380;
      32'h00000070: r_sin = 32'h00000384;
      32'h00000071: r_sin = 32'h00000388;
      32'h00000072: r_sin = 32'h0000038D;
      32'h00000073: r_sin = 32'h00000391;
      32'h00000074: r_sin = 32'h00000395;
      32'h00000075: r_sin = 32'h00000399;
      32'h00000076: r_sin = 32'h0000039D;
      32'h00000077: r_sin = 32'h000003A0;
      32'h00000078: r_sin = 32'h000003A4;
      32'h00000079: r_sin = 32'h000003A8;
      32'h0000007A: r_sin = 32'h000003AB;
      32'h0000007B: r_sin = 32'h000003AE;
      32'h0000007C: r_sin = 32'h000003B2;
      32'h0000007D: r_sin = 32'h000003B5;
      32'h0000007E: r_sin = 32'h000003B8;
      32'h0000007F: r_sin = 32'h000003BB;
      32'h00000080: r_sin = 32'h000003BE;
      32'h00000081: r_sin = 32'h000003C1;
      32'h00000082: r_sin = 32'h000003C4;
      32'h00000083: r_sin = 32'h000003C6;
      32'h00000084: r_sin = 32'h000003C9;
      32'h00000085: r_sin = 32'h000003CB;
      32'h00000086: r_sin = 32'h000003CD;
      32'h00000087: r_sin = 32'h000003D0;
      32'h00000088: r_sin = 32'h000003D2;
      32'h00000089: r_sin = 32'h000003D4;
      32'h0000008A: r_sin = 32'h000003D6;
      32'h0000008B: r_sin = 32'h000003D8;
      32'h0000008C: r_sin = 32'h000003D9;
      32'h0000008D: r_sin = 32'h000003DB;
      32'h0000008E: r_sin = 32'h000003DD;
      32'h0000008F: r_sin = 32'h000003DE;
      32'h00000090: r_sin = 32'h000003DF;
      32'h00000091: r_sin = 32'h000003E1;
      32'h00000092: r_sin = 32'h000003E2;
      32'h00000093: r_sin = 32'h000003E3;
      32'h00000094: r_sin = 32'h000003E4;
      32'h00000095: r_sin = 32'h000003E5;
      32'h00000096: r_sin = 32'h000003E5;
      32'h00000097: r_sin = 32'h000003E6;
      32'h00000098: r_sin = 32'h000003E7;
      32'h00000099: r_sin = 32'h000003E7;
      32'h0000009A: r_sin = 32'h000003E8;
      32'h0000009B: r_sin = 32'h000003E8;
      32'h0000009C: r_sin = 32'h000003E8;
      32'h0000009D: r_sin = 32'h000003E8;
      32'h0000009E: r_sin = 32'h000003E8;
      32'h0000009F: r_sin = 32'h000003E8;
      32'h000000A0: r_sin = 32'h000003E8;
      32'h000000A1: r_sin = 32'h000003E7;
      32'h000000A2: r_sin = 32'h000003E7;
      32'h000000A3: r_sin = 32'h000003E6;
      32'h000000A4: r_sin = 32'h000003E6;
      32'h000000A5: r_sin = 32'h000003E5;
      32'h000000A6: r_sin = 32'h000003E4;
      32'h000000A7: r_sin = 32'h000003E3;
      32'h000000A8: r_sin = 32'h000003E2;
      32'h000000A9: r_sin = 32'h000003E1;
      32'h000000AA: r_sin = 32'h000003E0;
      32'h000000AB: r_sin = 32'h000003DE;
      32'h000000AC: r_sin = 32'h000003DD;
      32'h000000AD: r_sin = 32'h000003DB;
      32'h000000AE: r_sin = 32'h000003DA;
      32'h000000AF: r_sin = 32'h000003D8;
      32'h000000B0: r_sin = 32'h000003D6;
      32'h000000B1: r_sin = 32'h000003D4;
      32'h000000B2: r_sin = 32'h000003D2;
      32'h000000B3: r_sin = 32'h000003D0;
      32'h000000B4: r_sin = 32'h000003CE;
      32'h000000B5: r_sin = 32'h000003CC;
      32'h000000B6: r_sin = 32'h000003C9;
      32'h000000B7: r_sin = 32'h000003C7;
      32'h000000B8: r_sin = 32'h000003C4;
      32'h000000B9: r_sin = 32'h000003C1;
      32'h000000BA: r_sin = 32'h000003BE;
      32'h000000BB: r_sin = 32'h000003BC;
      32'h000000BC: r_sin = 32'h000003B9;
      32'h000000BD: r_sin = 32'h000003B5;
      32'h000000BE: r_sin = 32'h000003B2;
      32'h000000BF: r_sin = 32'h000003AF;
      32'h000000C0: r_sin = 32'h000003AC;
      32'h000000C1: r_sin = 32'h000003A8;
      32'h000000C2: r_sin = 32'h000003A5;
      32'h000000C3: r_sin = 32'h000003A1;
      32'h000000C4: r_sin = 32'h0000039D;
      32'h000000C5: r_sin = 32'h00000399;
      32'h000000C6: r_sin = 32'h00000395;
      32'h000000C7: r_sin = 32'h00000391;
      32'h000000C8: r_sin = 32'h0000038D;
      32'h000000C9: r_sin = 32'h00000389;
      32'h000000CA: r_sin = 32'h00000385;
      32'h000000CB: r_sin = 32'h00000380;
      32'h000000CC: r_sin = 32'h0000037C;
      32'h000000CD: r_sin = 32'h00000377;
      32'h000000CE: r_sin = 32'h00000373;
      32'h000000CF: r_sin = 32'h0000036E;
      32'h000000D0: r_sin = 32'h00000369;
      32'h000000D1: r_sin = 32'h00000364;
      32'h000000D2: r_sin = 32'h0000035F;
      32'h000000D3: r_sin = 32'h0000035A;
      32'h000000D4: r_sin = 32'h00000355;
      32'h000000D5: r_sin = 32'h00000350;
      32'h000000D6: r_sin = 32'h0000034A;
      32'h000000D7: r_sin = 32'h00000345;
      32'h000000D8: r_sin = 32'h0000033F;
      32'h000000D9: r_sin = 32'h0000033A;
      32'h000000DA: r_sin = 32'h00000334;
      32'h000000DB: r_sin = 32'h0000032E;
      32'h000000DC: r_sin = 32'h00000328;
      32'h000000DD: r_sin = 32'h00000323;
      32'h000000DE: r_sin = 32'h0000031D;
      32'h000000DF: r_sin = 32'h00000316;
      32'h000000E0: r_sin = 32'h00000310;
      32'h000000E1: r_sin = 32'h0000030A;
      32'h000000E2: r_sin = 32'h00000304;
      32'h000000E3: r_sin = 32'h000002FD;
      32'h000000E4: r_sin = 32'h000002F7;
      32'h000000E5: r_sin = 32'h000002F0;
      32'h000000E6: r_sin = 32'h000002EA;
      32'h000000E7: r_sin = 32'h000002E3;
      32'h000000E8: r_sin = 32'h000002DC;
      32'h000000E9: r_sin = 32'h000002D5;
      32'h000000EA: r_sin = 32'h000002CE;
      32'h000000EB: r_sin = 32'h000002C7;
      32'h000000EC: r_sin = 32'h000002C0;
      32'h000000ED: r_sin = 32'h000002B9;
      32'h000000EE: r_sin = 32'h000002B2;
      32'h000000EF: r_sin = 32'h000002AB;
      32'h000000F0: r_sin = 32'h000002A3;
      32'h000000F1: r_sin = 32'h0000029C;
      32'h000000F2: r_sin = 32'h00000295;
      32'h000000F3: r_sin = 32'h0000028D;
      32'h000000F4: r_sin = 32'h00000285;
      32'h000000F5: r_sin = 32'h0000027E;
      32'h000000F6: r_sin = 32'h00000276;
      32'h000000F7: r_sin = 32'h0000026E;
      32'h000000F8: r_sin = 32'h00000266;
      32'h000000F9: r_sin = 32'h0000025E;
      32'h000000FA: r_sin = 32'h00000256;
      32'h000000FB: r_sin = 32'h0000024E;
      32'h000000FC: r_sin = 32'h00000246;
      32'h000000FD: r_sin = 32'h0000023E;
      32'h000000FE: r_sin = 32'h00000236;
      32'h000000FF: r_sin = 32'h0000022E;
      32'h00000100: r_sin = 32'h00000225;
      32'h00000101: r_sin = 32'h0000021D;
      32'h00000102: r_sin = 32'h00000215;
      32'h00000103: r_sin = 32'h0000020C;
      32'h00000104: r_sin = 32'h00000204;
      32'h00000105: r_sin = 32'h000001FB;
      32'h00000106: r_sin = 32'h000001F2;
      32'h00000107: r_sin = 32'h000001EA;
      32'h00000108: r_sin = 32'h000001E1;
      32'h00000109: r_sin = 32'h000001D8;
      32'h0000010A: r_sin = 32'h000001CF;
      32'h0000010B: r_sin = 32'h000001C6;
      32'h0000010C: r_sin = 32'h000001BD;
      32'h0000010D: r_sin = 32'h000001B4;
      32'h0000010E: r_sin = 32'h000001AB;
      32'h0000010F: r_sin = 32'h000001A2;
      32'h00000110: r_sin = 32'h00000199;
      32'h00000111: r_sin = 32'h00000190;
      32'h00000112: r_sin = 32'h00000187;
      32'h00000113: r_sin = 32'h0000017E;
      32'h00000114: r_sin = 32'h00000174;
      32'h00000115: r_sin = 32'h0000016B;
      32'h00000116: r_sin = 32'h00000162;
      32'h00000117: r_sin = 32'h00000158;
      32'h00000118: r_sin = 32'h0000014F;
      32'h00000119: r_sin = 32'h00000146;
      32'h0000011A: r_sin = 32'h0000013C;
      32'h0000011B: r_sin = 32'h00000133;
      32'h0000011C: r_sin = 32'h00000129;
      32'h0000011D: r_sin = 32'h0000011F;
      32'h0000011E: r_sin = 32'h00000116;
      32'h0000011F: r_sin = 32'h0000010C;
      32'h00000120: r_sin = 32'h00000103;
      32'h00000121: r_sin = 32'h000000F9;
      32'h00000122: r_sin = 32'h000000EF;
      32'h00000123: r_sin = 32'h000000E6;
      32'h00000124: r_sin = 32'h000000DC;
      32'h00000125: r_sin = 32'h000000D2;
      32'h00000126: r_sin = 32'h000000C8;
      32'h00000127: r_sin = 32'h000000BE;
      32'h00000128: r_sin = 32'h000000B5;
      32'h00000129: r_sin = 32'h000000AB;
      32'h0000012A: r_sin = 32'h000000A1;
      32'h0000012B: r_sin = 32'h00000097;
      32'h0000012C: r_sin = 32'h0000008D;
      32'h0000012D: r_sin = 32'h00000083;
      32'h0000012E: r_sin = 32'h00000079;
      32'h0000012F: r_sin = 32'h0000006F;
      32'h00000130: r_sin = 32'h00000065;
      32'h00000131: r_sin = 32'h0000005B;
      32'h00000132: r_sin = 32'h00000052;
      32'h00000133: r_sin = 32'h00000048;
      32'h00000134: r_sin = 32'h0000003E;
      32'h00000135: r_sin = 32'h00000034;
      32'h00000136: r_sin = 32'h0000002A;
      32'h00000137: r_sin = 32'h00000020;
      32'h00000138: r_sin = 32'h00000016;
      32'h00000139: r_sin = 32'h0000000C;
      32'h0000013A: r_sin = 32'h00000000;
      32'h0000013B: r_sin = 32'hFFFFFFF8;
      32'h0000013C: r_sin = 32'hFFFFFFEE;
      32'h0000013D: r_sin = 32'hFFFFFFE4;
      32'h0000013E: r_sin = 32'hFFFFFFDA;
      32'h0000013F: r_sin = 32'hFFFFFFD0;
      32'h00000140: r_sin = 32'hFFFFFFC6;
      32'h00000141: r_sin = 32'hFFFFFFBC;
      32'h00000142: r_sin = 32'hFFFFFFB2;
      32'h00000143: r_sin = 32'hFFFFFFA8;
      32'h00000144: r_sin = 32'hFFFFFF9E;
      32'h00000145: r_sin = 32'hFFFFFF94;
      32'h00000146: r_sin = 32'hFFFFFF8A;
      32'h00000147: r_sin = 32'hFFFFFF80;
      32'h00000148: r_sin = 32'hFFFFFF76;
      32'h00000149: r_sin = 32'hFFFFFF6C;
      32'h0000014A: r_sin = 32'hFFFFFF62;
      32'h0000014B: r_sin = 32'hFFFFFF58;
      32'h0000014C: r_sin = 32'hFFFFFF4F;
      32'h0000014D: r_sin = 32'hFFFFFF45;
      32'h0000014E: r_sin = 32'hFFFFFF3B;
      32'h0000014F: r_sin = 32'hFFFFFF31;
      32'h00000150: r_sin = 32'hFFFFFF27;
      32'h00000151: r_sin = 32'hFFFFFF1E;
      32'h00000152: r_sin = 32'hFFFFFF14;
      32'h00000153: r_sin = 32'hFFFFFF0A;
      32'h00000154: r_sin = 32'hFFFFFF00;
      32'h00000155: r_sin = 32'hFFFFFEF7;
      32'h00000156: r_sin = 32'hFFFFFEED;
      32'h00000157: r_sin = 32'hFFFFFEE4;
      32'h00000158: r_sin = 32'hFFFFFEDA;
      32'h00000159: r_sin = 32'hFFFFFED0;
      32'h0000015A: r_sin = 32'hFFFFFEC7;
      32'h0000015B: r_sin = 32'hFFFFFEBD;
      32'h0000015C: r_sin = 32'hFFFFFEB4;
      32'h0000015D: r_sin = 32'hFFFFFEAB;
      32'h0000015E: r_sin = 32'hFFFFFEA1;
      32'h0000015F: r_sin = 32'hFFFFFE98;
      32'h00000160: r_sin = 32'hFFFFFE8F;
      32'h00000161: r_sin = 32'hFFFFFE85;
      32'h00000162: r_sin = 32'hFFFFFE7C;
      32'h00000163: r_sin = 32'hFFFFFE73;
      32'h00000164: r_sin = 32'hFFFFFE6A;
      32'h00000165: r_sin = 32'hFFFFFE61;
      32'h00000166: r_sin = 32'hFFFFFE58;
      32'h00000167: r_sin = 32'hFFFFFE4E;
      32'h00000168: r_sin = 32'hFFFFFE45;
      32'h00000169: r_sin = 32'hFFFFFE3D;
      32'h0000016A: r_sin = 32'hFFFFFE34;
      32'h0000016B: r_sin = 32'hFFFFFE2B;
      32'h0000016C: r_sin = 32'hFFFFFE22;
      32'h0000016D: r_sin = 32'hFFFFFE19;
      32'h0000016E: r_sin = 32'hFFFFFE11;
      32'h0000016F: r_sin = 32'hFFFFFE08;
      32'h00000170: r_sin = 32'hFFFFFDFF;
      32'h00000171: r_sin = 32'hFFFFFDF7;
      32'h00000172: r_sin = 32'hFFFFFDEE;
      32'h00000173: r_sin = 32'hFFFFFDE6;
      32'h00000174: r_sin = 32'hFFFFFDDD;
      32'h00000175: r_sin = 32'hFFFFFDD5;
      32'h00000176: r_sin = 32'hFFFFFDCD;
      32'h00000177: r_sin = 32'hFFFFFDC4;
      32'h00000178: r_sin = 32'hFFFFFDBC;
      32'h00000179: r_sin = 32'hFFFFFDB4;
      32'h0000017A: r_sin = 32'hFFFFFDAC;
      32'h0000017B: r_sin = 32'hFFFFFDA4;
      32'h0000017C: r_sin = 32'hFFFFFD9C;
      32'h0000017D: r_sin = 32'hFFFFFD94;
      32'h0000017E: r_sin = 32'hFFFFFD8C;
      32'h0000017F: r_sin = 32'hFFFFFD85;
      32'h00000180: r_sin = 32'hFFFFFD7D;
      32'h00000181: r_sin = 32'hFFFFFD75;
      32'h00000182: r_sin = 32'hFFFFFD6E;
      32'h00000183: r_sin = 32'hFFFFFD66;
      32'h00000184: r_sin = 32'hFFFFFD5F;
      32'h00000185: r_sin = 32'hFFFFFD58;
      32'h00000186: r_sin = 32'hFFFFFD50;
      32'h00000187: r_sin = 32'hFFFFFD49;
      32'h00000188: r_sin = 32'hFFFFFD42;
      32'h00000189: r_sin = 32'hFFFFFD3B;
      32'h0000018A: r_sin = 32'hFFFFFD34;
      32'h0000018B: r_sin = 32'hFFFFFD2D;
      32'h0000018C: r_sin = 32'hFFFFFD26;
      32'h0000018D: r_sin = 32'hFFFFFD1F;
      32'h0000018E: r_sin = 32'hFFFFFD18;
      32'h0000018F: r_sin = 32'hFFFFFD12;
      32'h00000190: r_sin = 32'hFFFFFD0B;
      32'h00000191: r_sin = 32'hFFFFFD05;
      32'h00000192: r_sin = 32'hFFFFFCFE;
      32'h00000193: r_sin = 32'hFFFFFCF8;
      32'h00000194: r_sin = 32'hFFFFFCF2;
      32'h00000195: r_sin = 32'hFFFFFCEB;
      32'h00000196: r_sin = 32'hFFFFFCE5;
      32'h00000197: r_sin = 32'hFFFFFCDF;
      32'h00000198: r_sin = 32'hFFFFFCD9;
      32'h00000199: r_sin = 32'hFFFFFCD4;
      32'h0000019A: r_sin = 32'hFFFFFCCE;
      32'h0000019B: r_sin = 32'hFFFFFCC8;
      32'h0000019C: r_sin = 32'hFFFFFCC2;
      32'h0000019D: r_sin = 32'hFFFFFCBD;
      32'h0000019E: r_sin = 32'hFFFFFCB7;
      32'h0000019F: r_sin = 32'hFFFFFCB2;
      32'h000001A0: r_sin = 32'hFFFFFCAD;
      32'h000001A1: r_sin = 32'hFFFFFCA8;
      32'h000001A2: r_sin = 32'hFFFFFCA2;
      32'h000001A3: r_sin = 32'hFFFFFC9D;
      32'h000001A4: r_sin = 32'hFFFFFC98;
      32'h000001A5: r_sin = 32'hFFFFFC94;
      32'h000001A6: r_sin = 32'hFFFFFC8F;
      32'h000001A7: r_sin = 32'hFFFFFC8A;
      32'h000001A8: r_sin = 32'hFFFFFC86;
      32'h000001A9: r_sin = 32'hFFFFFC81;
      32'h000001AA: r_sin = 32'hFFFFFC7D;
      32'h000001AB: r_sin = 32'hFFFFFC78;
      32'h000001AC: r_sin = 32'hFFFFFC74;
      32'h000001AD: r_sin = 32'hFFFFFC70;
      32'h000001AE: r_sin = 32'hFFFFFC6C;
      32'h000001AF: r_sin = 32'hFFFFFC68;
      32'h000001B0: r_sin = 32'hFFFFFC64;
      32'h000001B1: r_sin = 32'hFFFFFC60;
      32'h000001B2: r_sin = 32'hFFFFFC5D;
      32'h000001B3: r_sin = 32'hFFFFFC59;
      32'h000001B4: r_sin = 32'hFFFFFC55;
      32'h000001B5: r_sin = 32'hFFFFFC52;
      32'h000001B6: r_sin = 32'hFFFFFC4F;
      32'h000001B7: r_sin = 32'hFFFFFC4C;
      32'h000001B8: r_sin = 32'hFFFFFC48;
      32'h000001B9: r_sin = 32'hFFFFFC45;
      32'h000001BA: r_sin = 32'hFFFFFC42;
      32'h000001BB: r_sin = 32'hFFFFFC40;
      32'h000001BC: r_sin = 32'hFFFFFC3D;
      32'h000001BD: r_sin = 32'hFFFFFC3A;
      32'h000001BE: r_sin = 32'hFFFFFC38;
      32'h000001BF: r_sin = 32'hFFFFFC35;
      32'h000001C0: r_sin = 32'hFFFFFC33;
      32'h000001C1: r_sin = 32'hFFFFFC31;
      32'h000001C2: r_sin = 32'hFFFFFC2E;
      32'h000001C3: r_sin = 32'hFFFFFC2C;
      32'h000001C4: r_sin = 32'hFFFFFC2A;
      32'h000001C5: r_sin = 32'hFFFFFC29;
      32'h000001C6: r_sin = 32'hFFFFFC27;
      32'h000001C7: r_sin = 32'hFFFFFC25;
      32'h000001C8: r_sin = 32'hFFFFFC24;
      32'h000001C9: r_sin = 32'hFFFFFC22;
      32'h000001CA: r_sin = 32'hFFFFFC21;
      32'h000001CB: r_sin = 32'hFFFFFC1F;
      32'h000001CC: r_sin = 32'hFFFFFC1E;
      32'h000001CD: r_sin = 32'hFFFFFC1D;
      32'h000001CE: r_sin = 32'hFFFFFC1C;
      32'h000001CF: r_sin = 32'hFFFFFC1B;
      32'h000001D0: r_sin = 32'hFFFFFC1B;
      32'h000001D1: r_sin = 32'hFFFFFC1A;
      32'h000001D2: r_sin = 32'hFFFFFC19;
      32'h000001D3: r_sin = 32'hFFFFFC19;
      32'h000001D4: r_sin = 32'hFFFFFC19;
      32'h000001D5: r_sin = 32'hFFFFFC18;
      32'h000001D6: r_sin = 32'hFFFFFC18;
      32'h000001D7: r_sin = 32'hFFFFFC18;
      32'h000001D8: r_sin = 32'hFFFFFC18;
      32'h000001D9: r_sin = 32'hFFFFFC18;
      32'h000001DA: r_sin = 32'hFFFFFC18;
      32'h000001DB: r_sin = 32'hFFFFFC19;
      32'h000001DC: r_sin = 32'hFFFFFC19;
      32'h000001DD: r_sin = 32'hFFFFFC1A;
      32'h000001DE: r_sin = 32'hFFFFFC1A;
      32'h000001DF: r_sin = 32'hFFFFFC1B;
      32'h000001E0: r_sin = 32'hFFFFFC1C;
      32'h000001E1: r_sin = 32'hFFFFFC1D;
      32'h000001E2: r_sin = 32'hFFFFFC1E;
      32'h000001E3: r_sin = 32'hFFFFFC1F;
      32'h000001E4: r_sin = 32'hFFFFFC20;
      32'h000001E5: r_sin = 32'hFFFFFC21;
      32'h000001E6: r_sin = 32'hFFFFFC23;
      32'h000001E7: r_sin = 32'hFFFFFC24;
      32'h000001E8: r_sin = 32'hFFFFFC26;
      32'h000001E9: r_sin = 32'hFFFFFC28;
      32'h000001EA: r_sin = 32'hFFFFFC2A;
      32'h000001EB: r_sin = 32'hFFFFFC2B;
      32'h000001EC: r_sin = 32'hFFFFFC2D;
      32'h000001ED: r_sin = 32'hFFFFFC30;
      32'h000001EE: r_sin = 32'hFFFFFC32;
      32'h000001EF: r_sin = 32'hFFFFFC34;
      32'h000001F0: r_sin = 32'hFFFFFC36;
      32'h000001F1: r_sin = 32'hFFFFFC39;
      32'h000001F2: r_sin = 32'hFFFFFC3C;
      32'h000001F3: r_sin = 32'hFFFFFC3E;
      32'h000001F4: r_sin = 32'hFFFFFC41;
      32'h000001F5: r_sin = 32'hFFFFFC44;
      32'h000001F6: r_sin = 32'hFFFFFC47;
      32'h000001F7: r_sin = 32'hFFFFFC4A;
      32'h000001F8: r_sin = 32'hFFFFFC4D;
      32'h000001F9: r_sin = 32'hFFFFFC50;
      32'h000001FA: r_sin = 32'hFFFFFC54;
      32'h000001FB: r_sin = 32'hFFFFFC57;
      32'h000001FC: r_sin = 32'hFFFFFC5B;
      32'h000001FD: r_sin = 32'hFFFFFC5E;
      32'h000001FE: r_sin = 32'hFFFFFC62;
      32'h000001FF: r_sin = 32'hFFFFFC66;
      32'h00000200: r_sin = 32'hFFFFFC6A;
      32'h00000201: r_sin = 32'hFFFFFC6E;
      32'h00000202: r_sin = 32'hFFFFFC72;
      32'h00000203: r_sin = 32'hFFFFFC76;
      32'h00000204: r_sin = 32'hFFFFFC7B;
      32'h00000205: r_sin = 32'hFFFFFC7F;
      32'h00000206: r_sin = 32'hFFFFFC83;
      32'h00000207: r_sin = 32'hFFFFFC88;
      32'h00000208: r_sin = 32'hFFFFFC8D;
      32'h00000209: r_sin = 32'hFFFFFC91;
      32'h0000020A: r_sin = 32'hFFFFFC96;
      32'h0000020B: r_sin = 32'hFFFFFC9B;
      32'h0000020C: r_sin = 32'hFFFFFCA0;
      32'h0000020D: r_sin = 32'hFFFFFCA5;
      32'h0000020E: r_sin = 32'hFFFFFCAA;
      32'h0000020F: r_sin = 32'hFFFFFCAF;
      32'h00000210: r_sin = 32'hFFFFFCB5;
      32'h00000211: r_sin = 32'hFFFFFCBA;
      32'h00000212: r_sin = 32'hFFFFFCC0;
      32'h00000213: r_sin = 32'hFFFFFCC5;
      32'h00000214: r_sin = 32'hFFFFFCCB;
      32'h00000215: r_sin = 32'hFFFFFCD1;
      32'h00000216: r_sin = 32'hFFFFFCD7;
      32'h00000217: r_sin = 32'hFFFFFCDC;
      32'h00000218: r_sin = 32'hFFFFFCE2;
      32'h00000219: r_sin = 32'hFFFFFCE9;
      32'h0000021A: r_sin = 32'hFFFFFCEF;
      32'h0000021B: r_sin = 32'hFFFFFCF5;
      32'h0000021C: r_sin = 32'hFFFFFCFB;
      32'h0000021D: r_sin = 32'hFFFFFD02;
      32'h0000021E: r_sin = 32'hFFFFFD08;
      32'h0000021F: r_sin = 32'hFFFFFD0F;
      32'h00000220: r_sin = 32'hFFFFFD15;
      32'h00000221: r_sin = 32'hFFFFFD1C;
      32'h00000222: r_sin = 32'hFFFFFD23;
      32'h00000223: r_sin = 32'hFFFFFD2A;
      32'h00000224: r_sin = 32'hFFFFFD30;
      32'h00000225: r_sin = 32'hFFFFFD37;
      32'h00000226: r_sin = 32'hFFFFFD3E;
      32'h00000227: r_sin = 32'hFFFFFD46;
      32'h00000228: r_sin = 32'hFFFFFD4D;
      32'h00000229: r_sin = 32'hFFFFFD54;
      32'h0000022A: r_sin = 32'hFFFFFD5B;
      32'h0000022B: r_sin = 32'hFFFFFD63;
      32'h0000022C: r_sin = 32'hFFFFFD6A;
      32'h0000022D: r_sin = 32'hFFFFFD72;
      32'h0000022E: r_sin = 32'hFFFFFD79;
      32'h0000022F: r_sin = 32'hFFFFFD81;
      32'h00000230: r_sin = 32'hFFFFFD89;
      32'h00000231: r_sin = 32'hFFFFFD91;
      32'h00000232: r_sin = 32'hFFFFFD98;
      32'h00000233: r_sin = 32'hFFFFFDA0;
      32'h00000234: r_sin = 32'hFFFFFDA8;
      32'h00000235: r_sin = 32'hFFFFFDB0;
      32'h00000236: r_sin = 32'hFFFFFDB8;
      32'h00000237: r_sin = 32'hFFFFFDC1;
      32'h00000238: r_sin = 32'hFFFFFDC9;
      32'h00000239: r_sin = 32'hFFFFFDD1;
      32'h0000023A: r_sin = 32'hFFFFFDD9;
      32'h0000023B: r_sin = 32'hFFFFFDE2;
      32'h0000023C: r_sin = 32'hFFFFFDEA;
      32'h0000023D: r_sin = 32'hFFFFFDF3;
      32'h0000023E: r_sin = 32'hFFFFFDFB;
      32'h0000023F: r_sin = 32'hFFFFFE04;
      32'h00000240: r_sin = 32'hFFFFFE0C;
      32'h00000241: r_sin = 32'hFFFFFE15;
      32'h00000242: r_sin = 32'hFFFFFE1E;
      32'h00000243: r_sin = 32'hFFFFFE27;
      32'h00000244: r_sin = 32'hFFFFFE2F;
      32'h00000245: r_sin = 32'hFFFFFE38;
      32'h00000246: r_sin = 32'hFFFFFE41;
      32'h00000247: r_sin = 32'hFFFFFE4A;
      32'h00000248: r_sin = 32'hFFFFFE53;
      32'h00000249: r_sin = 32'hFFFFFE5C;
      32'h0000024A: r_sin = 32'hFFFFFE65;
      32'h0000024B: r_sin = 32'hFFFFFE6E;
      32'h0000024C: r_sin = 32'hFFFFFE78;
      32'h0000024D: r_sin = 32'hFFFFFE81;
      32'h0000024E: r_sin = 32'hFFFFFE8A;
      32'h0000024F: r_sin = 32'hFFFFFE93;
      32'h00000250: r_sin = 32'hFFFFFE9D;
      32'h00000251: r_sin = 32'hFFFFFEA6;
      32'h00000252: r_sin = 32'hFFFFFEB0;
      32'h00000253: r_sin = 32'hFFFFFEB9;
      32'h00000254: r_sin = 32'hFFFFFEC2;
      32'h00000255: r_sin = 32'hFFFFFECC;
      32'h00000256: r_sin = 32'hFFFFFED5;
      32'h00000257: r_sin = 32'hFFFFFEDF;
      32'h00000258: r_sin = 32'hFFFFFEE9;
      32'h00000259: r_sin = 32'hFFFFFEF2;
      32'h0000025A: r_sin = 32'hFFFFFEFC;
      32'h0000025B: r_sin = 32'hFFFFFF06;
      32'h0000025C: r_sin = 32'hFFFFFF0F;
      32'h0000025D: r_sin = 32'hFFFFFF19;
      32'h0000025E: r_sin = 32'hFFFFFF23;
      32'h0000025F: r_sin = 32'hFFFFFF2C;
      32'h00000260: r_sin = 32'hFFFFFF36;
      32'h00000261: r_sin = 32'hFFFFFF40;
      32'h00000262: r_sin = 32'hFFFFFF4A;
      32'h00000263: r_sin = 32'hFFFFFF54;
      32'h00000264: r_sin = 32'hFFFFFF5E;
      32'h00000265: r_sin = 32'hFFFFFF67;
      32'h00000266: r_sin = 32'hFFFFFF71;
      32'h00000267: r_sin = 32'hFFFFFF7B;
      32'h00000268: r_sin = 32'hFFFFFF85;
      32'h00000269: r_sin = 32'hFFFFFF8F;
      32'h0000026A: r_sin = 32'hFFFFFF99;
      32'h0000026B: r_sin = 32'hFFFFFFA3;
      32'h0000026C: r_sin = 32'hFFFFFFAD;
      32'h0000026D: r_sin = 32'hFFFFFFB7;
      32'h0000026E: r_sin = 32'hFFFFFFC1;
      32'h0000026F: r_sin = 32'hFFFFFFCB;
      32'h00000270: r_sin = 32'hFFFFFFD5;
      32'h00000271: r_sin = 32'hFFFFFFDF;
      32'h00000272: r_sin = 32'hFFFFFFE9;
      32'h00000273: r_sin = 32'hFFFFFFF3;
      32'h00000274: r_sin = 32'hFFFFFFFD;
      default: r_sin = 32'h00000000;
endcase

case(i_theta)
      32'hFFFFFEC6: r_cos = 32'hFFFFFC18;
      32'hFFFFFEC7: r_cos = 32'hFFFFFC18;
      32'hFFFFFEC8: r_cos = 32'hFFFFFC18;
      32'hFFFFFEC9: r_cos = 32'hFFFFFC18;
      32'hFFFFFECA: r_cos = 32'hFFFFFC19;
      32'hFFFFFECB: r_cos = 32'hFFFFFC19;
      32'hFFFFFECC: r_cos = 32'hFFFFFC1A;
      32'hFFFFFECD: r_cos = 32'hFFFFFC1B;
      32'hFFFFFECE: r_cos = 32'hFFFFFC1B;
      32'hFFFFFECF: r_cos = 32'hFFFFFC1C;
      32'hFFFFFED0: r_cos = 32'hFFFFFC1D;
      32'hFFFFFED1: r_cos = 32'hFFFFFC1E;
      32'hFFFFFED2: r_cos = 32'hFFFFFC1F;
      32'hFFFFFED3: r_cos = 32'hFFFFFC21;
      32'hFFFFFED4: r_cos = 32'hFFFFFC22;
      32'hFFFFFED5: r_cos = 32'hFFFFFC23;
      32'hFFFFFED6: r_cos = 32'hFFFFFC25;
      32'hFFFFFED7: r_cos = 32'hFFFFFC27;
      32'hFFFFFED8: r_cos = 32'hFFFFFC28;
      32'hFFFFFED9: r_cos = 32'hFFFFFC2A;
      32'hFFFFFEDA: r_cos = 32'hFFFFFC2C;
      32'hFFFFFEDB: r_cos = 32'hFFFFFC2E;
      32'hFFFFFEDC: r_cos = 32'hFFFFFC30;
      32'hFFFFFEDD: r_cos = 32'hFFFFFC33;
      32'hFFFFFEDE: r_cos = 32'hFFFFFC35;
      32'hFFFFFEDF: r_cos = 32'hFFFFFC37;
      32'hFFFFFEE0: r_cos = 32'hFFFFFC3A;
      32'hFFFFFEE1: r_cos = 32'hFFFFFC3D;
      32'hFFFFFEE2: r_cos = 32'hFFFFFC3F;
      32'hFFFFFEE3: r_cos = 32'hFFFFFC42;
      32'hFFFFFEE4: r_cos = 32'hFFFFFC45;
      32'hFFFFFEE5: r_cos = 32'hFFFFFC48;
      32'hFFFFFEE6: r_cos = 32'hFFFFFC4B;
      32'hFFFFFEE7: r_cos = 32'hFFFFFC4E;
      32'hFFFFFEE8: r_cos = 32'hFFFFFC52;
      32'hFFFFFEE9: r_cos = 32'hFFFFFC55;
      32'hFFFFFEEA: r_cos = 32'hFFFFFC59;
      32'hFFFFFEEB: r_cos = 32'hFFFFFC5C;
      32'hFFFFFEEC: r_cos = 32'hFFFFFC60;
      32'hFFFFFEED: r_cos = 32'hFFFFFC64;
      32'hFFFFFEEE: r_cos = 32'hFFFFFC68;
      32'hFFFFFEEF: r_cos = 32'hFFFFFC6C;
      32'hFFFFFEF0: r_cos = 32'hFFFFFC70;
      32'hFFFFFEF1: r_cos = 32'hFFFFFC74;
      32'hFFFFFEF2: r_cos = 32'hFFFFFC78;
      32'hFFFFFEF3: r_cos = 32'hFFFFFC7C;
      32'hFFFFFEF4: r_cos = 32'hFFFFFC81;
      32'hFFFFFEF5: r_cos = 32'hFFFFFC85;
      32'hFFFFFEF6: r_cos = 32'hFFFFFC8A;
      32'hFFFFFEF7: r_cos = 32'hFFFFFC8E;
      32'hFFFFFEF8: r_cos = 32'hFFFFFC93;
      32'hFFFFFEF9: r_cos = 32'hFFFFFC98;
      32'hFFFFFEFA: r_cos = 32'hFFFFFC9D;
      32'hFFFFFEFB: r_cos = 32'hFFFFFCA2;
      32'hFFFFFEFC: r_cos = 32'hFFFFFCA7;
      32'hFFFFFEFD: r_cos = 32'hFFFFFCAC;
      32'hFFFFFEFE: r_cos = 32'hFFFFFCB2;
      32'hFFFFFEFF: r_cos = 32'hFFFFFCB7;
      32'hFFFFFF00: r_cos = 32'hFFFFFCBC;
      32'hFFFFFF01: r_cos = 32'hFFFFFCC2;
      32'hFFFFFF02: r_cos = 32'hFFFFFCC8;
      32'hFFFFFF03: r_cos = 32'hFFFFFCCD;
      32'hFFFFFF04: r_cos = 32'hFFFFFCD3;
      32'hFFFFFF05: r_cos = 32'hFFFFFCD9;
      32'hFFFFFF06: r_cos = 32'hFFFFFCDF;
      32'hFFFFFF07: r_cos = 32'hFFFFFCE5;
      32'hFFFFFF08: r_cos = 32'hFFFFFCEB;
      32'hFFFFFF09: r_cos = 32'hFFFFFCF1;
      32'hFFFFFF0A: r_cos = 32'hFFFFFCF7;
      32'hFFFFFF0B: r_cos = 32'hFFFFFCFE;
      32'hFFFFFF0C: r_cos = 32'hFFFFFD04;
      32'hFFFFFF0D: r_cos = 32'hFFFFFD0B;
      32'hFFFFFF0E: r_cos = 32'hFFFFFD11;
      32'hFFFFFF0F: r_cos = 32'hFFFFFD18;
      32'hFFFFFF10: r_cos = 32'hFFFFFD1F;
      32'hFFFFFF11: r_cos = 32'hFFFFFD25;
      32'hFFFFFF12: r_cos = 32'hFFFFFD2C;
      32'hFFFFFF13: r_cos = 32'hFFFFFD33;
      32'hFFFFFF14: r_cos = 32'hFFFFFD3A;
      32'hFFFFFF15: r_cos = 32'hFFFFFD41;
      32'hFFFFFF16: r_cos = 32'hFFFFFD48;
      32'hFFFFFF17: r_cos = 32'hFFFFFD50;
      32'hFFFFFF18: r_cos = 32'hFFFFFD57;
      32'hFFFFFF19: r_cos = 32'hFFFFFD5E;
      32'hFFFFFF1A: r_cos = 32'hFFFFFD66;
      32'hFFFFFF1B: r_cos = 32'hFFFFFD6D;
      32'hFFFFFF1C: r_cos = 32'hFFFFFD75;
      32'hFFFFFF1D: r_cos = 32'hFFFFFD7C;
      32'hFFFFFF1E: r_cos = 32'hFFFFFD84;
      32'hFFFFFF1F: r_cos = 32'hFFFFFD8C;
      32'hFFFFFF20: r_cos = 32'hFFFFFD94;
      32'hFFFFFF21: r_cos = 32'hFFFFFD9C;
      32'hFFFFFF22: r_cos = 32'hFFFFFDA3;
      32'hFFFFFF23: r_cos = 32'hFFFFFDAB;
      32'hFFFFFF24: r_cos = 32'hFFFFFDB3;
      32'hFFFFFF25: r_cos = 32'hFFFFFDBC;
      32'hFFFFFF26: r_cos = 32'hFFFFFDC4;
      32'hFFFFFF27: r_cos = 32'hFFFFFDCC;
      32'hFFFFFF28: r_cos = 32'hFFFFFDD4;
      32'hFFFFFF29: r_cos = 32'hFFFFFDDD;
      32'hFFFFFF2A: r_cos = 32'hFFFFFDE5;
      32'hFFFFFF2B: r_cos = 32'hFFFFFDED;
      32'hFFFFFF2C: r_cos = 32'hFFFFFDF6;
      32'hFFFFFF2D: r_cos = 32'hFFFFFDFF;
      32'hFFFFFF2E: r_cos = 32'hFFFFFE07;
      32'hFFFFFF2F: r_cos = 32'hFFFFFE10;
      32'hFFFFFF30: r_cos = 32'hFFFFFE19;
      32'hFFFFFF31: r_cos = 32'hFFFFFE21;
      32'hFFFFFF32: r_cos = 32'hFFFFFE2A;
      32'hFFFFFF33: r_cos = 32'hFFFFFE33;
      32'hFFFFFF34: r_cos = 32'hFFFFFE3C;
      32'hFFFFFF35: r_cos = 32'hFFFFFE45;
      32'hFFFFFF36: r_cos = 32'hFFFFFE4E;
      32'hFFFFFF37: r_cos = 32'hFFFFFE57;
      32'hFFFFFF38: r_cos = 32'hFFFFFE60;
      32'hFFFFFF39: r_cos = 32'hFFFFFE69;
      32'hFFFFFF3A: r_cos = 32'hFFFFFE72;
      32'hFFFFFF3B: r_cos = 32'hFFFFFE7B;
      32'hFFFFFF3C: r_cos = 32'hFFFFFE85;
      32'hFFFFFF3D: r_cos = 32'hFFFFFE8E;
      32'hFFFFFF3E: r_cos = 32'hFFFFFE97;
      32'hFFFFFF3F: r_cos = 32'hFFFFFEA0;
      32'hFFFFFF40: r_cos = 32'hFFFFFEAA;
      32'hFFFFFF41: r_cos = 32'hFFFFFEB3;
      32'hFFFFFF42: r_cos = 32'hFFFFFEBD;
      32'hFFFFFF43: r_cos = 32'hFFFFFEC6;
      32'hFFFFFF44: r_cos = 32'hFFFFFED0;
      32'hFFFFFF45: r_cos = 32'hFFFFFED9;
      32'hFFFFFF46: r_cos = 32'hFFFFFEE3;
      32'hFFFFFF47: r_cos = 32'hFFFFFEEC;
      32'hFFFFFF48: r_cos = 32'hFFFFFEF6;
      32'hFFFFFF49: r_cos = 32'hFFFFFF00;
      32'hFFFFFF4A: r_cos = 32'hFFFFFF09;
      32'hFFFFFF4B: r_cos = 32'hFFFFFF13;
      32'hFFFFFF4C: r_cos = 32'hFFFFFF1D;
      32'hFFFFFF4D: r_cos = 32'hFFFFFF27;
      32'hFFFFFF4E: r_cos = 32'hFFFFFF30;
      32'hFFFFFF4F: r_cos = 32'hFFFFFF3A;
      32'hFFFFFF50: r_cos = 32'hFFFFFF44;
      32'hFFFFFF51: r_cos = 32'hFFFFFF4E;
      32'hFFFFFF52: r_cos = 32'hFFFFFF58;
      32'hFFFFFF53: r_cos = 32'hFFFFFF61;
      32'hFFFFFF54: r_cos = 32'hFFFFFF6B;
      32'hFFFFFF55: r_cos = 32'hFFFFFF75;
      32'hFFFFFF56: r_cos = 32'hFFFFFF7F;
      32'hFFFFFF57: r_cos = 32'hFFFFFF89;
      32'hFFFFFF58: r_cos = 32'hFFFFFF93;
      32'hFFFFFF59: r_cos = 32'hFFFFFF9D;
      32'hFFFFFF5A: r_cos = 32'hFFFFFFA7;
      32'hFFFFFF5B: r_cos = 32'hFFFFFFB1;
      32'hFFFFFF5C: r_cos = 32'hFFFFFFBB;
      32'hFFFFFF5D: r_cos = 32'hFFFFFFC5;
      32'hFFFFFF5E: r_cos = 32'hFFFFFFCF;
      32'hFFFFFF5F: r_cos = 32'hFFFFFFD9;
      32'hFFFFFF60: r_cos = 32'hFFFFFFE3;
      32'hFFFFFF61: r_cos = 32'hFFFFFFED;
      32'hFFFFFF62: r_cos = 32'hFFFFFFF7;
      32'hFFFFFF63: r_cos = 32'h00000001;
      32'hFFFFFF64: r_cos = 32'h0000000B;
      32'hFFFFFF65: r_cos = 32'h00000015;
      32'hFFFFFF66: r_cos = 32'h0000001F;
      32'hFFFFFF67: r_cos = 32'h00000029;
      32'hFFFFFF68: r_cos = 32'h00000033;
      32'hFFFFFF69: r_cos = 32'h0000003D;
      32'hFFFFFF6A: r_cos = 32'h00000047;
      32'hFFFFFF6B: r_cos = 32'h00000051;
      32'hFFFFFF6C: r_cos = 32'h0000005B;
      32'hFFFFFF6D: r_cos = 32'h00000065;
      32'hFFFFFF6E: r_cos = 32'h0000006F;
      32'hFFFFFF6F: r_cos = 32'h00000079;
      32'hFFFFFF70: r_cos = 32'h00000082;
      32'hFFFFFF71: r_cos = 32'h0000008C;
      32'hFFFFFF72: r_cos = 32'h00000096;
      32'hFFFFFF73: r_cos = 32'h000000A0;
      32'hFFFFFF74: r_cos = 32'h000000AA;
      32'hFFFFFF75: r_cos = 32'h000000B4;
      32'hFFFFFF76: r_cos = 32'h000000BE;
      32'hFFFFFF77: r_cos = 32'h000000C7;
      32'hFFFFFF78: r_cos = 32'h000000D1;
      32'hFFFFFF79: r_cos = 32'h000000DB;
      32'hFFFFFF7A: r_cos = 32'h000000E5;
      32'hFFFFFF7B: r_cos = 32'h000000EE;
      32'hFFFFFF7C: r_cos = 32'h000000F8;
      32'hFFFFFF7D: r_cos = 32'h00000102;
      32'hFFFFFF7E: r_cos = 32'h0000010B;
      32'hFFFFFF7F: r_cos = 32'h00000115;
      32'hFFFFFF80: r_cos = 32'h0000011F;
      32'hFFFFFF81: r_cos = 32'h00000128;
      32'hFFFFFF82: r_cos = 32'h00000132;
      32'hFFFFFF83: r_cos = 32'h0000013B;
      32'hFFFFFF84: r_cos = 32'h00000145;
      32'hFFFFFF85: r_cos = 32'h0000014E;
      32'hFFFFFF86: r_cos = 32'h00000158;
      32'hFFFFFF87: r_cos = 32'h00000161;
      32'hFFFFFF88: r_cos = 32'h0000016A;
      32'hFFFFFF89: r_cos = 32'h00000174;
      32'hFFFFFF8A: r_cos = 32'h0000017D;
      32'hFFFFFF8B: r_cos = 32'h00000186;
      32'hFFFFFF8C: r_cos = 32'h0000018F;
      32'hFFFFFF8D: r_cos = 32'h00000198;
      32'hFFFFFF8E: r_cos = 32'h000001A2;
      32'hFFFFFF8F: r_cos = 32'h000001AB;
      32'hFFFFFF90: r_cos = 32'h000001B4;
      32'hFFFFFF91: r_cos = 32'h000001BD;
      32'hFFFFFF92: r_cos = 32'h000001C6;
      32'hFFFFFF93: r_cos = 32'h000001CE;
      32'hFFFFFF94: r_cos = 32'h000001D7;
      32'hFFFFFF95: r_cos = 32'h000001E0;
      32'hFFFFFF96: r_cos = 32'h000001E9;
      32'hFFFFFF97: r_cos = 32'h000001F2;
      32'hFFFFFF98: r_cos = 32'h000001FA;
      32'hFFFFFF99: r_cos = 32'h00000203;
      32'hFFFFFF9A: r_cos = 32'h0000020B;
      32'hFFFFFF9B: r_cos = 32'h00000214;
      32'hFFFFFF9C: r_cos = 32'h0000021C;
      32'hFFFFFF9D: r_cos = 32'h00000225;
      32'hFFFFFF9E: r_cos = 32'h0000022D;
      32'hFFFFFF9F: r_cos = 32'h00000235;
      32'hFFFFFFA0: r_cos = 32'h0000023E;
      32'hFFFFFFA1: r_cos = 32'h00000246;
      32'hFFFFFFA2: r_cos = 32'h0000024E;
      32'hFFFFFFA3: r_cos = 32'h00000256;
      32'hFFFFFFA4: r_cos = 32'h0000025E;
      32'hFFFFFFA5: r_cos = 32'h00000266;
      32'hFFFFFFA6: r_cos = 32'h0000026E;
      32'hFFFFFFA7: r_cos = 32'h00000275;
      32'hFFFFFFA8: r_cos = 32'h0000027D;
      32'hFFFFFFA9: r_cos = 32'h00000285;
      32'hFFFFFFAA: r_cos = 32'h0000028C;
      32'hFFFFFFAB: r_cos = 32'h00000294;
      32'hFFFFFFAC: r_cos = 32'h0000029B;
      32'hFFFFFFAD: r_cos = 32'h000002A3;
      32'hFFFFFFAE: r_cos = 32'h000002AA;
      32'hFFFFFFAF: r_cos = 32'h000002B1;
      32'hFFFFFFB0: r_cos = 32'h000002B9;
      32'hFFFFFFB1: r_cos = 32'h000002C0;
      32'hFFFFFFB2: r_cos = 32'h000002C7;
      32'hFFFFFFB3: r_cos = 32'h000002CE;
      32'hFFFFFFB4: r_cos = 32'h000002D5;
      32'hFFFFFFB5: r_cos = 32'h000002DC;
      32'hFFFFFFB6: r_cos = 32'h000002E2;
      32'hFFFFFFB7: r_cos = 32'h000002E9;
      32'hFFFFFFB8: r_cos = 32'h000002F0;
      32'hFFFFFFB9: r_cos = 32'h000002F6;
      32'hFFFFFFBA: r_cos = 32'h000002FD;
      32'hFFFFFFBB: r_cos = 32'h00000303;
      32'hFFFFFFBC: r_cos = 32'h0000030A;
      32'hFFFFFFBD: r_cos = 32'h00000310;
      32'hFFFFFFBE: r_cos = 32'h00000316;
      32'hFFFFFFBF: r_cos = 32'h0000031C;
      32'hFFFFFFC0: r_cos = 32'h00000322;
      32'hFFFFFFC1: r_cos = 32'h00000328;
      32'hFFFFFFC2: r_cos = 32'h0000032E;
      32'hFFFFFFC3: r_cos = 32'h00000334;
      32'hFFFFFFC4: r_cos = 32'h00000339;
      32'hFFFFFFC5: r_cos = 32'h0000033F;
      32'hFFFFFFC6: r_cos = 32'h00000344;
      32'hFFFFFFC7: r_cos = 32'h0000034A;
      32'hFFFFFFC8: r_cos = 32'h0000034F;
      32'hFFFFFFC9: r_cos = 32'h00000355;
      32'hFFFFFFCA: r_cos = 32'h0000035A;
      32'hFFFFFFCB: r_cos = 32'h0000035F;
      32'hFFFFFFCC: r_cos = 32'h00000364;
      32'hFFFFFFCD: r_cos = 32'h00000369;
      32'hFFFFFFCE: r_cos = 32'h0000036E;
      32'hFFFFFFCF: r_cos = 32'h00000372;
      32'hFFFFFFD0: r_cos = 32'h00000377;
      32'hFFFFFFD1: r_cos = 32'h0000037C;
      32'hFFFFFFD2: r_cos = 32'h00000380;
      32'hFFFFFFD3: r_cos = 32'h00000384;
      32'hFFFFFFD4: r_cos = 32'h00000389;
      32'hFFFFFFD5: r_cos = 32'h0000038D;
      32'hFFFFFFD6: r_cos = 32'h00000391;
      32'hFFFFFFD7: r_cos = 32'h00000395;
      32'hFFFFFFD8: r_cos = 32'h00000399;
      32'hFFFFFFD9: r_cos = 32'h0000039D;
      32'hFFFFFFDA: r_cos = 32'h000003A1;
      32'hFFFFFFDB: r_cos = 32'h000003A4;
      32'hFFFFFFDC: r_cos = 32'h000003A8;
      32'hFFFFFFDD: r_cos = 32'h000003AB;
      32'hFFFFFFDE: r_cos = 32'h000003AF;
      32'hFFFFFFDF: r_cos = 32'h000003B2;
      32'hFFFFFFE0: r_cos = 32'h000003B5;
      32'hFFFFFFE1: r_cos = 32'h000003B8;
      32'hFFFFFFE2: r_cos = 32'h000003BB;
      32'hFFFFFFE3: r_cos = 32'h000003BE;
      32'hFFFFFFE4: r_cos = 32'h000003C1;
      32'hFFFFFFE5: r_cos = 32'h000003C4;
      32'hFFFFFFE6: r_cos = 32'h000003C6;
      32'hFFFFFFE7: r_cos = 32'h000003C9;
      32'hFFFFFFE8: r_cos = 32'h000003CB;
      32'hFFFFFFE9: r_cos = 32'h000003CE;
      32'hFFFFFFEA: r_cos = 32'h000003D0;
      32'hFFFFFFEB: r_cos = 32'h000003D2;
      32'hFFFFFFEC: r_cos = 32'h000003D4;
      32'hFFFFFFED: r_cos = 32'h000003D6;
      32'hFFFFFFEE: r_cos = 32'h000003D8;
      32'hFFFFFFEF: r_cos = 32'h000003DA;
      32'hFFFFFFF0: r_cos = 32'h000003DB;
      32'hFFFFFFF1: r_cos = 32'h000003DD;
      32'hFFFFFFF2: r_cos = 32'h000003DE;
      32'hFFFFFFF3: r_cos = 32'h000003E0;
      32'hFFFFFFF4: r_cos = 32'h000003E1;
      32'hFFFFFFF5: r_cos = 32'h000003E2;
      32'hFFFFFFF6: r_cos = 32'h000003E3;
      32'hFFFFFFF7: r_cos = 32'h000003E4;
      32'hFFFFFFF8: r_cos = 32'h000003E5;
      32'hFFFFFFF9: r_cos = 32'h000003E6;
      32'hFFFFFFFA: r_cos = 32'h000003E6;
      32'hFFFFFFFB: r_cos = 32'h000003E7;
      32'hFFFFFFFC: r_cos = 32'h000003E7;
      32'hFFFFFFFD: r_cos = 32'h000003E8;
      32'hFFFFFFFE: r_cos = 32'h000003E8;
      32'hFFFFFFFF: r_cos = 32'h000003E8;
      32'h00000000: r_cos = 32'h000003E8;
      32'h00000001: r_cos = 32'h000003E8;
      32'h00000002: r_cos = 32'h000003E8;
      32'h00000003: r_cos = 32'h000003E8;
      32'h00000004: r_cos = 32'h000003E7;
      32'h00000005: r_cos = 32'h000003E7;
      32'h00000006: r_cos = 32'h000003E6;
      32'h00000007: r_cos = 32'h000003E6;
      32'h00000008: r_cos = 32'h000003E5;
      32'h00000009: r_cos = 32'h000003E4;
      32'h0000000A: r_cos = 32'h000003E3;
      32'h0000000B: r_cos = 32'h000003E2;
      32'h0000000C: r_cos = 32'h000003E1;
      32'h0000000D: r_cos = 32'h000003E0;
      32'h0000000E: r_cos = 32'h000003DE;
      32'h0000000F: r_cos = 32'h000003DD;
      32'h00000010: r_cos = 32'h000003DB;
      32'h00000011: r_cos = 32'h000003DA;
      32'h00000012: r_cos = 32'h000003D8;
      32'h00000013: r_cos = 32'h000003D6;
      32'h00000014: r_cos = 32'h000003D4;
      32'h00000015: r_cos = 32'h000003D2;
      32'h00000016: r_cos = 32'h000003D0;
      32'h00000017: r_cos = 32'h000003CE;
      32'h00000018: r_cos = 32'h000003CB;
      32'h00000019: r_cos = 32'h000003C9;
      32'h0000001A: r_cos = 32'h000003C6;
      32'h0000001B: r_cos = 32'h000003C4;
      32'h0000001C: r_cos = 32'h000003C1;
      32'h0000001D: r_cos = 32'h000003BE;
      32'h0000001E: r_cos = 32'h000003BB;
      32'h0000001F: r_cos = 32'h000003B8;
      32'h00000020: r_cos = 32'h000003B5;
      32'h00000021: r_cos = 32'h000003B2;
      32'h00000022: r_cos = 32'h000003AF;
      32'h00000023: r_cos = 32'h000003AB;
      32'h00000024: r_cos = 32'h000003A8;
      32'h00000025: r_cos = 32'h000003A4;
      32'h00000026: r_cos = 32'h000003A1;
      32'h00000027: r_cos = 32'h0000039D;
      32'h00000028: r_cos = 32'h00000399;
      32'h00000029: r_cos = 32'h00000395;
      32'h0000002A: r_cos = 32'h00000391;
      32'h0000002B: r_cos = 32'h0000038D;
      32'h0000002C: r_cos = 32'h00000389;
      32'h0000002D: r_cos = 32'h00000384;
      32'h0000002E: r_cos = 32'h00000380;
      32'h0000002F: r_cos = 32'h0000037C;
      32'h00000030: r_cos = 32'h00000377;
      32'h00000031: r_cos = 32'h00000372;
      32'h00000032: r_cos = 32'h0000036E;
      32'h00000033: r_cos = 32'h00000369;
      32'h00000034: r_cos = 32'h00000364;
      32'h00000035: r_cos = 32'h0000035F;
      32'h00000036: r_cos = 32'h0000035A;
      32'h00000037: r_cos = 32'h00000355;
      32'h00000038: r_cos = 32'h0000034F;
      32'h00000039: r_cos = 32'h0000034A;
      32'h0000003A: r_cos = 32'h00000344;
      32'h0000003B: r_cos = 32'h0000033F;
      32'h0000003C: r_cos = 32'h00000339;
      32'h0000003D: r_cos = 32'h00000334;
      32'h0000003E: r_cos = 32'h0000032E;
      32'h0000003F: r_cos = 32'h00000328;
      32'h00000040: r_cos = 32'h00000322;
      32'h00000041: r_cos = 32'h0000031C;
      32'h00000042: r_cos = 32'h00000316;
      32'h00000043: r_cos = 32'h00000310;
      32'h00000044: r_cos = 32'h0000030A;
      32'h00000045: r_cos = 32'h00000303;
      32'h00000046: r_cos = 32'h000002FD;
      32'h00000047: r_cos = 32'h000002F6;
      32'h00000048: r_cos = 32'h000002F0;
      32'h00000049: r_cos = 32'h000002E9;
      32'h0000004A: r_cos = 32'h000002E2;
      32'h0000004B: r_cos = 32'h000002DC;
      32'h0000004C: r_cos = 32'h000002D5;
      32'h0000004D: r_cos = 32'h000002CE;
      32'h0000004E: r_cos = 32'h000002C7;
      32'h0000004F: r_cos = 32'h000002C0;
      32'h00000050: r_cos = 32'h000002B9;
      32'h00000051: r_cos = 32'h000002B1;
      32'h00000052: r_cos = 32'h000002AA;
      32'h00000053: r_cos = 32'h000002A3;
      32'h00000054: r_cos = 32'h0000029B;
      32'h00000055: r_cos = 32'h00000294;
      32'h00000056: r_cos = 32'h0000028C;
      32'h00000057: r_cos = 32'h00000285;
      32'h00000058: r_cos = 32'h0000027D;
      32'h00000059: r_cos = 32'h00000275;
      32'h0000005A: r_cos = 32'h0000026E;
      32'h0000005B: r_cos = 32'h00000266;
      32'h0000005C: r_cos = 32'h0000025E;
      32'h0000005D: r_cos = 32'h00000256;
      32'h0000005E: r_cos = 32'h0000024E;
      32'h0000005F: r_cos = 32'h00000246;
      32'h00000060: r_cos = 32'h0000023E;
      32'h00000061: r_cos = 32'h00000235;
      32'h00000062: r_cos = 32'h0000022D;
      32'h00000063: r_cos = 32'h00000225;
      32'h00000064: r_cos = 32'h0000021C;
      32'h00000065: r_cos = 32'h00000214;
      32'h00000066: r_cos = 32'h0000020B;
      32'h00000067: r_cos = 32'h00000203;
      32'h00000068: r_cos = 32'h000001FA;
      32'h00000069: r_cos = 32'h000001F2;
      32'h0000006A: r_cos = 32'h000001E9;
      32'h0000006B: r_cos = 32'h000001E0;
      32'h0000006C: r_cos = 32'h000001D7;
      32'h0000006D: r_cos = 32'h000001CE;
      32'h0000006E: r_cos = 32'h000001C6;
      32'h0000006F: r_cos = 32'h000001BD;
      32'h00000070: r_cos = 32'h000001B4;
      32'h00000071: r_cos = 32'h000001AB;
      32'h00000072: r_cos = 32'h000001A2;
      32'h00000073: r_cos = 32'h00000198;
      32'h00000074: r_cos = 32'h0000018F;
      32'h00000075: r_cos = 32'h00000186;
      32'h00000076: r_cos = 32'h0000017D;
      32'h00000077: r_cos = 32'h00000174;
      32'h00000078: r_cos = 32'h0000016A;
      32'h00000079: r_cos = 32'h00000161;
      32'h0000007A: r_cos = 32'h00000158;
      32'h0000007B: r_cos = 32'h0000014E;
      32'h0000007C: r_cos = 32'h00000145;
      32'h0000007D: r_cos = 32'h0000013B;
      32'h0000007E: r_cos = 32'h00000132;
      32'h0000007F: r_cos = 32'h00000128;
      32'h00000080: r_cos = 32'h0000011F;
      32'h00000081: r_cos = 32'h00000115;
      32'h00000082: r_cos = 32'h0000010B;
      32'h00000083: r_cos = 32'h00000102;
      32'h00000084: r_cos = 32'h000000F8;
      32'h00000085: r_cos = 32'h000000EE;
      32'h00000086: r_cos = 32'h000000E5;
      32'h00000087: r_cos = 32'h000000DB;
      32'h00000088: r_cos = 32'h000000D1;
      32'h00000089: r_cos = 32'h000000C7;
      32'h0000008A: r_cos = 32'h000000BE;
      32'h0000008B: r_cos = 32'h000000B4;
      32'h0000008C: r_cos = 32'h000000AA;
      32'h0000008D: r_cos = 32'h000000A0;
      32'h0000008E: r_cos = 32'h00000096;
      32'h0000008F: r_cos = 32'h0000008C;
      32'h00000090: r_cos = 32'h00000082;
      32'h00000091: r_cos = 32'h00000079;
      32'h00000092: r_cos = 32'h0000006F;
      32'h00000093: r_cos = 32'h00000065;
      32'h00000094: r_cos = 32'h0000005B;
      32'h00000095: r_cos = 32'h00000051;
      32'h00000096: r_cos = 32'h00000047;
      32'h00000097: r_cos = 32'h0000003D;
      32'h00000098: r_cos = 32'h00000033;
      32'h00000099: r_cos = 32'h00000029;
      32'h0000009A: r_cos = 32'h0000001F;
      32'h0000009B: r_cos = 32'h00000015;
      32'h0000009C: r_cos = 32'h0000000B;
      32'h0000009D: r_cos = 32'h00000001;
      32'h0000009E: r_cos = 32'hFFFFFFF7;
      32'h0000009F: r_cos = 32'hFFFFFFED;
      32'h000000A0: r_cos = 32'hFFFFFFE3;
      32'h000000A1: r_cos = 32'hFFFFFFD9;
      32'h000000A2: r_cos = 32'hFFFFFFCF;
      32'h000000A3: r_cos = 32'hFFFFFFC5;
      32'h000000A4: r_cos = 32'hFFFFFFBB;
      32'h000000A5: r_cos = 32'hFFFFFFB1;
      32'h000000A6: r_cos = 32'hFFFFFFA7;
      32'h000000A7: r_cos = 32'hFFFFFF9D;
      32'h000000A8: r_cos = 32'hFFFFFF93;
      32'h000000A9: r_cos = 32'hFFFFFF89;
      32'h000000AA: r_cos = 32'hFFFFFF7F;
      32'h000000AB: r_cos = 32'hFFFFFF75;
      32'h000000AC: r_cos = 32'hFFFFFF6B;
      32'h000000AD: r_cos = 32'hFFFFFF61;
      32'h000000AE: r_cos = 32'hFFFFFF58;
      32'h000000AF: r_cos = 32'hFFFFFF4E;
      32'h000000B0: r_cos = 32'hFFFFFF44;
      32'h000000B1: r_cos = 32'hFFFFFF3A;
      32'h000000B2: r_cos = 32'hFFFFFF30;
      32'h000000B3: r_cos = 32'hFFFFFF27;
      32'h000000B4: r_cos = 32'hFFFFFF1D;
      32'h000000B5: r_cos = 32'hFFFFFF13;
      32'h000000B6: r_cos = 32'hFFFFFF09;
      32'h000000B7: r_cos = 32'hFFFFFF00;
      32'h000000B8: r_cos = 32'hFFFFFEF6;
      32'h000000B9: r_cos = 32'hFFFFFEEC;
      32'h000000BA: r_cos = 32'hFFFFFEE3;
      32'h000000BB: r_cos = 32'hFFFFFED9;
      32'h000000BC: r_cos = 32'hFFFFFED0;
      32'h000000BD: r_cos = 32'hFFFFFEC6;
      32'h000000BE: r_cos = 32'hFFFFFEBD;
      32'h000000BF: r_cos = 32'hFFFFFEB3;
      32'h000000C0: r_cos = 32'hFFFFFEAA;
      32'h000000C1: r_cos = 32'hFFFFFEA0;
      32'h000000C2: r_cos = 32'hFFFFFE97;
      32'h000000C3: r_cos = 32'hFFFFFE8E;
      32'h000000C4: r_cos = 32'hFFFFFE85;
      32'h000000C5: r_cos = 32'hFFFFFE7B;
      32'h000000C6: r_cos = 32'hFFFFFE72;
      32'h000000C7: r_cos = 32'hFFFFFE69;
      32'h000000C8: r_cos = 32'hFFFFFE60;
      32'h000000C9: r_cos = 32'hFFFFFE57;
      32'h000000CA: r_cos = 32'hFFFFFE4E;
      32'h000000CB: r_cos = 32'hFFFFFE45;
      32'h000000CC: r_cos = 32'hFFFFFE3C;
      32'h000000CD: r_cos = 32'hFFFFFE33;
      32'h000000CE: r_cos = 32'hFFFFFE2A;
      32'h000000CF: r_cos = 32'hFFFFFE21;
      32'h000000D0: r_cos = 32'hFFFFFE19;
      32'h000000D1: r_cos = 32'hFFFFFE10;
      32'h000000D2: r_cos = 32'hFFFFFE07;
      32'h000000D3: r_cos = 32'hFFFFFDFF;
      32'h000000D4: r_cos = 32'hFFFFFDF6;
      32'h000000D5: r_cos = 32'hFFFFFDED;
      32'h000000D6: r_cos = 32'hFFFFFDE5;
      32'h000000D7: r_cos = 32'hFFFFFDDD;
      32'h000000D8: r_cos = 32'hFFFFFDD4;
      32'h000000D9: r_cos = 32'hFFFFFDCC;
      32'h000000DA: r_cos = 32'hFFFFFDC4;
      32'h000000DB: r_cos = 32'hFFFFFDBC;
      32'h000000DC: r_cos = 32'hFFFFFDB3;
      32'h000000DD: r_cos = 32'hFFFFFDAB;
      32'h000000DE: r_cos = 32'hFFFFFDA3;
      32'h000000DF: r_cos = 32'hFFFFFD9C;
      32'h000000E0: r_cos = 32'hFFFFFD94;
      32'h000000E1: r_cos = 32'hFFFFFD8C;
      32'h000000E2: r_cos = 32'hFFFFFD84;
      32'h000000E3: r_cos = 32'hFFFFFD7C;
      32'h000000E4: r_cos = 32'hFFFFFD75;
      32'h000000E5: r_cos = 32'hFFFFFD6D;
      32'h000000E6: r_cos = 32'hFFFFFD66;
      32'h000000E7: r_cos = 32'hFFFFFD5E;
      32'h000000E8: r_cos = 32'hFFFFFD57;
      32'h000000E9: r_cos = 32'hFFFFFD50;
      32'h000000EA: r_cos = 32'hFFFFFD48;
      32'h000000EB: r_cos = 32'hFFFFFD41;
      32'h000000EC: r_cos = 32'hFFFFFD3A;
      32'h000000ED: r_cos = 32'hFFFFFD33;
      32'h000000EE: r_cos = 32'hFFFFFD2C;
      32'h000000EF: r_cos = 32'hFFFFFD25;
      32'h000000F0: r_cos = 32'hFFFFFD1F;
      32'h000000F1: r_cos = 32'hFFFFFD18;
      32'h000000F2: r_cos = 32'hFFFFFD11;
      32'h000000F3: r_cos = 32'hFFFFFD0B;
      32'h000000F4: r_cos = 32'hFFFFFD04;
      32'h000000F5: r_cos = 32'hFFFFFCFE;
      32'h000000F6: r_cos = 32'hFFFFFCF7;
      32'h000000F7: r_cos = 32'hFFFFFCF1;
      32'h000000F8: r_cos = 32'hFFFFFCEB;
      32'h000000F9: r_cos = 32'hFFFFFCE5;
      32'h000000FA: r_cos = 32'hFFFFFCDF;
      32'h000000FB: r_cos = 32'hFFFFFCD9;
      32'h000000FC: r_cos = 32'hFFFFFCD3;
      32'h000000FD: r_cos = 32'hFFFFFCCD;
      32'h000000FE: r_cos = 32'hFFFFFCC8;
      32'h000000FF: r_cos = 32'hFFFFFCC2;
      32'h00000100: r_cos = 32'hFFFFFCBC;
      32'h00000101: r_cos = 32'hFFFFFCB7;
      32'h00000102: r_cos = 32'hFFFFFCB2;
      32'h00000103: r_cos = 32'hFFFFFCAC;
      32'h00000104: r_cos = 32'hFFFFFCA7;
      32'h00000105: r_cos = 32'hFFFFFCA2;
      32'h00000106: r_cos = 32'hFFFFFC9D;
      32'h00000107: r_cos = 32'hFFFFFC98;
      32'h00000108: r_cos = 32'hFFFFFC93;
      32'h00000109: r_cos = 32'hFFFFFC8E;
      32'h0000010A: r_cos = 32'hFFFFFC8A;
      32'h0000010B: r_cos = 32'hFFFFFC85;
      32'h0000010C: r_cos = 32'hFFFFFC81;
      32'h0000010D: r_cos = 32'hFFFFFC7C;
      32'h0000010E: r_cos = 32'hFFFFFC78;
      32'h0000010F: r_cos = 32'hFFFFFC74;
      32'h00000110: r_cos = 32'hFFFFFC70;
      32'h00000111: r_cos = 32'hFFFFFC6C;
      32'h00000112: r_cos = 32'hFFFFFC68;
      32'h00000113: r_cos = 32'hFFFFFC64;
      32'h00000114: r_cos = 32'hFFFFFC60;
      32'h00000115: r_cos = 32'hFFFFFC5C;
      32'h00000116: r_cos = 32'hFFFFFC59;
      32'h00000117: r_cos = 32'hFFFFFC55;
      32'h00000118: r_cos = 32'hFFFFFC52;
      32'h00000119: r_cos = 32'hFFFFFC4E;
      32'h0000011A: r_cos = 32'hFFFFFC4B;
      32'h0000011B: r_cos = 32'hFFFFFC48;
      32'h0000011C: r_cos = 32'hFFFFFC45;
      32'h0000011D: r_cos = 32'hFFFFFC42;
      32'h0000011E: r_cos = 32'hFFFFFC3F;
      32'h0000011F: r_cos = 32'hFFFFFC3D;
      32'h00000120: r_cos = 32'hFFFFFC3A;
      32'h00000121: r_cos = 32'hFFFFFC37;
      32'h00000122: r_cos = 32'hFFFFFC35;
      32'h00000123: r_cos = 32'hFFFFFC33;
      32'h00000124: r_cos = 32'hFFFFFC30;
      32'h00000125: r_cos = 32'hFFFFFC2E;
      32'h00000126: r_cos = 32'hFFFFFC2C;
      32'h00000127: r_cos = 32'hFFFFFC2A;
      32'h00000128: r_cos = 32'hFFFFFC28;
      32'h00000129: r_cos = 32'hFFFFFC27;
      32'h0000012A: r_cos = 32'hFFFFFC25;
      32'h0000012B: r_cos = 32'hFFFFFC23;
      32'h0000012C: r_cos = 32'hFFFFFC22;
      32'h0000012D: r_cos = 32'hFFFFFC21;
      32'h0000012E: r_cos = 32'hFFFFFC1F;
      32'h0000012F: r_cos = 32'hFFFFFC1E;
      32'h00000130: r_cos = 32'hFFFFFC1D;
      32'h00000131: r_cos = 32'hFFFFFC1C;
      32'h00000132: r_cos = 32'hFFFFFC1B;
      32'h00000133: r_cos = 32'hFFFFFC1B;
      32'h00000134: r_cos = 32'hFFFFFC1A;
      32'h00000135: r_cos = 32'hFFFFFC19;
      32'h00000136: r_cos = 32'hFFFFFC19;
      32'h00000137: r_cos = 32'hFFFFFC18;
      32'h00000138: r_cos = 32'hFFFFFC18;
      32'h00000139: r_cos = 32'hFFFFFC18;
      32'h0000013A: r_cos = 32'hFFFFFC18;
      32'h0000013B: r_cos = 32'hFFFFFC18;
      32'h0000013C: r_cos = 32'hFFFFFC18;
      32'h0000013D: r_cos = 32'hFFFFFC18;
      32'h0000013E: r_cos = 32'hFFFFFC19;
      32'h0000013F: r_cos = 32'hFFFFFC19;
      32'h00000140: r_cos = 32'hFFFFFC1A;
      32'h00000141: r_cos = 32'hFFFFFC1A;
      32'h00000142: r_cos = 32'hFFFFFC1B;
      32'h00000143: r_cos = 32'hFFFFFC1C;
      32'h00000144: r_cos = 32'hFFFFFC1D;
      32'h00000145: r_cos = 32'hFFFFFC1E;
      32'h00000146: r_cos = 32'hFFFFFC1F;
      32'h00000147: r_cos = 32'hFFFFFC20;
      32'h00000148: r_cos = 32'hFFFFFC22;
      32'h00000149: r_cos = 32'hFFFFFC23;
      32'h0000014A: r_cos = 32'hFFFFFC25;
      32'h0000014B: r_cos = 32'hFFFFFC26;
      32'h0000014C: r_cos = 32'hFFFFFC28;
      32'h0000014D: r_cos = 32'hFFFFFC2A;
      32'h0000014E: r_cos = 32'hFFFFFC2C;
      32'h0000014F: r_cos = 32'hFFFFFC2E;
      32'h00000150: r_cos = 32'hFFFFFC30;
      32'h00000151: r_cos = 32'hFFFFFC32;
      32'h00000152: r_cos = 32'hFFFFFC34;
      32'h00000153: r_cos = 32'hFFFFFC37;
      32'h00000154: r_cos = 32'hFFFFFC39;
      32'h00000155: r_cos = 32'hFFFFFC3C;
      32'h00000156: r_cos = 32'hFFFFFC3F;
      32'h00000157: r_cos = 32'hFFFFFC41;
      32'h00000158: r_cos = 32'hFFFFFC44;
      32'h00000159: r_cos = 32'hFFFFFC47;
      32'h0000015A: r_cos = 32'hFFFFFC4A;
      32'h0000015B: r_cos = 32'hFFFFFC4D;
      32'h0000015C: r_cos = 32'hFFFFFC51;
      32'h0000015D: r_cos = 32'hFFFFFC54;
      32'h0000015E: r_cos = 32'hFFFFFC58;
      32'h0000015F: r_cos = 32'hFFFFFC5B;
      32'h00000160: r_cos = 32'hFFFFFC5F;
      32'h00000161: r_cos = 32'hFFFFFC62;
      32'h00000162: r_cos = 32'hFFFFFC66;
      32'h00000163: r_cos = 32'hFFFFFC6A;
      32'h00000164: r_cos = 32'hFFFFFC6E;
      32'h00000165: r_cos = 32'hFFFFFC72;
      32'h00000166: r_cos = 32'hFFFFFC77;
      32'h00000167: r_cos = 32'hFFFFFC7B;
      32'h00000168: r_cos = 32'hFFFFFC7F;
      32'h00000169: r_cos = 32'hFFFFFC84;
      32'h0000016A: r_cos = 32'hFFFFFC88;
      32'h0000016B: r_cos = 32'hFFFFFC8D;
      32'h0000016C: r_cos = 32'hFFFFFC92;
      32'h0000016D: r_cos = 32'hFFFFFC96;
      32'h0000016E: r_cos = 32'hFFFFFC9B;
      32'h0000016F: r_cos = 32'hFFFFFCA0;
      32'h00000170: r_cos = 32'hFFFFFCA5;
      32'h00000171: r_cos = 32'hFFFFFCAB;
      32'h00000172: r_cos = 32'hFFFFFCB0;
      32'h00000173: r_cos = 32'hFFFFFCB5;
      32'h00000174: r_cos = 32'hFFFFFCBB;
      32'h00000175: r_cos = 32'hFFFFFCC0;
      32'h00000176: r_cos = 32'hFFFFFCC6;
      32'h00000177: r_cos = 32'hFFFFFCCB;
      32'h00000178: r_cos = 32'hFFFFFCD1;
      32'h00000179: r_cos = 32'hFFFFFCD7;
      32'h0000017A: r_cos = 32'hFFFFFCDD;
      32'h0000017B: r_cos = 32'hFFFFFCE3;
      32'h0000017C: r_cos = 32'hFFFFFCE9;
      32'h0000017D: r_cos = 32'hFFFFFCEF;
      32'h0000017E: r_cos = 32'hFFFFFCF5;
      32'h0000017F: r_cos = 32'hFFFFFCFC;
      32'h00000180: r_cos = 32'hFFFFFD02;
      32'h00000181: r_cos = 32'hFFFFFD09;
      32'h00000182: r_cos = 32'hFFFFFD0F;
      32'h00000183: r_cos = 32'hFFFFFD16;
      32'h00000184: r_cos = 32'hFFFFFD1C;
      32'h00000185: r_cos = 32'hFFFFFD23;
      32'h00000186: r_cos = 32'hFFFFFD2A;
      32'h00000187: r_cos = 32'hFFFFFD31;
      32'h00000188: r_cos = 32'hFFFFFD38;
      32'h00000189: r_cos = 32'hFFFFFD3F;
      32'h0000018A: r_cos = 32'hFFFFFD46;
      32'h0000018B: r_cos = 32'hFFFFFD4D;
      32'h0000018C: r_cos = 32'hFFFFFD55;
      32'h0000018D: r_cos = 32'hFFFFFD5C;
      32'h0000018E: r_cos = 32'hFFFFFD63;
      32'h0000018F: r_cos = 32'hFFFFFD6B;
      32'h00000190: r_cos = 32'hFFFFFD72;
      32'h00000191: r_cos = 32'hFFFFFD7A;
      32'h00000192: r_cos = 32'hFFFFFD82;
      32'h00000193: r_cos = 32'hFFFFFD89;
      32'h00000194: r_cos = 32'hFFFFFD91;
      32'h00000195: r_cos = 32'hFFFFFD99;
      32'h00000196: r_cos = 32'hFFFFFDA1;
      32'h00000197: r_cos = 32'hFFFFFDA9;
      32'h00000198: r_cos = 32'hFFFFFDB1;
      32'h00000199: r_cos = 32'hFFFFFDB9;
      32'h0000019A: r_cos = 32'hFFFFFDC1;
      32'h0000019B: r_cos = 32'hFFFFFDC9;
      32'h0000019C: r_cos = 32'hFFFFFDD2;
      32'h0000019D: r_cos = 32'hFFFFFDDA;
      32'h0000019E: r_cos = 32'hFFFFFDE2;
      32'h0000019F: r_cos = 32'hFFFFFDEB;
      32'h000001A0: r_cos = 32'hFFFFFDF3;
      32'h000001A1: r_cos = 32'hFFFFFDFC;
      32'h000001A2: r_cos = 32'hFFFFFE04;
      32'h000001A3: r_cos = 32'hFFFFFE0D;
      32'h000001A4: r_cos = 32'hFFFFFE16;
      32'h000001A5: r_cos = 32'hFFFFFE1E;
      32'h000001A6: r_cos = 32'hFFFFFE27;
      32'h000001A7: r_cos = 32'hFFFFFE30;
      32'h000001A8: r_cos = 32'hFFFFFE39;
      32'h000001A9: r_cos = 32'hFFFFFE42;
      32'h000001AA: r_cos = 32'hFFFFFE4B;
      32'h000001AB: r_cos = 32'hFFFFFE54;
      32'h000001AC: r_cos = 32'hFFFFFE5D;
      32'h000001AD: r_cos = 32'hFFFFFE66;
      32'h000001AE: r_cos = 32'hFFFFFE6F;
      32'h000001AF: r_cos = 32'hFFFFFE78;
      32'h000001B0: r_cos = 32'hFFFFFE82;
      32'h000001B1: r_cos = 32'hFFFFFE8B;
      32'h000001B2: r_cos = 32'hFFFFFE94;
      32'h000001B3: r_cos = 32'hFFFFFE9D;
      32'h000001B4: r_cos = 32'hFFFFFEA7;
      32'h000001B5: r_cos = 32'hFFFFFEB0;
      32'h000001B6: r_cos = 32'hFFFFFEBA;
      32'h000001B7: r_cos = 32'hFFFFFEC3;
      32'h000001B8: r_cos = 32'hFFFFFECD;
      32'h000001B9: r_cos = 32'hFFFFFED6;
      32'h000001BA: r_cos = 32'hFFFFFEE0;
      32'h000001BB: r_cos = 32'hFFFFFEE9;
      32'h000001BC: r_cos = 32'hFFFFFEF3;
      32'h000001BD: r_cos = 32'hFFFFFEFD;
      32'h000001BE: r_cos = 32'hFFFFFF06;
      32'h000001BF: r_cos = 32'hFFFFFF10;
      32'h000001C0: r_cos = 32'hFFFFFF1A;
      32'h000001C1: r_cos = 32'hFFFFFF23;
      32'h000001C2: r_cos = 32'hFFFFFF2D;
      32'h000001C3: r_cos = 32'hFFFFFF37;
      32'h000001C4: r_cos = 32'hFFFFFF41;
      32'h000001C5: r_cos = 32'hFFFFFF4B;
      32'h000001C6: r_cos = 32'hFFFFFF54;
      32'h000001C7: r_cos = 32'hFFFFFF5E;
      32'h000001C8: r_cos = 32'hFFFFFF68;
      32'h000001C9: r_cos = 32'hFFFFFF72;
      32'h000001CA: r_cos = 32'hFFFFFF7C;
      32'h000001CB: r_cos = 32'hFFFFFF86;
      32'h000001CC: r_cos = 32'hFFFFFF90;
      32'h000001CD: r_cos = 32'hFFFFFF9A;
      32'h000001CE: r_cos = 32'hFFFFFFA4;
      32'h000001CF: r_cos = 32'hFFFFFFAE;
      32'h000001D0: r_cos = 32'hFFFFFFB8;
      32'h000001D1: r_cos = 32'hFFFFFFC2;
      32'h000001D2: r_cos = 32'hFFFFFFCC;
      32'h000001D3: r_cos = 32'hFFFFFFD6;
      32'h000001D4: r_cos = 32'hFFFFFFE0;
      32'h000001D5: r_cos = 32'hFFFFFFEA;
      32'h000001D6: r_cos = 32'hFFFFFFF4;
      32'h000001D7: r_cos = 32'hFFFFFFFE;
      32'h000001D8: r_cos = 32'h00000008;
      32'h000001D9: r_cos = 32'h00000012;
      32'h000001DA: r_cos = 32'h0000001C;
      32'h000001DB: r_cos = 32'h00000026;
      32'h000001DC: r_cos = 32'h00000030;
      32'h000001DD: r_cos = 32'h0000003A;
      32'h000001DE: r_cos = 32'h00000044;
      32'h000001DF: r_cos = 32'h0000004E;
      32'h000001E0: r_cos = 32'h00000057;
      32'h000001E1: r_cos = 32'h00000061;
      32'h000001E2: r_cos = 32'h0000006B;
      32'h000001E3: r_cos = 32'h00000075;
      32'h000001E4: r_cos = 32'h0000007F;
      32'h000001E5: r_cos = 32'h00000089;
      32'h000001E6: r_cos = 32'h00000093;
      32'h000001E7: r_cos = 32'h0000009D;
      32'h000001E8: r_cos = 32'h000000A7;
      32'h000001E9: r_cos = 32'h000000B1;
      32'h000001EA: r_cos = 32'h000000BB;
      32'h000001EB: r_cos = 32'h000000C4;
      32'h000001EC: r_cos = 32'h000000CE;
      32'h000001ED: r_cos = 32'h000000D8;
      32'h000001EE: r_cos = 32'h000000E2;
      32'h000001EF: r_cos = 32'h000000EB;
      32'h000001F0: r_cos = 32'h000000F5;
      32'h000001F1: r_cos = 32'h000000FF;
      32'h000001F2: r_cos = 32'h00000108;
      32'h000001F3: r_cos = 32'h00000112;
      32'h000001F4: r_cos = 32'h0000011C;
      32'h000001F5: r_cos = 32'h00000125;
      32'h000001F6: r_cos = 32'h0000012F;
      32'h000001F7: r_cos = 32'h00000138;
      32'h000001F8: r_cos = 32'h00000142;
      32'h000001F9: r_cos = 32'h0000014B;
      32'h000001FA: r_cos = 32'h00000155;
      32'h000001FB: r_cos = 32'h0000015E;
      32'h000001FC: r_cos = 32'h00000167;
      32'h000001FD: r_cos = 32'h00000171;
      32'h000001FE: r_cos = 32'h0000017A;
      32'h000001FF: r_cos = 32'h00000183;
      32'h00000200: r_cos = 32'h0000018C;
      32'h00000201: r_cos = 32'h00000196;
      32'h00000202: r_cos = 32'h0000019F;
      32'h00000203: r_cos = 32'h000001A8;
      32'h00000204: r_cos = 32'h000001B1;
      32'h00000205: r_cos = 32'h000001BA;
      32'h00000206: r_cos = 32'h000001C3;
      32'h00000207: r_cos = 32'h000001CC;
      32'h00000208: r_cos = 32'h000001D5;
      32'h00000209: r_cos = 32'h000001DD;
      32'h0000020A: r_cos = 32'h000001E6;
      32'h0000020B: r_cos = 32'h000001EF;
      32'h0000020C: r_cos = 32'h000001F7;
      32'h0000020D: r_cos = 32'h00000200;
      32'h0000020E: r_cos = 32'h00000209;
      32'h0000020F: r_cos = 32'h00000211;
      32'h00000210: r_cos = 32'h0000021A;
      32'h00000211: r_cos = 32'h00000222;
      32'h00000212: r_cos = 32'h0000022A;
      32'h00000213: r_cos = 32'h00000233;
      32'h00000214: r_cos = 32'h0000023B;
      32'h00000215: r_cos = 32'h00000243;
      32'h00000216: r_cos = 32'h0000024B;
      32'h00000217: r_cos = 32'h00000253;
      32'h00000218: r_cos = 32'h0000025B;
      32'h00000219: r_cos = 32'h00000263;
      32'h0000021A: r_cos = 32'h0000026B;
      32'h0000021B: r_cos = 32'h00000273;
      32'h0000021C: r_cos = 32'h0000027B;
      32'h0000021D: r_cos = 32'h00000282;
      32'h0000021E: r_cos = 32'h0000028A;
      32'h0000021F: r_cos = 32'h00000292;
      32'h00000220: r_cos = 32'h00000299;
      32'h00000221: r_cos = 32'h000002A1;
      32'h00000222: r_cos = 32'h000002A8;
      32'h00000223: r_cos = 32'h000002AF;
      32'h00000224: r_cos = 32'h000002B6;
      32'h00000225: r_cos = 32'h000002BE;
      32'h00000226: r_cos = 32'h000002C5;
      32'h00000227: r_cos = 32'h000002CC;
      32'h00000228: r_cos = 32'h000002D3;
      32'h00000229: r_cos = 32'h000002DA;
      32'h0000022A: r_cos = 32'h000002E0;
      32'h0000022B: r_cos = 32'h000002E7;
      32'h0000022C: r_cos = 32'h000002EE;
      32'h0000022D: r_cos = 32'h000002F4;
      32'h0000022E: r_cos = 32'h000002FB;
      32'h0000022F: r_cos = 32'h00000301;
      32'h00000230: r_cos = 32'h00000308;
      32'h00000231: r_cos = 32'h0000030E;
      32'h00000232: r_cos = 32'h00000314;
      32'h00000233: r_cos = 32'h0000031A;
      32'h00000234: r_cos = 32'h00000320;
      32'h00000235: r_cos = 32'h00000326;
      32'h00000236: r_cos = 32'h0000032C;
      32'h00000237: r_cos = 32'h00000332;
      32'h00000238: r_cos = 32'h00000338;
      32'h00000239: r_cos = 32'h0000033D;
      32'h0000023A: r_cos = 32'h00000343;
      32'h0000023B: r_cos = 32'h00000348;
      32'h0000023C: r_cos = 32'h0000034E;
      32'h0000023D: r_cos = 32'h00000353;
      32'h0000023E: r_cos = 32'h00000358;
      32'h0000023F: r_cos = 32'h0000035D;
      32'h00000240: r_cos = 32'h00000362;
      32'h00000241: r_cos = 32'h00000367;
      32'h00000242: r_cos = 32'h0000036C;
      32'h00000243: r_cos = 32'h00000371;
      32'h00000244: r_cos = 32'h00000376;
      32'h00000245: r_cos = 32'h0000037A;
      32'h00000246: r_cos = 32'h0000037F;
      32'h00000247: r_cos = 32'h00000383;
      32'h00000248: r_cos = 32'h00000387;
      32'h00000249: r_cos = 32'h0000038C;
      32'h0000024A: r_cos = 32'h00000390;
      32'h0000024B: r_cos = 32'h00000394;
      32'h0000024C: r_cos = 32'h00000398;
      32'h0000024D: r_cos = 32'h0000039C;
      32'h0000024E: r_cos = 32'h0000039F;
      32'h0000024F: r_cos = 32'h000003A3;
      32'h00000250: r_cos = 32'h000003A7;
      32'h00000251: r_cos = 32'h000003AA;
      32'h00000252: r_cos = 32'h000003AE;
      32'h00000253: r_cos = 32'h000003B1;
      32'h00000254: r_cos = 32'h000003B4;
      32'h00000255: r_cos = 32'h000003B7;
      32'h00000256: r_cos = 32'h000003BA;
      32'h00000257: r_cos = 32'h000003BD;
      32'h00000258: r_cos = 32'h000003C0;
      32'h00000259: r_cos = 32'h000003C3;
      32'h0000025A: r_cos = 32'h000003C6;
      32'h0000025B: r_cos = 32'h000003C8;
      32'h0000025C: r_cos = 32'h000003CB;
      32'h0000025D: r_cos = 32'h000003CD;
      32'h0000025E: r_cos = 32'h000003CF;
      32'h0000025F: r_cos = 32'h000003D1;
      32'h00000260: r_cos = 32'h000003D3;
      32'h00000261: r_cos = 32'h000003D5;
      32'h00000262: r_cos = 32'h000003D7;
      32'h00000263: r_cos = 32'h000003D9;
      32'h00000264: r_cos = 32'h000003DB;
      32'h00000265: r_cos = 32'h000003DC;
      32'h00000266: r_cos = 32'h000003DE;
      32'h00000267: r_cos = 32'h000003DF;
      32'h00000268: r_cos = 32'h000003E0;
      32'h00000269: r_cos = 32'h000003E2;
      32'h0000026A: r_cos = 32'h000003E3;
      32'h0000026B: r_cos = 32'h000003E4;
      32'h0000026C: r_cos = 32'h000003E5;
      32'h0000026D: r_cos = 32'h000003E5;
      32'h0000026E: r_cos = 32'h000003E6;
      32'h0000026F: r_cos = 32'h000003E7;
      32'h00000270: r_cos = 32'h000003E7;
      32'h00000271: r_cos = 32'h000003E7;
      32'h00000272: r_cos = 32'h000003E8;
      32'h00000273: r_cos = 32'h000003E8;
      32'h00000274: r_cos = 32'h000003E8;
      default: r_cos = 32'h00000000;
endcase

end


endmodule