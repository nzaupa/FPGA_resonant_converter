// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 15:05:49 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aMatLLfKUPCBwB6Z5+r8yOg6fkG7LzVMLxKNr5WedmPDfWeFp5XadQ/G7YyxnqhP
YhQhkVVF8OrhqLGF7VyOhD/CVsXdlQ+waUPdeQ61/sV1Miz2oB394EasLSst86XY
bl+JJH/C1Ayv9arKFjK8FyOxkj/ywEJeUpZ7vf/vHFs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9088)
8cCWZmJXvsxcGWRJeo8ZuBMSeYYGsRNB+54KoFG/ou1qQRRQcJV7v4Vp68m7Z9dp
NwM9XmUQntw6Fs60vNkv5K2n9v34t8VI4NCxV6BOHrcDOr2ofZNIDfR3qSogIzUs
c7jDXPtSW4TZzRhNk0zDKxgfP1RKuMpdiiC2KJWUQmmTXoQ3A/0SAhsXAlLdoJf1
3Bz+LKAOLjqlPziqwhbJ3DXcCtFt8NLGePTTeY+ZaGb2wATkR9S+F3OPc/5vRJEv
Sjg+MtIZIZPQR+F2YNWA8nmd0eEQu5kxVjuQJMPYGL44M18JziqoyhoLPtGgRntH
68Zq5/f8Xbe0+jiU7+Emkmvfv7MMJG/LtUOvEqXO8moL0kxDaaZHKkX0Ix0Yoa03
oaXtdwa6gYLHvxk8SX5+3vypw0j/5/KnEZV78P3Aa06uqL5nO5wkFNXHRj8+l2Jh
82URIf6H5ojXKWSpF6vIyVfScClzlMePG95AdbzOwr0HfyTqHjFH5zWMWv8BStlE
hs+uVnjJXwDvcvbYkXL4PnuCYmnaeVlS9TWb+Nu01GySjk+G0/24nY2oxQLUqiDy
wonGBpfsiPsz7+i/b9raQxYj/pnQyaGvXX8bMU/kqCdUVNssphR/vbgPnRjIoE24
NvddGuIs9LYSHjN2NTZ02e/A+nKnKw5wqMsB1HY2eui6E6k3U45RTe3vQ2+/6z/I
1/7b2Oam7CjraYqKFJwgKE5JbdoCguz1tTmfTm5LlhU5scG98cZrUsKotsZZcXRJ
VjuCFOJpBvYMuGbOd4p8N0YAIGJEDC+ZjfcA39KaIz7Lsd6a+jx+p8SHQ/M9jdsB
UbtT7yF9ydrYOi6wbRl8okiy62SuH/Hcjhgv6FRvzovW/2ozyYF/EZeJNLO5adh2
CEb0bKRHV1jNw64fE0+FMUsp1GAtDDDQHqhdKvYQgkSJRl144CIrVoMO8d8IrOce
Ui9Wght26zQYA7sYJ6VIHbHc7G4ig+XA9B79+8g8eVzLZE1swC/ov0ucjfp9MHAZ
QCbfHxyJMoi6UfT8dyPPxSVCdOQMdWeopRs3u5C+s4A0eZDck91D/t4b0ZYD020L
6MqYB1yqopp3FNqPp39RAkxsB20Zy2IEd5NczH2cQprkfjwTy0DvBNXBxqT6Yqyk
xNpRqf1p/ZvrSKwvGDwwoAT4iTXl2x55AMUzzaancIpBw9y2hs8U85ZquwFF7hC9
zjiyPRnGlep/PTtatZwJ1pD1OH7mZaix3oMRfdram1PCicb2TVEJFVRi9GzB09H3
ahdDg19NwjnKqNzvEkZ9Afh5F9QP7mgwVpXBaYwQP+lJwTplnjSRKmtqmz5zcbKq
TtGn4v400qP8rjCZzD8GY1NNYIpk2edCleua+D86e25afuQpW9a3uTGFAkl/hq49
hjyoFrguKQcrkcBNDV2exlQfOUh5ROtbif/LjyC91P+qeBeAhLfaJe6CLhkFBvUf
CJkbWKMAdlYG45kiQdR9OoTQDGuAcHWbnuc/hYwqFtv9AuSpp6XEyjGMrYJOT7Mr
KpEzAD0R+w95zB7SnU8Cjf2ZVjGG7T9MIEnPi4pbeYCFWWKpeR/KQlp5Wbc1trgI
T3j19OqyNhFT9+V8EjnVeB5FShJv4ltIaeW6cDJ0hPxCv11VqU4yheZP7tFMViyk
F4GKf02QMxxp1I53fbPXWXgR6aKtvXPevRC1xl7iyjswAbW8UIXRR2bQlN1wdyus
Oc+3/XfzS5TEIPUOQKNUNiUYft91BQJgOIT+1k5L9e2bsGVWFmjWGQ6LNq2yOhOi
jyvxSIk6rB2xeSuU1u3QkcnbBUDjcFcvqZxxZpsge6c93AxzaDNjEXgHJeEJs7qm
nMbDr4MnOmrqr4U7WATap0nT7lFtrBGGiyvfKMp7hsBQvC+IbR7g4OwFx8ZSCFfQ
p1ZRuCbagwlgPtJrqNjHKem2rmth0Aqcu0vnoMF0JHW4/b2bsxMUK7fxAdgsYK2Q
gR6fpt1WBnRXYM4Nh25S4vI6ntQ14sVrtMlDVZA8VKRKuLo33nalNU3kHqhvLurr
krTxRsh2SPb+DyMdVLTummRi4PemIQ3m14cZCH4jvxKk6ZLF/OHwRrBVxAEP+oQ3
hyyPU3Kgdjz6nVxQSFrSMEhFMMZk5lyba6gyLqdGqdIfMkCXojWhAOBeQSrk4X5P
MyrcFFHDtx8Ps1yGDEf4faSvv/PJTeabZyQx9Sp1VRJsxrQ4avf9TophoJrRP2lt
NenuFZmeAJS90pwYHxLkwhxHO1c9TMxRRWBaavQ8FW0vqUnWTcdlwublR1L8WHsg
mqOaxsECNqwXiue+21pcpblEA9nwz3+9zjGC13sjP50+TbPk/yCZWFhqBQDs0a7I
jbWBekTeS5VQ6NwpvmF6hylVTSvrQOgjFbAQ4RdNPTP8m2wixXP3vzke2vJPvuAV
VrFnBq6vMwSaApS3V7gZBKUma3YyVU4XDOGDonRsI30vbEuLF+l0Jz2DHsCoj9UQ
4oxGJ7LTNI4Vs95aAiPEfhKDrBTcP0VhiuDrWxZdbLJZ1u9LJ+GnvQGSp+fXhw7L
BTyRmAw3B8JI/uSIunNwrI5PbSoi5n2HehGRyu20NPq2iAM01y0fXgIrpGdPPbdP
bRHG1GQuwgIe/JQFlgnTD0ORYhCaqsXVNrRgMd6Lnvl00nHHbOY4ai6nTqFryBFU
Jo4Rr4M2OdVSYmvh4ONX0P3IjUqQHXzFh2rbIweYQ/jNxpZwPTWpm3AFi6W8kj11
736NjZBVhUsgkzt8M6rNdutCPqju4Qm9HoX2XQiW5ZuH4JyY3Vhd6Ied+1Qy370m
+mwDAVCDerZHIf4y4gxTQUDAfMDkHDxQ8Kl8V+fu7S+3UOePsGn2VYh0aPNuA7Hm
+58KEI/lAxR9NYZjaFax/wr8+rpYaPI+wkIQ3WfdJaEVGEetv01XNNlG428MiPLn
Vaa65v3rSYpGhhS+FZjqDCL15FtNsar0lsEoqzzat38vQj6s6hJ2Qs9oON1TiFUs
b0JudKUJkiLptcVk6vRlPFbHGsGjLgXsiY1bVb94FJCq4NGd9GyPP2Lixgcjuwcl
2ODI8X70ssp6Z2x+6OZvaaIL3P0hJL5aTfNK2CsQ99YO1GBc6wKgPCKFVtq7qYvg
CZO2gLLOmLLNFP6vbTqArCjLKxJZNMI75j+DU8oYjYCq1gRrFY3ZwzLFnFHblcCT
EMHYfqHind3X6ySeT+M8zJ41Ew3dXof4aQv/mFJVLdFca8HgpZ9Ra3/bLtAr83q6
qjYbDeaKUAWmNwfN/983EolD8ordUKuVpajW/PwbjPlyWcz6bio7WPIAdAbzDtiG
kNbQ4Qb1luuD8vfZNrY6r6dgReO31H9YpVxEuhTP/gFKjdzFbrG2Y1xizKkFNWY0
FYvMOoQOWs2vFU8yol2KZcBQ8+t+bwxgT7Bnkg+01kPbcdIyf45cYwlkctVHiQVo
mGtQFa9UdTj2cpKzgx8Kz77C2+0J9PkPdndklAnlh/BkeS05XNhW8UMqfnxcPYbh
qrk+IfWSXoZIEJirDOwiISZ4YWwlnZh4UltZ7n+BpsQmhgfgMPW67N7bTSS6d8pf
58CwxpWS4ClDTUcQl4c/NbLRIITXFjgEgRgzYrSStqGfZEnbbZL0aRGdiKj3whpa
CXhF8qNsTPvSvp4Ozm5yfPo/Qs/7X2ZLVJdc9kYDnaShiWLP5gsOEODZq803/Mup
POkHpJFpVkXSjTGdhBl0meWRrFzYdj8L8MwI+r1hXi5mVeORDMNeQPM6M9xODl67
Bm++KOQkXmjE49HPC2tGF+tLtThfg9wGxRMBgGwOtHT4czG1ZnOnVqWNRblxUbEi
yQGTOuIGC+kcVlOBkMLWFw8JiuJHFXmxxAtADuBNjiKIsPDQU/P6xK9+6XKoCb97
UvF0pp6Ac+fG3NFFmnTtMziSeazXwLjlxkkpFubeaHxEKgzl54Xjq2OwEAcFgxFV
1kYTOCfGGiZwThEHkO+x4V7Aa4vk6ZssZZJ0UwFD2qdgsYBW9oj98alofY1hSMBm
LltL35hGaTXKSFlK80WP3lURG6CKU630PbmdbXuZfInGuttvs5VjW9gelnwYVK+f
CFIr6hVlfYv5Sv3wvJIldeuN7KuKErGLy0YmKSgP+YwFZZ45VK2/xO2JNSdHWTLz
2CL7GNjAA4Hls2epJIyNhCpbruUSV4nZYo6odzO29gAYW0g/5TY4/uxm2X6fZV0a
FFuAHcE35SJAeLgfa9G0rJWb2cA9opwgE1NiryLzpqa9t83mm+AKmFDy6epfpQeG
PzeAau35H/N3QbiqEEdPwFjU+QUaCkiFXX2B7P8EsSRLY5c+IGnlDTX6FWjP2fRJ
Aa3fClOhku2LIkPu+jfydehYwLRJSVnqQG8pLKIhfyL1sDBC63CaRS6Pjyla6cpO
ggdznOYhXE8K9xdlLoNYJbOmiNC+RlH34iDYtLtX4xNPRGujEo2pll0ZmM1jTlm2
i/IJQaF0iBVPQ3SflUp+qEDKKSKWFbmdS28FLm/DJSnCX3GWCqQG3kJiOdcC3Dts
gjQvgAU3E2tfTZ0rsGeOZBI0uuZhPLIafoBC7taVdK+6k2b2ChPWFgJOA9kmF8/l
7K7WvdBGw6s69QhqzZwWO6a1f6HoFGAlXYT2MYj4iySLYInpOtKOYq6zdJnJ7nb7
C34wybB7NyOvoA/1yUSAWwaG0pCGB0ctcfltI8IVVsbU2/wvQVI+Ia35n3X82pWW
swzqqO4Glvt3zpAQ0U3DiU7dbtbcS+MhOG+hL2HUuOcRDYJ7dbFnO4eqBT/8UN0a
RVrGokWBao0/RJ5tXRNYkGQflLzj3gIyHDIeUED5Ms+GaAPBSoqEdUqkNxBMQQr0
zOKsRBz+tKWCDNUP/vZ07tjYr/P5+L4rmyurplJZE4fmi5lNr7h6SV1GcYSLTADR
c0UMVWD4yOhkuKks+SGvJTmOy0Divuuv22w6EFuPDyXk+DWqOh7Ce20lL62Mu+/z
o8Pu6VIlSsAK1gw1NwWoQoXnF2qTD0T6/0WU21HKvOaRFh56KGq8DehKehdCAFhg
BAIJVC2gIuA5YnssRGwdnyAvMDY9/bW44b7n+QdfNpIb2tC9XvrvAgrmGwaI2KBS
wSVZu/T8jhH+QRs/ZLCsp02+0pgnUsqCZKtI5xnFsdPwpxFEAzxcWZ2pq1N38F1i
4kb4OfoGFroRaBZaZExyAwKx1pcizgD7pXfa4PLHXBK2wn9kqPCmnZeViydr6LfA
qIjjzXAIEI96vYvVQUUrlNaTouRmlkXjozQT+BfCipHsxZR6wzeRdkq5BdZOqXGo
NOipqzP6wy5huSEFghohdDVY3RE8Z+XQO3g/C9FGds9ViEYKFH+ZQV8MyKQ3kAYn
yuHhzH3bOTiXX5GuA2cX/9K7wkll5b6LIXGMjP1lgrypImHu7SHxSP3el710dP43
OFn+DlRdb22W95YfRsCc1DJACG4C0S17O0Dr2VIgUkpDrNi1PCcuYaX7AfMTJtNl
FMktI2YD/gvDLKQ3lg5UxqI7YeUkVyjxHgb3yJotku0D+OKe1k7gFEgWNRKWBUYu
C57ie80/wmmigASw6+U+gV8SB8Pdx2uPnPncGsJxg1s3HC43cl2ziB0Esy5YZ8Tl
+ZERF+ge77gH1emiVXjSJ4ViAyn0eap8dOqNR0g8yzwTFAmyIQRA0r9BHEB2Hs11
ttVIxkDBdTCGX8uPMJ0pAxfpf/SvwIfeQuJcECCfcYxMz4/2rAMjz4utN9gOE05y
j18EYRP8pVZylBZm/QxLvF4ox0VeRmdVNMs5wkKhbE7vggoCWDzYcvLAF450NSkJ
iXxbWniL/9sCla/X7M1bk3O6oo0QREIiJyvSW6fuxUB5vSb5S2BoTzMcRSF1vyQu
QnDwXXIhf26Yg6cmi5W3P9Il6E6SX1DIK/hD07W9I5Jxm2v4HP3WU8xyyL8hm6sm
t+QjnLBzkHkX7NjtnITzXUX2VQsbhBDOh8hrSyzNZuXTq+E2H+fC3cz4veKE5xIr
GTH+3QfiMBx1Tt8Ell0jaYmuh2ArAPFIemAGZV+p+gQXm1017KCWnpNQOpdiyRSI
/VkzExoR5uoijpZQ3eqEGfMz1cEdXvRjFzpq2yotL0IHeAnPCSo30H37IQEkMIuk
TiI4lt5m7vzdvYHnd+8j4kOY1qeZ07eYzGEWMKmOvSi6tNGXoXF9yi4oszQIeCKC
MKI66Ndz7t2i3s9zLB613ol+Z4zPSKqsPvi1udQfgimG4XkyhikPPs42NmBSwdI0
VZH9XAJGNIy72wM0TZke1VrDOI3ctQGxvAM5ToSe5p/RFEiOgKOfgqxdeT5xpzUZ
iYXVXp1p29P2B1cu+inV1+Dk6gyp2XyTWKS6DeIPYgLgc2pnP+rBCrcyjenHJ+BL
EzLO2iI3NjVFRq6Z329EDdqmgAWMN41MelXofvlSI+QdCKb60YWYxCHuCt2NI9jC
0N6XSrHYSkf1GcsJL48kiRtX1QV25DRRbqNuGgzNciHzChz59k+XLozPKYz/o18L
oTU2MkVh4uTImnGIo5pSLa/pJIDDdkaGW+9T2TCp9+k4sDoi8ctPgJDg842A3DSM
oQtlmEW/LBGrrqGReRB5Dw9jEA5pAH2cwTm7NOtGWW00u7WcacUKhSPMTUfxiW2A
4BAV4Hmbb3O8cTHM0nLVMC4VggltByp4b0Y6R785V8T8eIthB9p1cacPcZp/0u6f
nGeS/tmfaWO29FSskGO79r1EIEtOacM7mXN0vFroykgjXnpIcel6C0AffdpyzGaW
MOJc8HodyTDcc1L05skG7KoqzLnwP2m7Or/dXrmruX+dCw1sFcrS0NQ+j/sU9zEk
swx7uwpsQP4vidbA5uXoR+/qiuZIYW3vKAD+Q1LwPcEJP+WC3KYHFVGzjTOlo4ZH
Ofv8R/PcsYhP+qnaa4rPxGp1m4mk0eZCk7Atzs2aA1QbASYf5jiiB8uHbLHsrKqh
atj7g+dlrW8YUYqIXJpESWUkDozu1PEQDm31NJzF6eMrEIoeZLL84HmRu8M7QDec
/laGFRJlgc1KOZ7SMDNodk/z4AVBsRDFS7P+q9pNHfth9WI82vVLFZoYkHPtZE+W
aDZugoTMZ7JjCAidGKSJZoIaaTVutxS3ipGLOpjLpUzdxKFLtsR8pjQwN09xQcIC
qfpG2mkiw2b/K01OAUHBpTlEXRGHgibHPx3yw+bG1b3A36wrYsfm99Q+M4RDA2Q0
4Kgi6wgoew007pCN675KUYaw67MzjO0mv6L1kAx7AoPGMSjHrRyV0EUWJFCFOjDW
KdYCGjuOn3XQRaSqknJQMkE9j+ro9oJvVsSU40V9XQ4lImXk1mINu9037rBvDX43
cEibvYmoq/Pwb1WRZAxsLYsTlzeHpp/MehxIRsmkhvyR6/Bm9mPF/BJbpoeNxh6m
MhTKwKlSgiLWOHS3mYyXJGTqFdpx7tWxE51TRTtMsYJ6Gw10K3ADm7Y92jgpaux+
O8jGk2kuWT2kj6kO/rSUMKT9BEjTcuPD41lKwMLCJL5NNZFTTY6K7U1Z+idOyV7U
oX5A57dVsEAzRUmAhBFWLL8ajiqEfkGuMlswGDWpVNoRinuxmBiElOqlB9t4TWe5
ACEvDni0ZiK6JaqLfquUvH7vBJuPdB8g7Y59XYAGs2ads0I558nT8B7jb6up0/tH
v93cSko1BGBdxBQomjKBtPMz3vKRsBbdZgAIA08xnfABhNN7bfiMlnHB+kBpw4YL
ixIv8rRwkjdzIuZDGxEsHVwRhWDCLzHYhQbdg1QYlZliMlTnG4FhIMdNq0GUJytj
nZllR+2xpFUkTQ7USW3Y0s4Yx/Z4u/e3Ef38ggc7mgeUXGdS22/CC7MQfq/dr/Ja
fmVWAohZIxVOh12iPqduFzPthXQWs9yHTRglv3g/6523rKlIPAvjD6F1eKmvo5GF
M4ySoprE4u6PRFyc8N/AP8sJIv4azG71QCazGsUV4ZwCc/aj9HvNz1y7+tujjyhS
uvg64tO2EuatWbTokLhVFLxO7T+K8VhqQxmF6p6dGKfRo4R2ImhPApbGw1OnICro
sU1F8rT//r69ae/+xmU9w1OTj055nvi8+0jzsc41qxXX7CEjwZ9cMr0F70X7Qr7h
ZryqzGiq+9dgY+sRQ3FR4WPKzOa7Sb8Op2QVWjeO2qPxQDQC+s3HrP+1YxKxR5hx
GBKF46YxndUb5OEPATKP6yuUFahKVHmobYcIB/cbO7EfPzFNjki4EUE4nhyldQDr
XaYPgebfsava3sVinN494UxDld8GSs/saB/wdBAe0NoSe7dbHa1tEZjQubt+MWqu
2QDGCECMwUmqxDUQfQoQsJjwe6OQGYca2MDSGvMR9sj1TdUWdYKQoI36p107hISs
BJ8ATMP83RmrZLWx7G2wyPhAS2j9n21TqhclGyGoDLn/Q4bCC+rch6X/WhhvVDYQ
fz4XS394yCvZbhUf2khRLfjCFAQdAmOpxRiks0AWxgy/n3bP3upiIjbIVUteJWHg
YdmDh8kISJr03OBBgwQWgwOsCw6qCi8oSHqiWCT0NZZJv7KQK604LgBklewHmgmD
PYoQK2u3eUg7n4W4JlPmHKzctqKIvy5gkiFzOGEBaDMvDiZr7ODxf3he2kViMPXn
aBd1VtxeB+GrYdVZ3ATe1YhtKxTkLK035/LGVhYRWRuCSgIsGof2ROiyqvQdVVUC
0hPDNKXGh9N2laQebpLQUt1w2CnEv4mK0WzyEsg4snpeEDTQxm5UKLbUvrBr9dD1
+qHjlb6MLoU+Of/7wR/qvDQ7loiDkJ6CUK/hfwyQ2s8AEfYOa4ySaYGUCesbu+oH
Nl9VraiTwuO1apl9orGkOZRCmWWO16/CKsIPZk1BLVT4uUG4FrFXi+7GET10EwMF
7ofm+Ryv7Kzm3WEVMzEaP9vbFv36rVnpTlfppjYeJoTBW8BPIxUbzpy5Roce3Qy5
eM8NgjNRjOWwYIlOpBTJam5yt6WzX1kfrFWq/r6SoQylp3d7SNwg9Jq5oVQqkVtl
v57rtL8WLR5vPvrDQxcZzkSWQ/UyuoL/lN/wLX7s48V/tAZKPujf6mRr+p4HSZcR
74zR8NEJSWs5fBYPlnGlhdG6v+zvx0p8atLaw8kaq7eJIRxSSxdCBTqApjOjEjxE
kM/8nfWPp5WbNdv8jZUtwc8skp8dDAvD73BzI6C1TP5gSqmy7d46+PmT+jkTV4Df
tLPF6ry7qdfvOIxxxzH9/OgfRbqLx3Xt8LW0pw3MUzRU9nMhkwsKXTQ/bhl1pm6O
RpQcCoy2lKc5e7JU3VLlRRrUdm/U1tkRvkb+CknIzUsG7Z7EvgXqnzHwY8b0bqcL
99Pvkiq19+JFb/O5JYCXJrIwkARZsI+knSN90NjgMst4sZS5BVnqZerst+DoiqMR
8JyEtT69if5QeZBYXe0Q+sILel/tfaT2o7Jo9M+aZDl4NjUGvey2n2t9PdLxmTzQ
xj1/L4ZwJ1xOttrXWvOw1cc2LNyYHGeLkOdb5LGSUqKpEc1xINWcT60TnSJtDpko
q0EuFsEKrKhZWqqNaaxGFx1+cl9hwRnNwLk4oNBOTA6spkvAZeN9Tl9b9+lsEyQM
QF+6TwP517WxC5e7d0MWjBqdwej6QoEPm/eNPUoAVNb+qCw9wRrbWB7t+jIf1InC
7X9q9tp0e+IzEGZNDLZUS71pamkJRPc2EdXtJMWEY/DpcYHH8xEcs2G3z18dulaR
cZAJY8E3rOKRa1CLyjQR0z4K95PtUBGhqJan4UV6IxkFCJ5/L0smj3daIHCawTFM
25KwykLMOyHik2LnXYJQ90RnFfNJUcGGa1ylHJiOfieE07XwSpBWcxM6iVgEZy/m
om9GLxokEoAI82Vcab8tWhuHwUyksrODPJ+t9jfZDhufIAemmKTt7yDT/NZGcbK4
QlyY1Weg14o7eoRP8AEhYeFNgRZcaiPHYkWWDsLLJmvBBmDR2DCMZppxEbJWRdBf
DZawOvkijZvH9EcZFz3Lcwnk1qkXSn4MR/gxwPfAnkPL6uaA+otPAsgqk4tm9aRu
jL9JDD4uzJss4bNUApI52aBS4/10aLs4kxiZhcK08OeLqvhrm2OQEq/1zX5l8PVT
POMCYvNkmLC+7HyKqPDYNNMcJe5AtnkgiraeY2xThlqMXpesjfGVF9UFk2Lda4Ni
3zdfDyDCXLdVQBh72Um2RamCA3QBd9iwqHcaDBMM15B5/tio5pwFHuCpnM3+9ZLk
rV0dHw4j6L/wpCFac+25Y3IPmIKYmeRFlLueedio6ycCnnUWPKdP4K5AEPevQzTk
/P7qHQYycOXq8FsV4HWsvTpp4ylKiTkOSWuMc+4mC4PuOiC21VSZXGfl+WEpF0P7
zFcT3g1Fz4Ng9w6wz/uytpIzmlcngwztq8QCuRVLK3oloYcgQxFCZztqc78Go6wS
feUel/TR1xcue8slF6wbA1YdSeGmBmTBwyk2RfJC//dPCLk7HECYjBwiPgIgpdsP
Az77lW5EDd6gF2OPVb3wf2ZgmWvBvmYGAeb+CoMLZrQngcvdgaGeMay1/kpW23OU
/fjeEVtR6fmPYVS1k0oHdSx7Qah/vGZqJqtxSvfHetJGoid73tyn0jL1AAHXH9s2
scOItgOWjsry4o57JTkZExL2SCEOTlndc+WbBMVn+PjUJW2KGdwrpc4oH3RFv1Uj
o4cO7l3zgOoNlzxLTy//4BvzyODkBrFYewxHB1OLS5RaMvmcnsAOZzGD72naH2kq
OoROy4a7YpYBydutJ3NR4dgXUksZD2dFFhzDHlyI8FGCuv0qwpOC5JyGj+3eVVC5
AbPisg0WzjjWdDirtuYV3Uef0gOdAbIuscD3lzKN+lOoSJxvdm7K+O8z1+z6cptY
YyrUvDN0BM5MFx86MU5Qj6AGrlRFOOwv6q5rX9tDVFoGpnc2QGd4TMbkMMlTBwHM
kb4YfVpYcf9OULOybG5/NcL19YehGG9FwNmMGvWSY0duOVP5+GGJJRqKZ4eLuw9B
RXd7OzigUtQp6XnhH3NgyJojgJAyf7qyoZl6PuP01Tspx40Wnc8zjJ8qkYFDX0mi
EIhz2yzHj7rbgqrrzeImvIlCcp6fCOORqdOSYcSN2gHQ/e/wow57Cbm9th4cci17
sUI20KkkMB+IBFtSNLWZRWY3yp9WBpMhv/9DO/WxKmPRa4a2rpFEakJHSe0fTVch
9gyWDLQ0NpZ4k/f8nN+ffwfSSo8OE3QYUhFa9m+Gj/jsgiiiZjiajVzOtOeVBvkQ
RWK1EkHNSF/IfUnHOdJZso09o35rh3UEeGUNa9kcwH2KHiPjE7cR5G1m1C97bBHf
F4zT94+C+wpWs9peGsClMqvHI/no4a1CruudYOqt3cjqDwqeCETZ8pjy94W4ndvX
GhmUvcU/dlkd2dyRjz5Wah17sEy1sx+cyHVs72St8oitXPRAw719mlTNyYL1U7mP
JukYDhWZl63000XHylJSmpC79/1NsE+i4gi/PpbTtzUvceZ0EhrRMOyVz6wsD8DZ
0yEFC5TSOzhFQ5708WioVTq4ue+LyI9K941wudGOJqcJHo2MpCSRJ6oVEI8uRX56
onCO72i5ASI4R8nm9XkMhvUQ6/HKAJw+h7/AMEaGshi/m3cmwaALPNum9FA7l3vA
MsyuPDH2RmHePPmeZi+0PH/3J2bnL7cZwaGQmopH1iDgRRScpIUFpkpeOkmT6uQN
cBew9iXTVun49Mnqi7fGEDtly6nJC8ZtyCFgs7iQrBxzALb/skvXjmvmtw2lrJit
fKKQ/g0nHfomyU/mAwAgqFwkh6crb6Tu3RgItL+BrONbz6PQYWVyR4LQKXPkjpYM
gnXY5IQS00DqeMmtL4DpOG05I0LSKhAJs+OPb/ZCItWsS2sxFf6LtJgvSl9xJNo7
AmhiVUkjKKXZq09/9UWkd/xyY7uQbJ7WqImA7ss9qtqvN7vXkyZxKdBF9gB1T+CU
UEd7X0BlnkdL+gDW8l7mP4T/v2i08+Wd3qOezeYoLVYEj67DmljXo793HN4VdVvl
rm0dewp4KKGgPf5f7KiQNGgHNQmxKTf7qG3O2oXp7OFipiJgiwOtWtHiS/pHhPEm
Ys1szWIOMkhoNafUkS7vpQ==
`pragma protect end_protected
