��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`w�z�5��#C�iL-G����=:�������~ʵi����]�n�xz��શ)���'�z�C]�w��{��|&('D���U���D�D�R�C�5)[{&�hUS5̹�W9�9�y�u�m��~3@^z���ɧ�{�@�RB byo��< ��{��$�
ѯ�$�%����?�}
�wɣhz����p���Lߜ�c�.3������p!��N�������u���3��p��e��X���Y3+�v	����a�,��[�k���7�:�o�^��vq��HoqҶ�Y�,S?�)�7�0�G�~S�
�rFϳ<�%Y�_���u6�l��h�� l�"FP4�6�֏�����p*�x�$��u�U1ub<���O���瘬G��$l��8�Ϟ]�N�=QC�����ɓ�AyD�cC��-�q��򱞓7�䶡�Z�s6���=\�{˱�F�R�e�P��F~Z-\��Q���Á�>�XGɽ�����q�ïl�?%u��6+˅^���f��f>���
���J���/&�(�Ş�J�֊��Pia`�C�V��o��t%@jV��k1�R��?����p#��o��K�OA�����W" ������
��	�.�l%��8��P��j5�{�{[�f/�D/��/�9�<]��.�hr�����h".p���|w���������R�=٫G�et#�R�� x��\E����8|DN!��V,�Gٜ�f�P[ǯ1�P,�_��h/q�C��t��o��F��QYT�B:�4p!�3�<�fz����p�u�>w�����lr,�h�H}Al��1�Ţ���C�� t5���u�r�X�oӧ�I�PG˂Bj��0�T�6�|���r�x��L�q���=�_դ�1(�0WRy���J���3#�[O��w�(��i�AX,��Ⱦ���Д48�ղYY��1ck�6�U��\D˯c�[r�Q�R���Vu��5�ԩ/�T��Q�_}�Z��[�9�)�:�x���2��C��:O�p����|K���L�`�%tY0��'GI�J�s����`��F�������'
g.�Y����\4A�e��Z3<�᷀�%F�T����ȴH*�A�;�5�Lp"0kI>�f��[������>ݭ&�V 4EºcCS�pс��.:#�����1�RS�s�JGh�
A�M�ĉ��3uC�nG;Kٟp[�XSҠ�I�1�L���F��������:��ׂ���j�1��?˂���%�-���r�&[�G��/%�x������o��ِ���+v�l^�Yoi�e���MW�|�4�2��[�פ����ҫa����%�<�i�g�+�j����E� @�R�Xˣ�����i���ز��0$�j����?\�}�9��朗?�X�j�r��p��Y?���;'je�kv�I^ԿR�� �U��h#�Q�eBxH 00�^%�Nc���3TYt�g�~"�0�śܣ>��^	�V� 
n�����׆��L�4���n�1t��s5w?��ȨL�-{���,;u�vO?_