//------------------------------------------------------------
// Project: HYBRID_CONTROL
// Author: Nicola Zaupa
// Date: (2022/02/23) (10:20:49)
// File: trigonometry_deg.v
//------------------------------------------------------------
// Description:
//
// Compuation of sine and cosine of an angle [-180,360]
// angle  x 1
// output x 1000
//------------------------------------------------------------


`timescale 1 ns / 1 ps
//`default_nettype none


module trigonometry_deg (
   o_cos,    // cosine of the input
   o_sin,    // sine of the input
   i_theta   // input angle
);

output [31:0] o_sin;
output [31:0] o_cos;
input  [31:0] i_theta;

// output  signed [31:0] o_sin;
// output  signed [31:0] o_cos;
// input   signed [31:0] i_theta;

// wire [31:0] o_sin;
// wire [31:0] o_cos;
// wire [31:0] i_theta;

reg [31:0] r_sin;
reg [31:0] r_cos;

assign o_sin = r_sin;
assign o_cos = r_cos;


always @ ( i_theta )
begin

// computation of sine and cosine using integers
// taking advanatges of look-up-table
// input angle is multiplied by x100
// trigonometric output is multiplied by x1000

case(i_theta)
      32'hFFFFFF4C: r_sin = 32'h00000000;
      32'hFFFFFF4D: r_sin = 32'hFFFFFFEF;
      32'hFFFFFF4E: r_sin = 32'hFFFFFFDD;
      32'hFFFFFF4F: r_sin = 32'hFFFFFFCC;
      32'hFFFFFF50: r_sin = 32'hFFFFFFBA;
      32'hFFFFFF51: r_sin = 32'hFFFFFFA9;
      32'hFFFFFF52: r_sin = 32'hFFFFFF97;
      32'hFFFFFF53: r_sin = 32'hFFFFFF86;
      32'hFFFFFF54: r_sin = 32'hFFFFFF75;
      32'hFFFFFF55: r_sin = 32'hFFFFFF64;
      32'hFFFFFF56: r_sin = 32'hFFFFFF52;
      32'hFFFFFF57: r_sin = 32'hFFFFFF41;
      32'hFFFFFF58: r_sin = 32'hFFFFFF30;
      32'hFFFFFF59: r_sin = 32'hFFFFFF1F;
      32'hFFFFFF5A: r_sin = 32'hFFFFFF0E;
      32'hFFFFFF5B: r_sin = 32'hFFFFFEFD;
      32'hFFFFFF5C: r_sin = 32'hFFFFFEEC;
      32'hFFFFFF5D: r_sin = 32'hFFFFFEDC;
      32'hFFFFFF5E: r_sin = 32'hFFFFFECB;
      32'hFFFFFF5F: r_sin = 32'hFFFFFEBA;
      32'hFFFFFF60: r_sin = 32'hFFFFFEAA;
      32'hFFFFFF61: r_sin = 32'hFFFFFE9A;
      32'hFFFFFF62: r_sin = 32'hFFFFFE89;
      32'hFFFFFF63: r_sin = 32'hFFFFFE79;
      32'hFFFFFF64: r_sin = 32'hFFFFFE69;
      32'hFFFFFF65: r_sin = 32'hFFFFFE59;
      32'hFFFFFF66: r_sin = 32'hFFFFFE4A;
      32'hFFFFFF67: r_sin = 32'hFFFFFE3A;
      32'hFFFFFF68: r_sin = 32'hFFFFFE2B;
      32'hFFFFFF69: r_sin = 32'hFFFFFE1B;
      32'hFFFFFF6A: r_sin = 32'hFFFFFE0C;
      32'hFFFFFF6B: r_sin = 32'hFFFFFDFD;
      32'hFFFFFF6C: r_sin = 32'hFFFFFDEE;
      32'hFFFFFF6D: r_sin = 32'hFFFFFDDF;
      32'hFFFFFF6E: r_sin = 32'hFFFFFDD1;
      32'hFFFFFF6F: r_sin = 32'hFFFFFDC2;
      32'hFFFFFF70: r_sin = 32'hFFFFFDB4;
      32'hFFFFFF71: r_sin = 32'hFFFFFDA6;
      32'hFFFFFF72: r_sin = 32'hFFFFFD98;
      32'hFFFFFF73: r_sin = 32'hFFFFFD8B;
      32'hFFFFFF74: r_sin = 32'hFFFFFD7D;
      32'hFFFFFF75: r_sin = 32'hFFFFFD70;
      32'hFFFFFF76: r_sin = 32'hFFFFFD63;
      32'hFFFFFF77: r_sin = 32'hFFFFFD56;
      32'hFFFFFF78: r_sin = 32'hFFFFFD49;
      32'hFFFFFF79: r_sin = 32'hFFFFFD3D;
      32'hFFFFFF7A: r_sin = 32'hFFFFFD31;
      32'hFFFFFF7B: r_sin = 32'hFFFFFD25;
      32'hFFFFFF7C: r_sin = 32'hFFFFFD19;
      32'hFFFFFF7D: r_sin = 32'hFFFFFD0D;
      32'hFFFFFF7E: r_sin = 32'hFFFFFD02;
      32'hFFFFFF7F: r_sin = 32'hFFFFFCF7;
      32'hFFFFFF80: r_sin = 32'hFFFFFCEC;
      32'hFFFFFF81: r_sin = 32'hFFFFFCE1;
      32'hFFFFFF82: r_sin = 32'hFFFFFCD7;
      32'hFFFFFF83: r_sin = 32'hFFFFFCCD;
      32'hFFFFFF84: r_sin = 32'hFFFFFCC3;
      32'hFFFFFF85: r_sin = 32'hFFFFFCB9;
      32'hFFFFFF86: r_sin = 32'hFFFFFCB0;
      32'hFFFFFF87: r_sin = 32'hFFFFFCA7;
      32'hFFFFFF88: r_sin = 32'hFFFFFC9E;
      32'hFFFFFF89: r_sin = 32'hFFFFFC95;
      32'hFFFFFF8A: r_sin = 32'hFFFFFC8D;
      32'hFFFFFF8B: r_sin = 32'hFFFFFC85;
      32'hFFFFFF8C: r_sin = 32'hFFFFFC7D;
      32'hFFFFFF8D: r_sin = 32'hFFFFFC76;
      32'hFFFFFF8E: r_sin = 32'hFFFFFC6E;
      32'hFFFFFF8F: r_sin = 32'hFFFFFC67;
      32'hFFFFFF90: r_sin = 32'hFFFFFC61;
      32'hFFFFFF91: r_sin = 32'hFFFFFC5A;
      32'hFFFFFF92: r_sin = 32'hFFFFFC54;
      32'hFFFFFF93: r_sin = 32'hFFFFFC4E;
      32'hFFFFFF94: r_sin = 32'hFFFFFC49;
      32'hFFFFFF95: r_sin = 32'hFFFFFC44;
      32'hFFFFFF96: r_sin = 32'hFFFFFC3F;
      32'hFFFFFF97: r_sin = 32'hFFFFFC3A;
      32'hFFFFFF98: r_sin = 32'hFFFFFC36;
      32'hFFFFFF99: r_sin = 32'hFFFFFC32;
      32'hFFFFFF9A: r_sin = 32'hFFFFFC2E;
      32'hFFFFFF9B: r_sin = 32'hFFFFFC2A;
      32'hFFFFFF9C: r_sin = 32'hFFFFFC27;
      32'hFFFFFF9D: r_sin = 32'hFFFFFC24;
      32'hFFFFFF9E: r_sin = 32'hFFFFFC22;
      32'hFFFFFF9F: r_sin = 32'hFFFFFC1F;
      32'hFFFFFFA0: r_sin = 32'hFFFFFC1D;
      32'hFFFFFFA1: r_sin = 32'hFFFFFC1C;
      32'hFFFFFFA2: r_sin = 32'hFFFFFC1A;
      32'hFFFFFFA3: r_sin = 32'hFFFFFC19;
      32'hFFFFFFA4: r_sin = 32'hFFFFFC19;
      32'hFFFFFFA5: r_sin = 32'hFFFFFC18;
      32'hFFFFFFA6: r_sin = 32'hFFFFFC18;
      32'hFFFFFFA7: r_sin = 32'hFFFFFC18;
      32'hFFFFFFA8: r_sin = 32'hFFFFFC19;
      32'hFFFFFFA9: r_sin = 32'hFFFFFC19;
      32'hFFFFFFAA: r_sin = 32'hFFFFFC1A;
      32'hFFFFFFAB: r_sin = 32'hFFFFFC1C;
      32'hFFFFFFAC: r_sin = 32'hFFFFFC1D;
      32'hFFFFFFAD: r_sin = 32'hFFFFFC1F;
      32'hFFFFFFAE: r_sin = 32'hFFFFFC22;
      32'hFFFFFFAF: r_sin = 32'hFFFFFC24;
      32'hFFFFFFB0: r_sin = 32'hFFFFFC27;
      32'hFFFFFFB1: r_sin = 32'hFFFFFC2A;
      32'hFFFFFFB2: r_sin = 32'hFFFFFC2E;
      32'hFFFFFFB3: r_sin = 32'hFFFFFC32;
      32'hFFFFFFB4: r_sin = 32'hFFFFFC36;
      32'hFFFFFFB5: r_sin = 32'hFFFFFC3A;
      32'hFFFFFFB6: r_sin = 32'hFFFFFC3F;
      32'hFFFFFFB7: r_sin = 32'hFFFFFC44;
      32'hFFFFFFB8: r_sin = 32'hFFFFFC49;
      32'hFFFFFFB9: r_sin = 32'hFFFFFC4E;
      32'hFFFFFFBA: r_sin = 32'hFFFFFC54;
      32'hFFFFFFBB: r_sin = 32'hFFFFFC5A;
      32'hFFFFFFBC: r_sin = 32'hFFFFFC61;
      32'hFFFFFFBD: r_sin = 32'hFFFFFC67;
      32'hFFFFFFBE: r_sin = 32'hFFFFFC6E;
      32'hFFFFFFBF: r_sin = 32'hFFFFFC76;
      32'hFFFFFFC0: r_sin = 32'hFFFFFC7D;
      32'hFFFFFFC1: r_sin = 32'hFFFFFC85;
      32'hFFFFFFC2: r_sin = 32'hFFFFFC8D;
      32'hFFFFFFC3: r_sin = 32'hFFFFFC95;
      32'hFFFFFFC4: r_sin = 32'hFFFFFC9E;
      32'hFFFFFFC5: r_sin = 32'hFFFFFCA7;
      32'hFFFFFFC6: r_sin = 32'hFFFFFCB0;
      32'hFFFFFFC7: r_sin = 32'hFFFFFCB9;
      32'hFFFFFFC8: r_sin = 32'hFFFFFCC3;
      32'hFFFFFFC9: r_sin = 32'hFFFFFCCD;
      32'hFFFFFFCA: r_sin = 32'hFFFFFCD7;
      32'hFFFFFFCB: r_sin = 32'hFFFFFCE1;
      32'hFFFFFFCC: r_sin = 32'hFFFFFCEC;
      32'hFFFFFFCD: r_sin = 32'hFFFFFCF7;
      32'hFFFFFFCE: r_sin = 32'hFFFFFD02;
      32'hFFFFFFCF: r_sin = 32'hFFFFFD0D;
      32'hFFFFFFD0: r_sin = 32'hFFFFFD19;
      32'hFFFFFFD1: r_sin = 32'hFFFFFD25;
      32'hFFFFFFD2: r_sin = 32'hFFFFFD31;
      32'hFFFFFFD3: r_sin = 32'hFFFFFD3D;
      32'hFFFFFFD4: r_sin = 32'hFFFFFD49;
      32'hFFFFFFD5: r_sin = 32'hFFFFFD56;
      32'hFFFFFFD6: r_sin = 32'hFFFFFD63;
      32'hFFFFFFD7: r_sin = 32'hFFFFFD70;
      32'hFFFFFFD8: r_sin = 32'hFFFFFD7D;
      32'hFFFFFFD9: r_sin = 32'hFFFFFD8B;
      32'hFFFFFFDA: r_sin = 32'hFFFFFD98;
      32'hFFFFFFDB: r_sin = 32'hFFFFFDA6;
      32'hFFFFFFDC: r_sin = 32'hFFFFFDB4;
      32'hFFFFFFDD: r_sin = 32'hFFFFFDC2;
      32'hFFFFFFDE: r_sin = 32'hFFFFFDD1;
      32'hFFFFFFDF: r_sin = 32'hFFFFFDDF;
      32'hFFFFFFE0: r_sin = 32'hFFFFFDEE;
      32'hFFFFFFE1: r_sin = 32'hFFFFFDFD;
      32'hFFFFFFE2: r_sin = 32'hFFFFFE0C;
      32'hFFFFFFE3: r_sin = 32'hFFFFFE1B;
      32'hFFFFFFE4: r_sin = 32'hFFFFFE2B;
      32'hFFFFFFE5: r_sin = 32'hFFFFFE3A;
      32'hFFFFFFE6: r_sin = 32'hFFFFFE4A;
      32'hFFFFFFE7: r_sin = 32'hFFFFFE59;
      32'hFFFFFFE8: r_sin = 32'hFFFFFE69;
      32'hFFFFFFE9: r_sin = 32'hFFFFFE79;
      32'hFFFFFFEA: r_sin = 32'hFFFFFE89;
      32'hFFFFFFEB: r_sin = 32'hFFFFFE9A;
      32'hFFFFFFEC: r_sin = 32'hFFFFFEAA;
      32'hFFFFFFED: r_sin = 32'hFFFFFEBA;
      32'hFFFFFFEE: r_sin = 32'hFFFFFECB;
      32'hFFFFFFEF: r_sin = 32'hFFFFFEDC;
      32'hFFFFFFF0: r_sin = 32'hFFFFFEEC;
      32'hFFFFFFF1: r_sin = 32'hFFFFFEFD;
      32'hFFFFFFF2: r_sin = 32'hFFFFFF0E;
      32'hFFFFFFF3: r_sin = 32'hFFFFFF1F;
      32'hFFFFFFF4: r_sin = 32'hFFFFFF30;
      32'hFFFFFFF5: r_sin = 32'hFFFFFF41;
      32'hFFFFFFF6: r_sin = 32'hFFFFFF52;
      32'hFFFFFFF7: r_sin = 32'hFFFFFF64;
      32'hFFFFFFF8: r_sin = 32'hFFFFFF75;
      32'hFFFFFFF9: r_sin = 32'hFFFFFF86;
      32'hFFFFFFFA: r_sin = 32'hFFFFFF97;
      32'hFFFFFFFB: r_sin = 32'hFFFFFFA9;
      32'hFFFFFFFC: r_sin = 32'hFFFFFFBA;
      32'hFFFFFFFD: r_sin = 32'hFFFFFFCC;
      32'hFFFFFFFE: r_sin = 32'hFFFFFFDD;
      32'hFFFFFFFF: r_sin = 32'hFFFFFFEF;
      32'h00000000: r_sin = 32'h00000000;
      32'h00000001: r_sin = 32'h00000011;
      32'h00000002: r_sin = 32'h00000023;
      32'h00000003: r_sin = 32'h00000034;
      32'h00000004: r_sin = 32'h00000046;
      32'h00000005: r_sin = 32'h00000057;
      32'h00000006: r_sin = 32'h00000069;
      32'h00000007: r_sin = 32'h0000007A;
      32'h00000008: r_sin = 32'h0000008B;
      32'h00000009: r_sin = 32'h0000009C;
      32'h0000000A: r_sin = 32'h000000AE;
      32'h0000000B: r_sin = 32'h000000BF;
      32'h0000000C: r_sin = 32'h000000D0;
      32'h0000000D: r_sin = 32'h000000E1;
      32'h0000000E: r_sin = 32'h000000F2;
      32'h0000000F: r_sin = 32'h00000103;
      32'h00000010: r_sin = 32'h00000114;
      32'h00000011: r_sin = 32'h00000124;
      32'h00000012: r_sin = 32'h00000135;
      32'h00000013: r_sin = 32'h00000146;
      32'h00000014: r_sin = 32'h00000156;
      32'h00000015: r_sin = 32'h00000166;
      32'h00000016: r_sin = 32'h00000177;
      32'h00000017: r_sin = 32'h00000187;
      32'h00000018: r_sin = 32'h00000197;
      32'h00000019: r_sin = 32'h000001A7;
      32'h0000001A: r_sin = 32'h000001B6;
      32'h0000001B: r_sin = 32'h000001C6;
      32'h0000001C: r_sin = 32'h000001D5;
      32'h0000001D: r_sin = 32'h000001E5;
      32'h0000001E: r_sin = 32'h000001F4;
      32'h0000001F: r_sin = 32'h00000203;
      32'h00000020: r_sin = 32'h00000212;
      32'h00000021: r_sin = 32'h00000221;
      32'h00000022: r_sin = 32'h0000022F;
      32'h00000023: r_sin = 32'h0000023E;
      32'h00000024: r_sin = 32'h0000024C;
      32'h00000025: r_sin = 32'h0000025A;
      32'h00000026: r_sin = 32'h00000268;
      32'h00000027: r_sin = 32'h00000275;
      32'h00000028: r_sin = 32'h00000283;
      32'h00000029: r_sin = 32'h00000290;
      32'h0000002A: r_sin = 32'h0000029D;
      32'h0000002B: r_sin = 32'h000002AA;
      32'h0000002C: r_sin = 32'h000002B7;
      32'h0000002D: r_sin = 32'h000002C3;
      32'h0000002E: r_sin = 32'h000002CF;
      32'h0000002F: r_sin = 32'h000002DB;
      32'h00000030: r_sin = 32'h000002E7;
      32'h00000031: r_sin = 32'h000002F3;
      32'h00000032: r_sin = 32'h000002FE;
      32'h00000033: r_sin = 32'h00000309;
      32'h00000034: r_sin = 32'h00000314;
      32'h00000035: r_sin = 32'h0000031F;
      32'h00000036: r_sin = 32'h00000329;
      32'h00000037: r_sin = 32'h00000333;
      32'h00000038: r_sin = 32'h0000033D;
      32'h00000039: r_sin = 32'h00000347;
      32'h0000003A: r_sin = 32'h00000350;
      32'h0000003B: r_sin = 32'h00000359;
      32'h0000003C: r_sin = 32'h00000362;
      32'h0000003D: r_sin = 32'h0000036B;
      32'h0000003E: r_sin = 32'h00000373;
      32'h0000003F: r_sin = 32'h0000037B;
      32'h00000040: r_sin = 32'h00000383;
      32'h00000041: r_sin = 32'h0000038A;
      32'h00000042: r_sin = 32'h00000392;
      32'h00000043: r_sin = 32'h00000399;
      32'h00000044: r_sin = 32'h0000039F;
      32'h00000045: r_sin = 32'h000003A6;
      32'h00000046: r_sin = 32'h000003AC;
      32'h00000047: r_sin = 32'h000003B2;
      32'h00000048: r_sin = 32'h000003B7;
      32'h00000049: r_sin = 32'h000003BC;
      32'h0000004A: r_sin = 32'h000003C1;
      32'h0000004B: r_sin = 32'h000003C6;
      32'h0000004C: r_sin = 32'h000003CA;
      32'h0000004D: r_sin = 32'h000003CE;
      32'h0000004E: r_sin = 32'h000003D2;
      32'h0000004F: r_sin = 32'h000003D6;
      32'h00000050: r_sin = 32'h000003D9;
      32'h00000051: r_sin = 32'h000003DC;
      32'h00000052: r_sin = 32'h000003DE;
      32'h00000053: r_sin = 32'h000003E1;
      32'h00000054: r_sin = 32'h000003E3;
      32'h00000055: r_sin = 32'h000003E4;
      32'h00000056: r_sin = 32'h000003E6;
      32'h00000057: r_sin = 32'h000003E7;
      32'h00000058: r_sin = 32'h000003E7;
      32'h00000059: r_sin = 32'h000003E8;
      32'h0000005A: r_sin = 32'h000003E8;
      32'h0000005B: r_sin = 32'h000003E8;
      32'h0000005C: r_sin = 32'h000003E7;
      32'h0000005D: r_sin = 32'h000003E7;
      32'h0000005E: r_sin = 32'h000003E6;
      32'h0000005F: r_sin = 32'h000003E4;
      32'h00000060: r_sin = 32'h000003E3;
      32'h00000061: r_sin = 32'h000003E1;
      32'h00000062: r_sin = 32'h000003DE;
      32'h00000063: r_sin = 32'h000003DC;
      32'h00000064: r_sin = 32'h000003D9;
      32'h00000065: r_sin = 32'h000003D6;
      32'h00000066: r_sin = 32'h000003D2;
      32'h00000067: r_sin = 32'h000003CE;
      32'h00000068: r_sin = 32'h000003CA;
      32'h00000069: r_sin = 32'h000003C6;
      32'h0000006A: r_sin = 32'h000003C1;
      32'h0000006B: r_sin = 32'h000003BC;
      32'h0000006C: r_sin = 32'h000003B7;
      32'h0000006D: r_sin = 32'h000003B2;
      32'h0000006E: r_sin = 32'h000003AC;
      32'h0000006F: r_sin = 32'h000003A6;
      32'h00000070: r_sin = 32'h0000039F;
      32'h00000071: r_sin = 32'h00000399;
      32'h00000072: r_sin = 32'h00000392;
      32'h00000073: r_sin = 32'h0000038A;
      32'h00000074: r_sin = 32'h00000383;
      32'h00000075: r_sin = 32'h0000037B;
      32'h00000076: r_sin = 32'h00000373;
      32'h00000077: r_sin = 32'h0000036B;
      32'h00000078: r_sin = 32'h00000362;
      32'h00000079: r_sin = 32'h00000359;
      32'h0000007A: r_sin = 32'h00000350;
      32'h0000007B: r_sin = 32'h00000347;
      32'h0000007C: r_sin = 32'h0000033D;
      32'h0000007D: r_sin = 32'h00000333;
      32'h0000007E: r_sin = 32'h00000329;
      32'h0000007F: r_sin = 32'h0000031F;
      32'h00000080: r_sin = 32'h00000314;
      32'h00000081: r_sin = 32'h00000309;
      32'h00000082: r_sin = 32'h000002FE;
      32'h00000083: r_sin = 32'h000002F3;
      32'h00000084: r_sin = 32'h000002E7;
      32'h00000085: r_sin = 32'h000002DB;
      32'h00000086: r_sin = 32'h000002CF;
      32'h00000087: r_sin = 32'h000002C3;
      32'h00000088: r_sin = 32'h000002B7;
      32'h00000089: r_sin = 32'h000002AA;
      32'h0000008A: r_sin = 32'h0000029D;
      32'h0000008B: r_sin = 32'h00000290;
      32'h0000008C: r_sin = 32'h00000283;
      32'h0000008D: r_sin = 32'h00000275;
      32'h0000008E: r_sin = 32'h00000268;
      32'h0000008F: r_sin = 32'h0000025A;
      32'h00000090: r_sin = 32'h0000024C;
      32'h00000091: r_sin = 32'h0000023E;
      32'h00000092: r_sin = 32'h0000022F;
      32'h00000093: r_sin = 32'h00000221;
      32'h00000094: r_sin = 32'h00000212;
      32'h00000095: r_sin = 32'h00000203;
      32'h00000096: r_sin = 32'h000001F4;
      32'h00000097: r_sin = 32'h000001E5;
      32'h00000098: r_sin = 32'h000001D5;
      32'h00000099: r_sin = 32'h000001C6;
      32'h0000009A: r_sin = 32'h000001B6;
      32'h0000009B: r_sin = 32'h000001A7;
      32'h0000009C: r_sin = 32'h00000197;
      32'h0000009D: r_sin = 32'h00000187;
      32'h0000009E: r_sin = 32'h00000177;
      32'h0000009F: r_sin = 32'h00000166;
      32'h000000A0: r_sin = 32'h00000156;
      32'h000000A1: r_sin = 32'h00000146;
      32'h000000A2: r_sin = 32'h00000135;
      32'h000000A3: r_sin = 32'h00000124;
      32'h000000A4: r_sin = 32'h00000114;
      32'h000000A5: r_sin = 32'h00000103;
      32'h000000A6: r_sin = 32'h000000F2;
      32'h000000A7: r_sin = 32'h000000E1;
      32'h000000A8: r_sin = 32'h000000D0;
      32'h000000A9: r_sin = 32'h000000BF;
      32'h000000AA: r_sin = 32'h000000AE;
      32'h000000AB: r_sin = 32'h0000009C;
      32'h000000AC: r_sin = 32'h0000008B;
      32'h000000AD: r_sin = 32'h0000007A;
      32'h000000AE: r_sin = 32'h00000069;
      32'h000000AF: r_sin = 32'h00000057;
      32'h000000B0: r_sin = 32'h00000046;
      32'h000000B1: r_sin = 32'h00000034;
      32'h000000B2: r_sin = 32'h00000023;
      32'h000000B3: r_sin = 32'h00000011;
      32'h000000B4: r_sin = 32'h00000000;
      32'h000000B5: r_sin = 32'hFFFFFFEF;
      32'h000000B6: r_sin = 32'hFFFFFFDD;
      32'h000000B7: r_sin = 32'hFFFFFFCC;
      32'h000000B8: r_sin = 32'hFFFFFFBA;
      32'h000000B9: r_sin = 32'hFFFFFFA9;
      32'h000000BA: r_sin = 32'hFFFFFF97;
      32'h000000BB: r_sin = 32'hFFFFFF86;
      32'h000000BC: r_sin = 32'hFFFFFF75;
      32'h000000BD: r_sin = 32'hFFFFFF64;
      32'h000000BE: r_sin = 32'hFFFFFF52;
      32'h000000BF: r_sin = 32'hFFFFFF41;
      32'h000000C0: r_sin = 32'hFFFFFF30;
      32'h000000C1: r_sin = 32'hFFFFFF1F;
      32'h000000C2: r_sin = 32'hFFFFFF0E;
      32'h000000C3: r_sin = 32'hFFFFFEFD;
      32'h000000C4: r_sin = 32'hFFFFFEEC;
      32'h000000C5: r_sin = 32'hFFFFFEDC;
      32'h000000C6: r_sin = 32'hFFFFFECB;
      32'h000000C7: r_sin = 32'hFFFFFEBA;
      32'h000000C8: r_sin = 32'hFFFFFEAA;
      32'h000000C9: r_sin = 32'hFFFFFE9A;
      32'h000000CA: r_sin = 32'hFFFFFE89;
      32'h000000CB: r_sin = 32'hFFFFFE79;
      32'h000000CC: r_sin = 32'hFFFFFE69;
      32'h000000CD: r_sin = 32'hFFFFFE59;
      32'h000000CE: r_sin = 32'hFFFFFE4A;
      32'h000000CF: r_sin = 32'hFFFFFE3A;
      32'h000000D0: r_sin = 32'hFFFFFE2B;
      32'h000000D1: r_sin = 32'hFFFFFE1B;
      32'h000000D2: r_sin = 32'hFFFFFE0C;
      32'h000000D3: r_sin = 32'hFFFFFDFD;
      32'h000000D4: r_sin = 32'hFFFFFDEE;
      32'h000000D5: r_sin = 32'hFFFFFDDF;
      32'h000000D6: r_sin = 32'hFFFFFDD1;
      32'h000000D7: r_sin = 32'hFFFFFDC2;
      32'h000000D8: r_sin = 32'hFFFFFDB4;
      32'h000000D9: r_sin = 32'hFFFFFDA6;
      32'h000000DA: r_sin = 32'hFFFFFD98;
      32'h000000DB: r_sin = 32'hFFFFFD8B;
      32'h000000DC: r_sin = 32'hFFFFFD7D;
      32'h000000DD: r_sin = 32'hFFFFFD70;
      32'h000000DE: r_sin = 32'hFFFFFD63;
      32'h000000DF: r_sin = 32'hFFFFFD56;
      32'h000000E0: r_sin = 32'hFFFFFD49;
      32'h000000E1: r_sin = 32'hFFFFFD3D;
      32'h000000E2: r_sin = 32'hFFFFFD31;
      32'h000000E3: r_sin = 32'hFFFFFD25;
      32'h000000E4: r_sin = 32'hFFFFFD19;
      32'h000000E5: r_sin = 32'hFFFFFD0D;
      32'h000000E6: r_sin = 32'hFFFFFD02;
      32'h000000E7: r_sin = 32'hFFFFFCF7;
      32'h000000E8: r_sin = 32'hFFFFFCEC;
      32'h000000E9: r_sin = 32'hFFFFFCE1;
      32'h000000EA: r_sin = 32'hFFFFFCD7;
      32'h000000EB: r_sin = 32'hFFFFFCCD;
      32'h000000EC: r_sin = 32'hFFFFFCC3;
      32'h000000ED: r_sin = 32'hFFFFFCB9;
      32'h000000EE: r_sin = 32'hFFFFFCB0;
      32'h000000EF: r_sin = 32'hFFFFFCA7;
      32'h000000F0: r_sin = 32'hFFFFFC9E;
      32'h000000F1: r_sin = 32'hFFFFFC95;
      32'h000000F2: r_sin = 32'hFFFFFC8D;
      32'h000000F3: r_sin = 32'hFFFFFC85;
      32'h000000F4: r_sin = 32'hFFFFFC7D;
      32'h000000F5: r_sin = 32'hFFFFFC76;
      32'h000000F6: r_sin = 32'hFFFFFC6E;
      32'h000000F7: r_sin = 32'hFFFFFC67;
      32'h000000F8: r_sin = 32'hFFFFFC61;
      32'h000000F9: r_sin = 32'hFFFFFC5A;
      32'h000000FA: r_sin = 32'hFFFFFC54;
      32'h000000FB: r_sin = 32'hFFFFFC4E;
      32'h000000FC: r_sin = 32'hFFFFFC49;
      32'h000000FD: r_sin = 32'hFFFFFC44;
      32'h000000FE: r_sin = 32'hFFFFFC3F;
      32'h000000FF: r_sin = 32'hFFFFFC3A;
      32'h00000100: r_sin = 32'hFFFFFC36;
      32'h00000101: r_sin = 32'hFFFFFC32;
      32'h00000102: r_sin = 32'hFFFFFC2E;
      32'h00000103: r_sin = 32'hFFFFFC2A;
      32'h00000104: r_sin = 32'hFFFFFC27;
      32'h00000105: r_sin = 32'hFFFFFC24;
      32'h00000106: r_sin = 32'hFFFFFC22;
      32'h00000107: r_sin = 32'hFFFFFC1F;
      32'h00000108: r_sin = 32'hFFFFFC1D;
      32'h00000109: r_sin = 32'hFFFFFC1C;
      32'h0000010A: r_sin = 32'hFFFFFC1A;
      32'h0000010B: r_sin = 32'hFFFFFC19;
      32'h0000010C: r_sin = 32'hFFFFFC19;
      32'h0000010D: r_sin = 32'hFFFFFC18;
      32'h0000010E: r_sin = 32'hFFFFFC18;
      32'h0000010F: r_sin = 32'hFFFFFC18;
      32'h00000110: r_sin = 32'hFFFFFC19;
      32'h00000111: r_sin = 32'hFFFFFC19;
      32'h00000112: r_sin = 32'hFFFFFC1A;
      32'h00000113: r_sin = 32'hFFFFFC1C;
      32'h00000114: r_sin = 32'hFFFFFC1D;
      32'h00000115: r_sin = 32'hFFFFFC1F;
      32'h00000116: r_sin = 32'hFFFFFC22;
      32'h00000117: r_sin = 32'hFFFFFC24;
      32'h00000118: r_sin = 32'hFFFFFC27;
      32'h00000119: r_sin = 32'hFFFFFC2A;
      32'h0000011A: r_sin = 32'hFFFFFC2E;
      32'h0000011B: r_sin = 32'hFFFFFC32;
      32'h0000011C: r_sin = 32'hFFFFFC36;
      32'h0000011D: r_sin = 32'hFFFFFC3A;
      32'h0000011E: r_sin = 32'hFFFFFC3F;
      32'h0000011F: r_sin = 32'hFFFFFC44;
      32'h00000120: r_sin = 32'hFFFFFC49;
      32'h00000121: r_sin = 32'hFFFFFC4E;
      32'h00000122: r_sin = 32'hFFFFFC54;
      32'h00000123: r_sin = 32'hFFFFFC5A;
      32'h00000124: r_sin = 32'hFFFFFC61;
      32'h00000125: r_sin = 32'hFFFFFC67;
      32'h00000126: r_sin = 32'hFFFFFC6E;
      32'h00000127: r_sin = 32'hFFFFFC76;
      32'h00000128: r_sin = 32'hFFFFFC7D;
      32'h00000129: r_sin = 32'hFFFFFC85;
      32'h0000012A: r_sin = 32'hFFFFFC8D;
      32'h0000012B: r_sin = 32'hFFFFFC95;
      32'h0000012C: r_sin = 32'hFFFFFC9E;
      32'h0000012D: r_sin = 32'hFFFFFCA7;
      32'h0000012E: r_sin = 32'hFFFFFCB0;
      32'h0000012F: r_sin = 32'hFFFFFCB9;
      32'h00000130: r_sin = 32'hFFFFFCC3;
      32'h00000131: r_sin = 32'hFFFFFCCD;
      32'h00000132: r_sin = 32'hFFFFFCD7;
      32'h00000133: r_sin = 32'hFFFFFCE1;
      32'h00000134: r_sin = 32'hFFFFFCEC;
      32'h00000135: r_sin = 32'hFFFFFCF7;
      32'h00000136: r_sin = 32'hFFFFFD02;
      32'h00000137: r_sin = 32'hFFFFFD0D;
      32'h00000138: r_sin = 32'hFFFFFD19;
      32'h00000139: r_sin = 32'hFFFFFD25;
      32'h0000013A: r_sin = 32'hFFFFFD31;
      32'h0000013B: r_sin = 32'hFFFFFD3D;
      32'h0000013C: r_sin = 32'hFFFFFD49;
      32'h0000013D: r_sin = 32'hFFFFFD56;
      32'h0000013E: r_sin = 32'hFFFFFD63;
      32'h0000013F: r_sin = 32'hFFFFFD70;
      32'h00000140: r_sin = 32'hFFFFFD7D;
      32'h00000141: r_sin = 32'hFFFFFD8B;
      32'h00000142: r_sin = 32'hFFFFFD98;
      32'h00000143: r_sin = 32'hFFFFFDA6;
      32'h00000144: r_sin = 32'hFFFFFDB4;
      32'h00000145: r_sin = 32'hFFFFFDC2;
      32'h00000146: r_sin = 32'hFFFFFDD1;
      32'h00000147: r_sin = 32'hFFFFFDDF;
      32'h00000148: r_sin = 32'hFFFFFDEE;
      32'h00000149: r_sin = 32'hFFFFFDFD;
      32'h0000014A: r_sin = 32'hFFFFFE0C;
      32'h0000014B: r_sin = 32'hFFFFFE1B;
      32'h0000014C: r_sin = 32'hFFFFFE2B;
      32'h0000014D: r_sin = 32'hFFFFFE3A;
      32'h0000014E: r_sin = 32'hFFFFFE4A;
      32'h0000014F: r_sin = 32'hFFFFFE59;
      32'h00000150: r_sin = 32'hFFFFFE69;
      32'h00000151: r_sin = 32'hFFFFFE79;
      32'h00000152: r_sin = 32'hFFFFFE89;
      32'h00000153: r_sin = 32'hFFFFFE9A;
      32'h00000154: r_sin = 32'hFFFFFEAA;
      32'h00000155: r_sin = 32'hFFFFFEBA;
      32'h00000156: r_sin = 32'hFFFFFECB;
      32'h00000157: r_sin = 32'hFFFFFEDC;
      32'h00000158: r_sin = 32'hFFFFFEEC;
      32'h00000159: r_sin = 32'hFFFFFEFD;
      32'h0000015A: r_sin = 32'hFFFFFF0E;
      32'h0000015B: r_sin = 32'hFFFFFF1F;
      32'h0000015C: r_sin = 32'hFFFFFF30;
      32'h0000015D: r_sin = 32'hFFFFFF41;
      32'h0000015E: r_sin = 32'hFFFFFF52;
      32'h0000015F: r_sin = 32'hFFFFFF64;
      32'h00000160: r_sin = 32'hFFFFFF75;
      32'h00000161: r_sin = 32'hFFFFFF86;
      32'h00000162: r_sin = 32'hFFFFFF97;
      32'h00000163: r_sin = 32'hFFFFFFA9;
      32'h00000164: r_sin = 32'hFFFFFFBA;
      32'h00000165: r_sin = 32'hFFFFFFCC;
      32'h00000166: r_sin = 32'hFFFFFFDD;
      32'h00000167: r_sin = 32'hFFFFFFEF;
      32'h00000168: r_sin = 32'h00000000;
      default:      r_sin = 32'h00000000;
endcase

case(i_theta)
      32'hFFFFFF4C: r_cos = 32'hFFFFFC18;
      32'hFFFFFF4D: r_cos = 32'hFFFFFC18;
      32'hFFFFFF4E: r_cos = 32'hFFFFFC19;
      32'hFFFFFF4F: r_cos = 32'hFFFFFC19;
      32'hFFFFFF50: r_cos = 32'hFFFFFC1A;
      32'hFFFFFF51: r_cos = 32'hFFFFFC1C;
      32'hFFFFFF52: r_cos = 32'hFFFFFC1D;
      32'hFFFFFF53: r_cos = 32'hFFFFFC1F;
      32'hFFFFFF54: r_cos = 32'hFFFFFC22;
      32'hFFFFFF55: r_cos = 32'hFFFFFC24;
      32'hFFFFFF56: r_cos = 32'hFFFFFC27;
      32'hFFFFFF57: r_cos = 32'hFFFFFC2A;
      32'hFFFFFF58: r_cos = 32'hFFFFFC2E;
      32'hFFFFFF59: r_cos = 32'hFFFFFC32;
      32'hFFFFFF5A: r_cos = 32'hFFFFFC36;
      32'hFFFFFF5B: r_cos = 32'hFFFFFC3A;
      32'hFFFFFF5C: r_cos = 32'hFFFFFC3F;
      32'hFFFFFF5D: r_cos = 32'hFFFFFC44;
      32'hFFFFFF5E: r_cos = 32'hFFFFFC49;
      32'hFFFFFF5F: r_cos = 32'hFFFFFC4E;
      32'hFFFFFF60: r_cos = 32'hFFFFFC54;
      32'hFFFFFF61: r_cos = 32'hFFFFFC5A;
      32'hFFFFFF62: r_cos = 32'hFFFFFC61;
      32'hFFFFFF63: r_cos = 32'hFFFFFC67;
      32'hFFFFFF64: r_cos = 32'hFFFFFC6E;
      32'hFFFFFF65: r_cos = 32'hFFFFFC76;
      32'hFFFFFF66: r_cos = 32'hFFFFFC7D;
      32'hFFFFFF67: r_cos = 32'hFFFFFC85;
      32'hFFFFFF68: r_cos = 32'hFFFFFC8D;
      32'hFFFFFF69: r_cos = 32'hFFFFFC95;
      32'hFFFFFF6A: r_cos = 32'hFFFFFC9E;
      32'hFFFFFF6B: r_cos = 32'hFFFFFCA7;
      32'hFFFFFF6C: r_cos = 32'hFFFFFCB0;
      32'hFFFFFF6D: r_cos = 32'hFFFFFCB9;
      32'hFFFFFF6E: r_cos = 32'hFFFFFCC3;
      32'hFFFFFF6F: r_cos = 32'hFFFFFCCD;
      32'hFFFFFF70: r_cos = 32'hFFFFFCD7;
      32'hFFFFFF71: r_cos = 32'hFFFFFCE1;
      32'hFFFFFF72: r_cos = 32'hFFFFFCEC;
      32'hFFFFFF73: r_cos = 32'hFFFFFCF7;
      32'hFFFFFF74: r_cos = 32'hFFFFFD02;
      32'hFFFFFF75: r_cos = 32'hFFFFFD0D;
      32'hFFFFFF76: r_cos = 32'hFFFFFD19;
      32'hFFFFFF77: r_cos = 32'hFFFFFD25;
      32'hFFFFFF78: r_cos = 32'hFFFFFD31;
      32'hFFFFFF79: r_cos = 32'hFFFFFD3D;
      32'hFFFFFF7A: r_cos = 32'hFFFFFD49;
      32'hFFFFFF7B: r_cos = 32'hFFFFFD56;
      32'hFFFFFF7C: r_cos = 32'hFFFFFD63;
      32'hFFFFFF7D: r_cos = 32'hFFFFFD70;
      32'hFFFFFF7E: r_cos = 32'hFFFFFD7D;
      32'hFFFFFF7F: r_cos = 32'hFFFFFD8B;
      32'hFFFFFF80: r_cos = 32'hFFFFFD98;
      32'hFFFFFF81: r_cos = 32'hFFFFFDA6;
      32'hFFFFFF82: r_cos = 32'hFFFFFDB4;
      32'hFFFFFF83: r_cos = 32'hFFFFFDC2;
      32'hFFFFFF84: r_cos = 32'hFFFFFDD1;
      32'hFFFFFF85: r_cos = 32'hFFFFFDDF;
      32'hFFFFFF86: r_cos = 32'hFFFFFDEE;
      32'hFFFFFF87: r_cos = 32'hFFFFFDFD;
      32'hFFFFFF88: r_cos = 32'hFFFFFE0C;
      32'hFFFFFF89: r_cos = 32'hFFFFFE1B;
      32'hFFFFFF8A: r_cos = 32'hFFFFFE2B;
      32'hFFFFFF8B: r_cos = 32'hFFFFFE3A;
      32'hFFFFFF8C: r_cos = 32'hFFFFFE4A;
      32'hFFFFFF8D: r_cos = 32'hFFFFFE59;
      32'hFFFFFF8E: r_cos = 32'hFFFFFE69;
      32'hFFFFFF8F: r_cos = 32'hFFFFFE79;
      32'hFFFFFF90: r_cos = 32'hFFFFFE89;
      32'hFFFFFF91: r_cos = 32'hFFFFFE9A;
      32'hFFFFFF92: r_cos = 32'hFFFFFEAA;
      32'hFFFFFF93: r_cos = 32'hFFFFFEBA;
      32'hFFFFFF94: r_cos = 32'hFFFFFECB;
      32'hFFFFFF95: r_cos = 32'hFFFFFEDC;
      32'hFFFFFF96: r_cos = 32'hFFFFFEEC;
      32'hFFFFFF97: r_cos = 32'hFFFFFEFD;
      32'hFFFFFF98: r_cos = 32'hFFFFFF0E;
      32'hFFFFFF99: r_cos = 32'hFFFFFF1F;
      32'hFFFFFF9A: r_cos = 32'hFFFFFF30;
      32'hFFFFFF9B: r_cos = 32'hFFFFFF41;
      32'hFFFFFF9C: r_cos = 32'hFFFFFF52;
      32'hFFFFFF9D: r_cos = 32'hFFFFFF64;
      32'hFFFFFF9E: r_cos = 32'hFFFFFF75;
      32'hFFFFFF9F: r_cos = 32'hFFFFFF86;
      32'hFFFFFFA0: r_cos = 32'hFFFFFF97;
      32'hFFFFFFA1: r_cos = 32'hFFFFFFA9;
      32'hFFFFFFA2: r_cos = 32'hFFFFFFBA;
      32'hFFFFFFA3: r_cos = 32'hFFFFFFCC;
      32'hFFFFFFA4: r_cos = 32'hFFFFFFDD;
      32'hFFFFFFA5: r_cos = 32'hFFFFFFEF;
      32'hFFFFFFA6: r_cos = 32'h00000000;
      32'hFFFFFFA7: r_cos = 32'h00000011;
      32'hFFFFFFA8: r_cos = 32'h00000023;
      32'hFFFFFFA9: r_cos = 32'h00000034;
      32'hFFFFFFAA: r_cos = 32'h00000046;
      32'hFFFFFFAB: r_cos = 32'h00000057;
      32'hFFFFFFAC: r_cos = 32'h00000069;
      32'hFFFFFFAD: r_cos = 32'h0000007A;
      32'hFFFFFFAE: r_cos = 32'h0000008B;
      32'hFFFFFFAF: r_cos = 32'h0000009C;
      32'hFFFFFFB0: r_cos = 32'h000000AE;
      32'hFFFFFFB1: r_cos = 32'h000000BF;
      32'hFFFFFFB2: r_cos = 32'h000000D0;
      32'hFFFFFFB3: r_cos = 32'h000000E1;
      32'hFFFFFFB4: r_cos = 32'h000000F2;
      32'hFFFFFFB5: r_cos = 32'h00000103;
      32'hFFFFFFB6: r_cos = 32'h00000114;
      32'hFFFFFFB7: r_cos = 32'h00000124;
      32'hFFFFFFB8: r_cos = 32'h00000135;
      32'hFFFFFFB9: r_cos = 32'h00000146;
      32'hFFFFFFBA: r_cos = 32'h00000156;
      32'hFFFFFFBB: r_cos = 32'h00000166;
      32'hFFFFFFBC: r_cos = 32'h00000177;
      32'hFFFFFFBD: r_cos = 32'h00000187;
      32'hFFFFFFBE: r_cos = 32'h00000197;
      32'hFFFFFFBF: r_cos = 32'h000001A7;
      32'hFFFFFFC0: r_cos = 32'h000001B6;
      32'hFFFFFFC1: r_cos = 32'h000001C6;
      32'hFFFFFFC2: r_cos = 32'h000001D5;
      32'hFFFFFFC3: r_cos = 32'h000001E5;
      32'hFFFFFFC4: r_cos = 32'h000001F4;
      32'hFFFFFFC5: r_cos = 32'h00000203;
      32'hFFFFFFC6: r_cos = 32'h00000212;
      32'hFFFFFFC7: r_cos = 32'h00000221;
      32'hFFFFFFC8: r_cos = 32'h0000022F;
      32'hFFFFFFC9: r_cos = 32'h0000023E;
      32'hFFFFFFCA: r_cos = 32'h0000024C;
      32'hFFFFFFCB: r_cos = 32'h0000025A;
      32'hFFFFFFCC: r_cos = 32'h00000268;
      32'hFFFFFFCD: r_cos = 32'h00000275;
      32'hFFFFFFCE: r_cos = 32'h00000283;
      32'hFFFFFFCF: r_cos = 32'h00000290;
      32'hFFFFFFD0: r_cos = 32'h0000029D;
      32'hFFFFFFD1: r_cos = 32'h000002AA;
      32'hFFFFFFD2: r_cos = 32'h000002B7;
      32'hFFFFFFD3: r_cos = 32'h000002C3;
      32'hFFFFFFD4: r_cos = 32'h000002CF;
      32'hFFFFFFD5: r_cos = 32'h000002DB;
      32'hFFFFFFD6: r_cos = 32'h000002E7;
      32'hFFFFFFD7: r_cos = 32'h000002F3;
      32'hFFFFFFD8: r_cos = 32'h000002FE;
      32'hFFFFFFD9: r_cos = 32'h00000309;
      32'hFFFFFFDA: r_cos = 32'h00000314;
      32'hFFFFFFDB: r_cos = 32'h0000031F;
      32'hFFFFFFDC: r_cos = 32'h00000329;
      32'hFFFFFFDD: r_cos = 32'h00000333;
      32'hFFFFFFDE: r_cos = 32'h0000033D;
      32'hFFFFFFDF: r_cos = 32'h00000347;
      32'hFFFFFFE0: r_cos = 32'h00000350;
      32'hFFFFFFE1: r_cos = 32'h00000359;
      32'hFFFFFFE2: r_cos = 32'h00000362;
      32'hFFFFFFE3: r_cos = 32'h0000036B;
      32'hFFFFFFE4: r_cos = 32'h00000373;
      32'hFFFFFFE5: r_cos = 32'h0000037B;
      32'hFFFFFFE6: r_cos = 32'h00000383;
      32'hFFFFFFE7: r_cos = 32'h0000038A;
      32'hFFFFFFE8: r_cos = 32'h00000392;
      32'hFFFFFFE9: r_cos = 32'h00000399;
      32'hFFFFFFEA: r_cos = 32'h0000039F;
      32'hFFFFFFEB: r_cos = 32'h000003A6;
      32'hFFFFFFEC: r_cos = 32'h000003AC;
      32'hFFFFFFED: r_cos = 32'h000003B2;
      32'hFFFFFFEE: r_cos = 32'h000003B7;
      32'hFFFFFFEF: r_cos = 32'h000003BC;
      32'hFFFFFFF0: r_cos = 32'h000003C1;
      32'hFFFFFFF1: r_cos = 32'h000003C6;
      32'hFFFFFFF2: r_cos = 32'h000003CA;
      32'hFFFFFFF3: r_cos = 32'h000003CE;
      32'hFFFFFFF4: r_cos = 32'h000003D2;
      32'hFFFFFFF5: r_cos = 32'h000003D6;
      32'hFFFFFFF6: r_cos = 32'h000003D9;
      32'hFFFFFFF7: r_cos = 32'h000003DC;
      32'hFFFFFFF8: r_cos = 32'h000003DE;
      32'hFFFFFFF9: r_cos = 32'h000003E1;
      32'hFFFFFFFA: r_cos = 32'h000003E3;
      32'hFFFFFFFB: r_cos = 32'h000003E4;
      32'hFFFFFFFC: r_cos = 32'h000003E6;
      32'hFFFFFFFD: r_cos = 32'h000003E7;
      32'hFFFFFFFE: r_cos = 32'h000003E7;
      32'hFFFFFFFF: r_cos = 32'h000003E8;
      32'h00000000: r_cos = 32'h000003E8;
      32'h00000001: r_cos = 32'h000003E8;
      32'h00000002: r_cos = 32'h000003E7;
      32'h00000003: r_cos = 32'h000003E7;
      32'h00000004: r_cos = 32'h000003E6;
      32'h00000005: r_cos = 32'h000003E4;
      32'h00000006: r_cos = 32'h000003E3;
      32'h00000007: r_cos = 32'h000003E1;
      32'h00000008: r_cos = 32'h000003DE;
      32'h00000009: r_cos = 32'h000003DC;
      32'h0000000A: r_cos = 32'h000003D9;
      32'h0000000B: r_cos = 32'h000003D6;
      32'h0000000C: r_cos = 32'h000003D2;
      32'h0000000D: r_cos = 32'h000003CE;
      32'h0000000E: r_cos = 32'h000003CA;
      32'h0000000F: r_cos = 32'h000003C6;
      32'h00000010: r_cos = 32'h000003C1;
      32'h00000011: r_cos = 32'h000003BC;
      32'h00000012: r_cos = 32'h000003B7;
      32'h00000013: r_cos = 32'h000003B2;
      32'h00000014: r_cos = 32'h000003AC;
      32'h00000015: r_cos = 32'h000003A6;
      32'h00000016: r_cos = 32'h0000039F;
      32'h00000017: r_cos = 32'h00000399;
      32'h00000018: r_cos = 32'h00000392;
      32'h00000019: r_cos = 32'h0000038A;
      32'h0000001A: r_cos = 32'h00000383;
      32'h0000001B: r_cos = 32'h0000037B;
      32'h0000001C: r_cos = 32'h00000373;
      32'h0000001D: r_cos = 32'h0000036B;
      32'h0000001E: r_cos = 32'h00000362;
      32'h0000001F: r_cos = 32'h00000359;
      32'h00000020: r_cos = 32'h00000350;
      32'h00000021: r_cos = 32'h00000347;
      32'h00000022: r_cos = 32'h0000033D;
      32'h00000023: r_cos = 32'h00000333;
      32'h00000024: r_cos = 32'h00000329;
      32'h00000025: r_cos = 32'h0000031F;
      32'h00000026: r_cos = 32'h00000314;
      32'h00000027: r_cos = 32'h00000309;
      32'h00000028: r_cos = 32'h000002FE;
      32'h00000029: r_cos = 32'h000002F3;
      32'h0000002A: r_cos = 32'h000002E7;
      32'h0000002B: r_cos = 32'h000002DB;
      32'h0000002C: r_cos = 32'h000002CF;
      32'h0000002D: r_cos = 32'h000002C3;
      32'h0000002E: r_cos = 32'h000002B7;
      32'h0000002F: r_cos = 32'h000002AA;
      32'h00000030: r_cos = 32'h0000029D;
      32'h00000031: r_cos = 32'h00000290;
      32'h00000032: r_cos = 32'h00000283;
      32'h00000033: r_cos = 32'h00000275;
      32'h00000034: r_cos = 32'h00000268;
      32'h00000035: r_cos = 32'h0000025A;
      32'h00000036: r_cos = 32'h0000024C;
      32'h00000037: r_cos = 32'h0000023E;
      32'h00000038: r_cos = 32'h0000022F;
      32'h00000039: r_cos = 32'h00000221;
      32'h0000003A: r_cos = 32'h00000212;
      32'h0000003B: r_cos = 32'h00000203;
      32'h0000003C: r_cos = 32'h000001F4;
      32'h0000003D: r_cos = 32'h000001E5;
      32'h0000003E: r_cos = 32'h000001D5;
      32'h0000003F: r_cos = 32'h000001C6;
      32'h00000040: r_cos = 32'h000001B6;
      32'h00000041: r_cos = 32'h000001A7;
      32'h00000042: r_cos = 32'h00000197;
      32'h00000043: r_cos = 32'h00000187;
      32'h00000044: r_cos = 32'h00000177;
      32'h00000045: r_cos = 32'h00000166;
      32'h00000046: r_cos = 32'h00000156;
      32'h00000047: r_cos = 32'h00000146;
      32'h00000048: r_cos = 32'h00000135;
      32'h00000049: r_cos = 32'h00000124;
      32'h0000004A: r_cos = 32'h00000114;
      32'h0000004B: r_cos = 32'h00000103;
      32'h0000004C: r_cos = 32'h000000F2;
      32'h0000004D: r_cos = 32'h000000E1;
      32'h0000004E: r_cos = 32'h000000D0;
      32'h0000004F: r_cos = 32'h000000BF;
      32'h00000050: r_cos = 32'h000000AE;
      32'h00000051: r_cos = 32'h0000009C;
      32'h00000052: r_cos = 32'h0000008B;
      32'h00000053: r_cos = 32'h0000007A;
      32'h00000054: r_cos = 32'h00000069;
      32'h00000055: r_cos = 32'h00000057;
      32'h00000056: r_cos = 32'h00000046;
      32'h00000057: r_cos = 32'h00000034;
      32'h00000058: r_cos = 32'h00000023;
      32'h00000059: r_cos = 32'h00000011;
      32'h0000005A: r_cos = 32'h00000000;
      32'h0000005B: r_cos = 32'hFFFFFFEF;
      32'h0000005C: r_cos = 32'hFFFFFFDD;
      32'h0000005D: r_cos = 32'hFFFFFFCC;
      32'h0000005E: r_cos = 32'hFFFFFFBA;
      32'h0000005F: r_cos = 32'hFFFFFFA9;
      32'h00000060: r_cos = 32'hFFFFFF97;
      32'h00000061: r_cos = 32'hFFFFFF86;
      32'h00000062: r_cos = 32'hFFFFFF75;
      32'h00000063: r_cos = 32'hFFFFFF64;
      32'h00000064: r_cos = 32'hFFFFFF52;
      32'h00000065: r_cos = 32'hFFFFFF41;
      32'h00000066: r_cos = 32'hFFFFFF30;
      32'h00000067: r_cos = 32'hFFFFFF1F;
      32'h00000068: r_cos = 32'hFFFFFF0E;
      32'h00000069: r_cos = 32'hFFFFFEFD;
      32'h0000006A: r_cos = 32'hFFFFFEEC;
      32'h0000006B: r_cos = 32'hFFFFFEDC;
      32'h0000006C: r_cos = 32'hFFFFFECB;
      32'h0000006D: r_cos = 32'hFFFFFEBA;
      32'h0000006E: r_cos = 32'hFFFFFEAA;
      32'h0000006F: r_cos = 32'hFFFFFE9A;
      32'h00000070: r_cos = 32'hFFFFFE89;
      32'h00000071: r_cos = 32'hFFFFFE79;
      32'h00000072: r_cos = 32'hFFFFFE69;
      32'h00000073: r_cos = 32'hFFFFFE59;
      32'h00000074: r_cos = 32'hFFFFFE4A;
      32'h00000075: r_cos = 32'hFFFFFE3A;
      32'h00000076: r_cos = 32'hFFFFFE2B;
      32'h00000077: r_cos = 32'hFFFFFE1B;
      32'h00000078: r_cos = 32'hFFFFFE0C;
      32'h00000079: r_cos = 32'hFFFFFDFD;
      32'h0000007A: r_cos = 32'hFFFFFDEE;
      32'h0000007B: r_cos = 32'hFFFFFDDF;
      32'h0000007C: r_cos = 32'hFFFFFDD1;
      32'h0000007D: r_cos = 32'hFFFFFDC2;
      32'h0000007E: r_cos = 32'hFFFFFDB4;
      32'h0000007F: r_cos = 32'hFFFFFDA6;
      32'h00000080: r_cos = 32'hFFFFFD98;
      32'h00000081: r_cos = 32'hFFFFFD8B;
      32'h00000082: r_cos = 32'hFFFFFD7D;
      32'h00000083: r_cos = 32'hFFFFFD70;
      32'h00000084: r_cos = 32'hFFFFFD63;
      32'h00000085: r_cos = 32'hFFFFFD56;
      32'h00000086: r_cos = 32'hFFFFFD49;
      32'h00000087: r_cos = 32'hFFFFFD3D;
      32'h00000088: r_cos = 32'hFFFFFD31;
      32'h00000089: r_cos = 32'hFFFFFD25;
      32'h0000008A: r_cos = 32'hFFFFFD19;
      32'h0000008B: r_cos = 32'hFFFFFD0D;
      32'h0000008C: r_cos = 32'hFFFFFD02;
      32'h0000008D: r_cos = 32'hFFFFFCF7;
      32'h0000008E: r_cos = 32'hFFFFFCEC;
      32'h0000008F: r_cos = 32'hFFFFFCE1;
      32'h00000090: r_cos = 32'hFFFFFCD7;
      32'h00000091: r_cos = 32'hFFFFFCCD;
      32'h00000092: r_cos = 32'hFFFFFCC3;
      32'h00000093: r_cos = 32'hFFFFFCB9;
      32'h00000094: r_cos = 32'hFFFFFCB0;
      32'h00000095: r_cos = 32'hFFFFFCA7;
      32'h00000096: r_cos = 32'hFFFFFC9E;
      32'h00000097: r_cos = 32'hFFFFFC95;
      32'h00000098: r_cos = 32'hFFFFFC8D;
      32'h00000099: r_cos = 32'hFFFFFC85;
      32'h0000009A: r_cos = 32'hFFFFFC7D;
      32'h0000009B: r_cos = 32'hFFFFFC76;
      32'h0000009C: r_cos = 32'hFFFFFC6E;
      32'h0000009D: r_cos = 32'hFFFFFC67;
      32'h0000009E: r_cos = 32'hFFFFFC61;
      32'h0000009F: r_cos = 32'hFFFFFC5A;
      32'h000000A0: r_cos = 32'hFFFFFC54;
      32'h000000A1: r_cos = 32'hFFFFFC4E;
      32'h000000A2: r_cos = 32'hFFFFFC49;
      32'h000000A3: r_cos = 32'hFFFFFC44;
      32'h000000A4: r_cos = 32'hFFFFFC3F;
      32'h000000A5: r_cos = 32'hFFFFFC3A;
      32'h000000A6: r_cos = 32'hFFFFFC36;
      32'h000000A7: r_cos = 32'hFFFFFC32;
      32'h000000A8: r_cos = 32'hFFFFFC2E;
      32'h000000A9: r_cos = 32'hFFFFFC2A;
      32'h000000AA: r_cos = 32'hFFFFFC27;
      32'h000000AB: r_cos = 32'hFFFFFC24;
      32'h000000AC: r_cos = 32'hFFFFFC22;
      32'h000000AD: r_cos = 32'hFFFFFC1F;
      32'h000000AE: r_cos = 32'hFFFFFC1D;
      32'h000000AF: r_cos = 32'hFFFFFC1C;
      32'h000000B0: r_cos = 32'hFFFFFC1A;
      32'h000000B1: r_cos = 32'hFFFFFC19;
      32'h000000B2: r_cos = 32'hFFFFFC19;
      32'h000000B3: r_cos = 32'hFFFFFC18;
      32'h000000B4: r_cos = 32'hFFFFFC18;
      32'h000000B5: r_cos = 32'hFFFFFC18;
      32'h000000B6: r_cos = 32'hFFFFFC19;
      32'h000000B7: r_cos = 32'hFFFFFC19;
      32'h000000B8: r_cos = 32'hFFFFFC1A;
      32'h000000B9: r_cos = 32'hFFFFFC1C;
      32'h000000BA: r_cos = 32'hFFFFFC1D;
      32'h000000BB: r_cos = 32'hFFFFFC1F;
      32'h000000BC: r_cos = 32'hFFFFFC22;
      32'h000000BD: r_cos = 32'hFFFFFC24;
      32'h000000BE: r_cos = 32'hFFFFFC27;
      32'h000000BF: r_cos = 32'hFFFFFC2A;
      32'h000000C0: r_cos = 32'hFFFFFC2E;
      32'h000000C1: r_cos = 32'hFFFFFC32;
      32'h000000C2: r_cos = 32'hFFFFFC36;
      32'h000000C3: r_cos = 32'hFFFFFC3A;
      32'h000000C4: r_cos = 32'hFFFFFC3F;
      32'h000000C5: r_cos = 32'hFFFFFC44;
      32'h000000C6: r_cos = 32'hFFFFFC49;
      32'h000000C7: r_cos = 32'hFFFFFC4E;
      32'h000000C8: r_cos = 32'hFFFFFC54;
      32'h000000C9: r_cos = 32'hFFFFFC5A;
      32'h000000CA: r_cos = 32'hFFFFFC61;
      32'h000000CB: r_cos = 32'hFFFFFC67;
      32'h000000CC: r_cos = 32'hFFFFFC6E;
      32'h000000CD: r_cos = 32'hFFFFFC76;
      32'h000000CE: r_cos = 32'hFFFFFC7D;
      32'h000000CF: r_cos = 32'hFFFFFC85;
      32'h000000D0: r_cos = 32'hFFFFFC8D;
      32'h000000D1: r_cos = 32'hFFFFFC95;
      32'h000000D2: r_cos = 32'hFFFFFC9E;
      32'h000000D3: r_cos = 32'hFFFFFCA7;
      32'h000000D4: r_cos = 32'hFFFFFCB0;
      32'h000000D5: r_cos = 32'hFFFFFCB9;
      32'h000000D6: r_cos = 32'hFFFFFCC3;
      32'h000000D7: r_cos = 32'hFFFFFCCD;
      32'h000000D8: r_cos = 32'hFFFFFCD7;
      32'h000000D9: r_cos = 32'hFFFFFCE1;
      32'h000000DA: r_cos = 32'hFFFFFCEC;
      32'h000000DB: r_cos = 32'hFFFFFCF7;
      32'h000000DC: r_cos = 32'hFFFFFD02;
      32'h000000DD: r_cos = 32'hFFFFFD0D;
      32'h000000DE: r_cos = 32'hFFFFFD19;
      32'h000000DF: r_cos = 32'hFFFFFD25;
      32'h000000E0: r_cos = 32'hFFFFFD31;
      32'h000000E1: r_cos = 32'hFFFFFD3D;
      32'h000000E2: r_cos = 32'hFFFFFD49;
      32'h000000E3: r_cos = 32'hFFFFFD56;
      32'h000000E4: r_cos = 32'hFFFFFD63;
      32'h000000E5: r_cos = 32'hFFFFFD70;
      32'h000000E6: r_cos = 32'hFFFFFD7D;
      32'h000000E7: r_cos = 32'hFFFFFD8B;
      32'h000000E8: r_cos = 32'hFFFFFD98;
      32'h000000E9: r_cos = 32'hFFFFFDA6;
      32'h000000EA: r_cos = 32'hFFFFFDB4;
      32'h000000EB: r_cos = 32'hFFFFFDC2;
      32'h000000EC: r_cos = 32'hFFFFFDD1;
      32'h000000ED: r_cos = 32'hFFFFFDDF;
      32'h000000EE: r_cos = 32'hFFFFFDEE;
      32'h000000EF: r_cos = 32'hFFFFFDFD;
      32'h000000F0: r_cos = 32'hFFFFFE0C;
      32'h000000F1: r_cos = 32'hFFFFFE1B;
      32'h000000F2: r_cos = 32'hFFFFFE2B;
      32'h000000F3: r_cos = 32'hFFFFFE3A;
      32'h000000F4: r_cos = 32'hFFFFFE4A;
      32'h000000F5: r_cos = 32'hFFFFFE59;
      32'h000000F6: r_cos = 32'hFFFFFE69;
      32'h000000F7: r_cos = 32'hFFFFFE79;
      32'h000000F8: r_cos = 32'hFFFFFE89;
      32'h000000F9: r_cos = 32'hFFFFFE9A;
      32'h000000FA: r_cos = 32'hFFFFFEAA;
      32'h000000FB: r_cos = 32'hFFFFFEBA;
      32'h000000FC: r_cos = 32'hFFFFFECB;
      32'h000000FD: r_cos = 32'hFFFFFEDC;
      32'h000000FE: r_cos = 32'hFFFFFEEC;
      32'h000000FF: r_cos = 32'hFFFFFEFD;
      32'h00000100: r_cos = 32'hFFFFFF0E;
      32'h00000101: r_cos = 32'hFFFFFF1F;
      32'h00000102: r_cos = 32'hFFFFFF30;
      32'h00000103: r_cos = 32'hFFFFFF41;
      32'h00000104: r_cos = 32'hFFFFFF52;
      32'h00000105: r_cos = 32'hFFFFFF64;
      32'h00000106: r_cos = 32'hFFFFFF75;
      32'h00000107: r_cos = 32'hFFFFFF86;
      32'h00000108: r_cos = 32'hFFFFFF97;
      32'h00000109: r_cos = 32'hFFFFFFA9;
      32'h0000010A: r_cos = 32'hFFFFFFBA;
      32'h0000010B: r_cos = 32'hFFFFFFCC;
      32'h0000010C: r_cos = 32'hFFFFFFDD;
      32'h0000010D: r_cos = 32'hFFFFFFEF;
      32'h0000010E: r_cos = 32'h00000000;
      32'h0000010F: r_cos = 32'h00000011;
      32'h00000110: r_cos = 32'h00000023;
      32'h00000111: r_cos = 32'h00000034;
      32'h00000112: r_cos = 32'h00000046;
      32'h00000113: r_cos = 32'h00000057;
      32'h00000114: r_cos = 32'h00000069;
      32'h00000115: r_cos = 32'h0000007A;
      32'h00000116: r_cos = 32'h0000008B;
      32'h00000117: r_cos = 32'h0000009C;
      32'h00000118: r_cos = 32'h000000AE;
      32'h00000119: r_cos = 32'h000000BF;
      32'h0000011A: r_cos = 32'h000000D0;
      32'h0000011B: r_cos = 32'h000000E1;
      32'h0000011C: r_cos = 32'h000000F2;
      32'h0000011D: r_cos = 32'h00000103;
      32'h0000011E: r_cos = 32'h00000114;
      32'h0000011F: r_cos = 32'h00000124;
      32'h00000120: r_cos = 32'h00000135;
      32'h00000121: r_cos = 32'h00000146;
      32'h00000122: r_cos = 32'h00000156;
      32'h00000123: r_cos = 32'h00000166;
      32'h00000124: r_cos = 32'h00000177;
      32'h00000125: r_cos = 32'h00000187;
      32'h00000126: r_cos = 32'h00000197;
      32'h00000127: r_cos = 32'h000001A7;
      32'h00000128: r_cos = 32'h000001B6;
      32'h00000129: r_cos = 32'h000001C6;
      32'h0000012A: r_cos = 32'h000001D5;
      32'h0000012B: r_cos = 32'h000001E5;
      32'h0000012C: r_cos = 32'h000001F4;
      32'h0000012D: r_cos = 32'h00000203;
      32'h0000012E: r_cos = 32'h00000212;
      32'h0000012F: r_cos = 32'h00000221;
      32'h00000130: r_cos = 32'h0000022F;
      32'h00000131: r_cos = 32'h0000023E;
      32'h00000132: r_cos = 32'h0000024C;
      32'h00000133: r_cos = 32'h0000025A;
      32'h00000134: r_cos = 32'h00000268;
      32'h00000135: r_cos = 32'h00000275;
      32'h00000136: r_cos = 32'h00000283;
      32'h00000137: r_cos = 32'h00000290;
      32'h00000138: r_cos = 32'h0000029D;
      32'h00000139: r_cos = 32'h000002AA;
      32'h0000013A: r_cos = 32'h000002B7;
      32'h0000013B: r_cos = 32'h000002C3;
      32'h0000013C: r_cos = 32'h000002CF;
      32'h0000013D: r_cos = 32'h000002DB;
      32'h0000013E: r_cos = 32'h000002E7;
      32'h0000013F: r_cos = 32'h000002F3;
      32'h00000140: r_cos = 32'h000002FE;
      32'h00000141: r_cos = 32'h00000309;
      32'h00000142: r_cos = 32'h00000314;
      32'h00000143: r_cos = 32'h0000031F;
      32'h00000144: r_cos = 32'h00000329;
      32'h00000145: r_cos = 32'h00000333;
      32'h00000146: r_cos = 32'h0000033D;
      32'h00000147: r_cos = 32'h00000347;
      32'h00000148: r_cos = 32'h00000350;
      32'h00000149: r_cos = 32'h00000359;
      32'h0000014A: r_cos = 32'h00000362;
      32'h0000014B: r_cos = 32'h0000036B;
      32'h0000014C: r_cos = 32'h00000373;
      32'h0000014D: r_cos = 32'h0000037B;
      32'h0000014E: r_cos = 32'h00000383;
      32'h0000014F: r_cos = 32'h0000038A;
      32'h00000150: r_cos = 32'h00000392;
      32'h00000151: r_cos = 32'h00000399;
      32'h00000152: r_cos = 32'h0000039F;
      32'h00000153: r_cos = 32'h000003A6;
      32'h00000154: r_cos = 32'h000003AC;
      32'h00000155: r_cos = 32'h000003B2;
      32'h00000156: r_cos = 32'h000003B7;
      32'h00000157: r_cos = 32'h000003BC;
      32'h00000158: r_cos = 32'h000003C1;
      32'h00000159: r_cos = 32'h000003C6;
      32'h0000015A: r_cos = 32'h000003CA;
      32'h0000015B: r_cos = 32'h000003CE;
      32'h0000015C: r_cos = 32'h000003D2;
      32'h0000015D: r_cos = 32'h000003D6;
      32'h0000015E: r_cos = 32'h000003D9;
      32'h0000015F: r_cos = 32'h000003DC;
      32'h00000160: r_cos = 32'h000003DE;
      32'h00000161: r_cos = 32'h000003E1;
      32'h00000162: r_cos = 32'h000003E3;
      32'h00000163: r_cos = 32'h000003E4;
      32'h00000164: r_cos = 32'h000003E6;
      32'h00000165: r_cos = 32'h000003E7;
      32'h00000166: r_cos = 32'h000003E7;
      32'h00000167: r_cos = 32'h000003E8;
      32'h00000168: r_cos = 32'h000003E8; // 360deg
      default:      r_cos = 32'h00000000;
endcase

end


endmodule