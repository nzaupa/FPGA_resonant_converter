// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
jRUPhLmqH2VHmNicFybkd60oOzUUEW3Isas/71nABSyc0XKTZlMo66KLqYcHwBhw7IEfLGccQDm0
FfIHsjoDSY4abTlwBTtZ46gIsDsYzeHJDt6YjMgHHEXfOJQ3t4sPNy56oB9vUUlwtpMC0XeeRiBl
Cd7oziv/cUJl0qdWXThQNcn7opP92n8fQqqmqYpYUPn3FO/Bsg8xdsQdm5qyemaXlby151VJ8g1P
I6X1LPYtcYOIMCzXFREjvSze1UVkP1A1zBB+pRdAfk467nV8T7+omj8mQwvdT8DwDkI1mm4VcIAK
7bZrZiS6FEvrgEs3SP8e7UQZZqav1aKbyViPkw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3024)
Bp7NFmyWe35mQlwkYS465vNhiScgnjpfGQUVSg23QPPYEWI12GnTqS5xoL8CXrWyMebPCdgz8E2m
OnU8ndCi1s9Jzr/BpvwHKITR9VEyo6dz4EVIPjrF6PYIdxL08XKDitg0SZHcD+eSqSPZhGvd5vJ3
XSdma0RbyK8IDb2PaFISHuNFFSjeDAKGT+ICv7Erlx0wo8q5sZWDXJt/RNyTIzO73gNnzcB98Qr5
+Eqvq3L2u+ID6GZgJp8Jh8p03/S6lw6KCVXfRsf4Rx2VXEIJfcPV7sIDVvmYVUkEQ9RLO0+kcYvl
1bjSvGruFsHKm3I33yfywtkyhDymayPAo/bL8zuwPJouAbR25zRTa7e5PSf52rtQZqVaYc0s54Sv
jubSD7JLTwIDOmwtzosfA+9ZeD/nlPVjfQBZHRVKGfcXWuFPLVhAHC00DwU+SvY5zdsHgWpeYBuv
cVKHaA/Ao7+SBK28xf0FtZ8t3IaeaJ0PbcHP1BgI0U8RIxXKYEgXvXKcXGsw1oSMtKKztwqEbsgL
Yk7Ww6Fx0t8ihac6XLnA7YARGt3E3Enp3LwqPNEAMePF5hyVoTHbBc7+xJRZtdhyeBs8KcDAUc0I
3UpkZ9PBZx6O9hHwCjYv+MsZ3T3UiRtq3UcCzLGMvb4ZY474XVWBUFEUtaNcs803JHHtCHbe6HU9
dlwcZb2JezlDTr/RWrUEJzeZe9ncbdV1Ge0tVZo9xkHyn4OGFiyWj4VhKk0rYzR16o+kCn22ALfT
gYuzxAxypgYTFCrLM66/55FVlaUB6u+8unoCL0efYFKVyTOIoqrPFG0IVd5cVueoD3tAwCnSDv6F
HsGFvYtLBB4qMGn8MqQMw6+hnV0DOdIpzAQTar8wXmTybYT+V9SUrzuy8DMerAjWw56eZm/Mj0ZD
r60ecC/MUx3FDlelZBzVg5MyFQQRfcJBRnCaX7WrvCNqp52k97CfJEItIsv0bYOEH2AgSgXkJh8z
t4iN4DOmdPEgWdVWEhPwKeuIyMBYLIAgN+VPbctxxENmDlLgODXNifNehOdz21a396ZTu+5f7oLS
ULHbqDGeKcBIKu83yLxmcfZbfPl9gf/e0tHA9K9a47CYcg+FSjoYekUEH/BMLYTcE352n+5DQ6Hk
5hoBhyvi8l7N6kWD3h9e3Gn3mIvzWazNV6lLlezUtiHyuVjTpHiTe6AWwTj/hcINAOf8FFciUNdi
Qi8eL8wz6wPhl96v96IUWEvsjvwK3C35B7Coas3onzs3JfiPGQcctu1iWHDYnES/Q7Va4WtMjk+I
PsVZ0mpm33XmLYhDBxy0m4vxLQOdCFZNOIwNMMsDniffLgEm1/w8XDXX/q4+hWMRNWIdLwcPAkm3
Y9Ix98hn1j7ja6PjfzCOluDYXXhmfTUxgL0SrtN1AFsN0CAIfSaZhjPaoEmubS5/fPzq8XDlbvKi
AMK1IqSzeF6pb27Ntzg52SUaKOm7b29FmhyDIUIzIWC0fuZ9XJM10ALd/LKXzsSaCNTDnilxYHMp
j0RgjGRzAneyA9ZwhFQUGjuqZjQkXDkN9FgKcQdWvt7s6i2YQ5CvBjcXkhj89L776w0RxR8tYaB6
JHUW+cI+KM4OtxWfTwZ7nEuyymSl5iU0DoIvqS2DL6dxBXg231h2rjtTAurS3k3p+UhZVP8RgH7u
GbE41ckP4SL+dpO6/DG5kczBeDph0Pm086UD6t5ucF44YWW2Gh8D9Ev88evxoMMH/6RD0qH3fHAg
7SsGSk/w3mIe77ruDdzlKWcg4t865uxllm4uaUPm5daGvas8TiTUWw29wlxOrfAZ7qLrPmRzINs7
KeIjA+6lx+DIPO/L/EjglniFYw+91Tq+3+CwUUaUZ4uBXwqjiRDStWV9GpZt+jCLFd7Ma056EpJq
FczrwB1Aayve0FxiXiqHpE23WpdY0g1QtNfwanRAK9AIuspYS6ruEgDZraLsrlOhUDufiTHXFHU3
ydeZ8apLSWhKND5zQt781bX19NUzJI0DYHywNyfNNNMaaaJDNy+iFjyQXFRANuqOHEKeMmTVEzo6
b/+IFyrh0UwyXgYZDzmnuQKnesJegvyTvZuG1YUMOe41aKWYpnLWahLzDE0bAwKgHEiShKYTMNnX
lrokrwdsM/eeGTPWubMWZM332yLf7Zg34oyhzBXZFkfDlqGHRRXj4IZSLpWXEm6UbLbUCQWCWeRJ
Fch6l9IEreZbBQtZ3/GvuUArDvLkBrJjV/+J9lN+ff4jFQHhVAZ3m6lIbHPrOB9LcR09yOMiTbrh
Y4VVpuURi1r6SWVggRyrhuT/BWHYIlQ88K7JcVVkG+n39O6QblvVV6k4hvck/K77EvUxdNiYLPe/
aP9hH3STPZkJJuD7SaCN26OI0SQHSJnsU4xv9q704eHwiQjfqbxaPjSCR7xkFSC/pXGrrs9Jia7Y
CssPmMZcjjcG+3ouyhQ4P3T0fc6jzDN0Qh1gW1YWwRoUWiK82q9rr2C/zHPu/Zz7DWmmLB0p5M60
nTAwgNK2B8Aio0THdZsPee5f0G9BLiqevNZOE0NG4Uq9qXyx+QEqlD4ifSJUdQFBIQOGPTjcoPpt
G10lxz4ViWjjhvnD7wEjoEjzq4VEpe+laqdIsQJQQTvSDsmvRp23neh4boxrbUUfONq/Hd9a6IEP
xM/W6x/tsaRgAv6GfsLozUoC8SsDgssazFBvZzu05C6WWpvRzinFJQiQOYpds6LssKC1XzXkEMmd
NxWzwNohpjHtwtrQFfHVESmvxB4FIy5CE6Adzgohxb/zpmtslFBBaRMbXnq4PD8bAhO1HlOUhBwT
qlNvV/QiAxD/VAJBCohDOq8vZZgQBjD8XJRuT2wx1GebwurROh7QqxU+gXDav/nCG8IH93WuBPjr
nP6M3teqylKT78eAUcZrSEgCBQpLC7wCS9YAvVVA1HFJE1f6uFtPpLbKgn1IlAdHqVPOlZAnc8bZ
nvsZsz+tmBBKFK75gZUL80FukophLHUtlUIG0EYEqmu0kgYva0qn0S7htXFeSWI410OxrLOFi5SS
O/YXZmnlzeblFkt9e63BxUgVC9QH2U4wLFdWUhBSVrePRFVCc1X0E8gzLhxxRKZhBi1RNxjytbVY
aP9dpmnQ5fIzNzfrkqQf2Jh6/FcSyPB4CB4Alxa1JCcjtcpz0NLMD3Izl7Ezq0lrx4xuaW5un1DG
inhTT3VyHL0+yBU7SvTfKDNeDjTZNBYTwAaWZO2A45r7+4pINpo+qRZPOiqGZFCufU8r7yCkJV3n
nj7ttrcYzN/nqexOQyYVfGGXwJ5iuvlTW0FotzhVtFcoaYP892n4lK67vcntjrhze6JJIkWAN8tv
MhYTJlsF5LDSIWKOrUKYVdLkZf0VDpzoUvSFoxChEOUk4rWvzNmYVfYdZUI6Iy7E+hQ4b6BTYmRA
sxFABRouBUDHKwKRtcRz0pB74HHWyo16OgICbL8TFRnyNpPrVt9nbSOHrJ3BQT5NxzXqARF9AC2b
N7aTleWb4HlfebIDoWKU8lDg8p6jv7FqJsy7p36frTL+nT1fshRI+WjY/EghlnP+iTe75RoSFSj9
e7bKW5eaDMWfADxqVuI46QthKTA22EKPZRx/r+1I4AE5Suv5wYjSpbUCf74dP3E17NtSK8Q75QEe
cr51NTWsZQZpji/QpdHz+uc0PEGocdRm7RNcq1hJDF6Am6lunMRmz4ZovZJMem+kebeLFyUxbCfH
IKMmeZ5GbPOb46Hxmz8uIFUFLv4VaKVgekc+HMR8U3+juiw+vvvDUSvzxEGfbWPy2sY5j2cK4THZ
OsBMaDV1uWJpKyXXdO6McuizW+urOuVAAcFWM2N6Tlnhk6AUb40fDru3bTPZOKQfD6Lb3X60e6g+
bY73iLpte+gKZDWP+W7hPndF/XKa+Y3pZ/KYFq8HzlJQj88MeKI6kLkarVh8Cnvc8QE+xkcs5OkJ
U6Rc6ZNaUSeQC9dqwe6u7Vj1zQCFoZbFKwo+rmjdj3KmQ9Y8hhXFyLa0C4uIfWg6sObfkzRdxIt0
YgXA
`pragma protect end_protected
