// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 15:05:45 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pNVVqlhnvsyeplILC/ytCYpouQ6gRTQp1DZNT4scfLJ64Q+F0QSdvAnfuvsdlrow
qrf/QcWi+icZjmNVI4hbu7ylSzjVWGXCYU4JSaFB0mu1VVyLvrjnOWLBBhABEfF3
bxksuCweWxGsYVFY8DFlpbAAd0PH+ydpiOw0ZaqI8oU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24512)
mxLsL01NAsBhsNGH6/v6/iibxPcChc/TgLc58XTw1K5Qu5OJ5VUn3z9vd9e62k9a
Y1MY1l0lla33PrxYaKTxLAhjkzGvEPungqOcriLrGRSNFXbOQD5XdapLr+B9oq8V
LgB946ENDyCjv+yPjNyove60iaMTvkV3QnzLX8Aoj+MY5Rm1HNIIHiiQUAAmD8XS
Zk8T8kl0v2JtnZ8Ey892p0/D0wocx9JsEiaFcultLeTQJEL2qsyj1WqcwSmqmj7g
naA6bEAbEsjjq7iw6HSfIAu3cZaHKup3yQn21CaCR6l0Q5xX53Q8oUwkVRD/Aazl
j6ZazMxaFzGoYz3stdwVVNCcc26oMVQjNCEi57bYT6fy2Plf7Ipvujtrm64APncB
9FepHZdpX48BtBiLNhZUrEEoYGgfxDD9gGBkVspJUvWM19ogT7AQyZBXZb7Q+vtQ
Z2PWImiU4MyV03rqn5GN1nKwNTwor+8Z+GFTQ7hE1s/X0dAutG02mjEJsxvC5MZQ
vEiruKU8daz2MlzsBjvjHM5a2c+/9X0bVUsYgJby4X84LceOVbJ2Q8ECqSoVZdBk
RgqkjqFX6AYd981cgYsKHS64VGxOztHdIXX/sOfLyMvYDCxBX5GeUbPHp7COGLL7
ddyWXuomkFa2bFltZ9dghcpVtpY+8Kntbu8S3+DlM7KnlQBurPrDz4MzoJy9cOHs
9r0Sj3xpxh5Ur+YTII7x1LXFZ8E/TgHsGZCwRvwwB9KLVZlP2bzB0kqRLXQ7r9RT
W1dhgJNNVsLFI443P74mhef302OkIL7SRi8KKNkjyj0TF2+FzoRNR1VqYsp1b6nP
Ftong+r+8ieii+wglmk0yqAFFh4gHtgi3UH5DbROR/wiq9WRkGKf7I20YWg9d0OU
uQ+w/QUStjuYo2ASz1FTqYdINHCknq+KBA/TA1eYmCrJ/xxDeoN/aKygNYH1LqOk
6BVRjRZ+mGNk4uiQ7lma2wjGsq3Gs3jYUy2uy5XnsO7GWnNCaqvS4brCeqKjA8FD
w0EkwUU7RCMbw/6LV5SZydcTRdLjydz3qsUMRvDxXZjRwQF1Es9oPCEf+vUlWzTJ
y+gbi+LvbzLzuJBTWgDrFDoMa3K3C17byiG2ulFLQ671R/jUXhzrmqR2Dr4/eMIC
YBuKzWVG3B8dYa0vvRhnEJhcQ5Sh8EMe1JvHPmig1jmOLJNf1sh7kGt0kRW3Gdko
PJU+yJStyQBboJ/cZnRwAiOCtEO65t0/6G7zJ1IZZ5a52GfrR7OMRxjKQJO5oEyu
HNUVBb2Z7qTjq+i67uf47qd47afMZaHu/Tm/pKzaQ5nYHZ2clfKCiclKxfi04X3a
pu3NaLTlA2HnWY2PY1kNv7eXrlpgCalQEnAWn1WpgAafSRYRgsx4uOUcAzThffLk
rIYOCdv097loxmd91cPYE0vpzkvoYJlXndYO76qr0OxWF/DpKnYcFhvY6mCWod8g
9Sos5Zxlt3FG3jN/9A/QpDOmDoqOQ8y7+vlEYu+njtoA+9aJg4VFY1zISvCG8xjn
ylP6LZz1vWFWPQvrcy14REMnBGKr/uzxyyxZnm+RmpKOAdhhm8qCXo678KHmUARe
sFjpJltOgsU8KINrCDC24D98NJjsHb6xLzqGjPot/GTfWLiHjrzMeBHQ4vRpDuOx
cQmsxRZEu+/tFYN9Op2TRLrCXTjzEvUW5HXYRkoXUn5em9D8hmV5v+iH24cOiH76
gwmtFDcSJL0PzDjCpm6iARGS0HwIAkIn0WNkA/AYLE3vKa6It8yk8DFEu3VJIGjQ
7NXXH+2rUSVaXfxx+8biULbEs0qn0BatB4OG8QSZMklBW0FPwtNDdQwFvaIAy+P0
y7EFnypT5Vc9qMQh1NRzqkOkqnz+tIUF4kui1abA0SKpmdaPqvGDd7IWJerkvLiX
CPyb5PjODsMdEiwWRHBLr7oRHT84FRFxoFduI2nqh9Ef6RSDl50WXfXkmv1OdA3t
wUU/RuXq2p0B6SGPaQ9u/AZB+3WX+gL07SKvW8x/kBtJvunjpVetLNLrNaUwffze
aXGvTigbC0DlRCLU5eQI/bV+wp0EM1z4N7175BEUQlX4diUWHrzDQRWAIfbJ1J4A
dVNN/nhMrGjjr+m6MI82C4CnDghZnq6VBlL2YhJxXFAAgn7Tpk3Nrev3xluCpH/D
hpeemA0x0sidA8iRz5B+GbWpZZFjfaQqlwImN+RZcvpmlLRet9gep5uPA15YkwQj
39A8mJba57F0/fuPzLB3Ax96sM8yRyXEHOnnHkfhDuHTLMyX1QiLcDoJNe6fTmpx
2ROC4Q25dDtRVcf5TY8L/qia41HcWxpZPt26fmlSJs4+C9s2rIqNAP+AjRZ7oHkL
xuLPTwjGRNPQGDGIx+SE4HEwwOl6XXTBwve7xT0RBNciMFBHF9B3fhak5lFg+IvR
05jd10M/sq3pwQxsaIAnMzSimUcPjCbYQuSPTFCrIhoCfyjU7PshDff0SlZ2l07O
U+gNWi7F1C+PRCzdAsQGqmodBCN9QgclPoXCj+KS8x/5Qn/8YJtLbD1rVoxeTqq5
fq0dO3YUIBdO4niz6MaNNYfJh6KRSB9iVnycEQg75bFKZFXyHclEPtseErUH6zVs
0F4By3VJnKfzkofn3k+8CZd44xnKO/TEJmO6/yBZHD7y6kpjjZOnoR4zYjlYzq9E
PBIQp/udMmByH2CatRw2eT+hh0UHQjsZi5ekHIhZ9lhCOjVKGKdU464mLRsdeLYL
V2HhKPHgy0wcjhD3tK7y9VtRzYPPciSXFFMHP/0O/ANoKSw2CdKmp5fjTNhAN0Yl
H9mpwRIKCayEwZRvEGhQtQmFT/hJZN6YBFGCnfvPuQ1cRkiJnMGr8bFa1WCRNyfM
KDMK0G6GDuOSND2T57qPIyd3O2C5QWzyxZY62qZcrfo0e20hpnrRe4Vwcgsrl/W8
OnbnPMh/Ch6PeWfNl7GO/zSILN3+7ZzZ74scF2RkxrnrPXoVsk4KBc+OUzl4mLdE
sHHu8ns/3ys8UfRusIyU0xkVByCvUfp/Y8vBPBDz2rQsZbzU0mouWH6IK97tJ/DM
idN0k0lF64GV+NhB+dh6HnOb2x8vqLgapa2GfAxItdLzNyCxuyisXy/ocdbD7Y3A
lBWG5tFH6d8a7j0ngI3XMY0EO0RG4VCEZcAt2Tql2L/Que6olewZfB0RNydBDgHB
rsxrhL8Nsg9dcgY17R8D6r2/GbPqrN7QF/hmOzk+mapl+D0o6jbmmEGmQEWJerOm
P4b/MYUqQ1PuJGZcAqAHxILxnQvf/kkxGORmJtRU5VTEB/mQLPftYXioKww8gs5Y
y83cVNy/0uuNlaI5SxCURiEsVW4VmYfEP5Twl3+v9mr1He2x6PwPVC4DdogizSsG
v6yMLAH8R215FVY4mF5346JUs/3tl0+GiDpf1EwD8DEdJ9s8VZQHPU/eLifISRjg
MiSjpBohuwK8GTQUtiWkfW7h9Dlou5Ga61yYdSZNb2yQiex0sQS+Lk/MB0SknAGK
TLlPDvt7ZJMqbqN1XIf2AghNCQ++uJaLWVQBgexJ0yscFPJTFubCO5kfzMrI6FH6
++nBamuAX4tsNmtnX9WZHypxIrslvU2zePKGhQ6vtFK/AjHSTCdMDGJMz+x+bmLr
VT+tGWKVv55yNUsFzE6WBEqd0E/Y1r+o9T06aYLR0FxLnFRiETGkLF4NcI8WMYjC
kQkGXr+C/cHXasFjspNff3g1jFHWHp6UGaNo09VmikvfncVNSlSlPwIt9cKg9MCA
mbEUFsO0zpaMoSa3CzZt50ZX9bcOoBDmd+Y6++M6CWKCxttp52DpAdOcRG3aajpm
gPszD+M2u6pvC12OYUNL57W5xZCLSrzPFn+UFfoWpeTCNnc2PoWZ9n6MxvocJT9M
IafpALRu7SN+k1oAkIPIRSLDBzkiynxIPFheu7679ZEH6R31T2wU3QPyM8/UFGbm
W9snkdp4QWLedeDrYT6CdQBSrdvJBM77fFEaEfa1gu2rhYAL2Sz2n6n6YiaDS7qs
qk1ZM5UHhWCEZ1+zszfYzl6ADKPnkhBIPRb7RlFM7YRhgXMTzrBSLDnIKmNrNxTz
dXB1R4xYycDQhegP7Mm2ll8lbzi+C/uvSe3EwxCBmofr30xjvEJmrRGp27QrdPXB
CMDZnT6vxHImLzSyPe1KPYUxDiLPZ//mPyzGA20UFEeyUcWvACUlhCJ2OOyPpoWP
PVMEjUvQGqVeUfaTsniim5nb4UGc9aAcLiyren/gr7j75Xe1YcfFUfGpKgGKWTfT
y1AUddeQ9OmdeDig+MlhjUlwygFMEbeRBjbBWTTly7sbapgdA4aqgIkgaZquEw3Y
AlsFmOSnOF5o5FbshKiz+B1uTJTX/qoY0ni+j3z0Z4YvsH+CgVpfrm76KhJQIJ7+
QmHzQQUfiED2k8Xw+ufDHvjUXEuikQfC+sNSXwpslq9Au07wYNt1ceVfAbQsv/hy
ruEmlVOQ6nq8q7jBsnA8GguuTVQ68I1EPXm0dDO3iFGREeqJrhXqoHKP6ju9PVFA
86jzKqmyxwNqm2rXWXI3ichNm937zbV6VIpLqHIFmq3F7VBGwBAMkf1LRY/WURpN
ZJ4AB+5pbeyY8KI4AwECRT0UdLgHMLYkFNzDYh469RvMvGiaoRnUsvnyFEjT+z3N
JQlfLquvlo69tP1twvMChiBYeFEVDEw4+vGxL2HBoFKQ4NP8fs1suAVk+vf9NpFz
zmAnDsrZdOUyqXvCZzspUnnKEnkytXFDjj8cg/2Uugcht5Bt0D7KtocTuBeF5EbY
e6tp05fngPPqSYjmolMLJ9CXglPxNgLfkQTBoVK5D0fbHMKwBJ2DYD/gZDeDP0xN
XGxqj9bZCDEkNBm29bRXMA7uWDCaXqxnfzcCTrKXuoZZfVPUxJ5ueJXD+esK+rty
96K+0Cns1Zn/VZvTsKovV18N0hGzDJbVajGq5fxNYmWwCGsKTEHm+2WeFqPzFJSY
ExFJXaKr4gzEEnTqDmVT7q+w4f6zLOkFF3hS4eCFB2LCjceg5Gp97zozF1BfwDvQ
5/cAQLAbIPvDXAAGWFu/q/UwtJTzueQlAhAeokpfaGbzx0XdRZNR/P3vCy7CTQz+
Z/lX3JohAYQdpKcXKat5yQbw6VqvgJk2GyFpPJa+MDkVpvL6t5igW+wQSzBojJZ7
So3RNR/XgTnxQ4MeenFoXti4RZt3rJJQxiSZnckeXGpqOa7He8PHwSz2PkEzhkk+
dsNQyRzMEgA37f9a9t2lEOepmnVurlJDYIR1OuXiNoz01cmC5DmF3S+5rCAQZtLY
6JuTWCG3RsTtrOMv8r4arbcGCfdnW1+fasWiG1mIzVs6bW1hA5XLK9henDK7c8Bw
aVI9OE7jz3KOiWWmI4gQZP2Fv6Pu1mw7yXH8NZiVgVRFcXtoA12Fp0sXco2Us0hY
VkmaW/9o3P/qRUBGPoiIwd8pv3tAW52SvUx2HFhv1aaIloVnXvl8mHnwppiShgYX
Qk7zkCcbyd1oHZ26uF+KEUe2A2b888X72AQGLlJ5TxmRfara6ixnekXvltVRzc6d
40RFkXAA6Z7fNcUa4xtLBcGlt70aWxAYMJ05Sriwd4uCavrwJHk856r/RYFwY67z
gf3E6CL+wle1xjA7XHx73IeobnEnXcXjE/qUzZM9Zcl/3zHiTaYHFyUpqZ+O6yA7
TmoupTw8U4hhpl/AoY4TR41FnFM4Z0zlfaeLY/fgliBoprvHRxVAzJKQ46P2XfV8
GPttuZt7HUA7L1XS2ZYv0nKgt0nTuzqogbw6D27YqDTSrGIMlIEIE+xYHkLtg4qe
7yj9zoKeOEwLK0Yc9J3UYD5JSA58rwqN6Gh6SzU7RkrMDq47CbV6C5F2CqCA201o
g+KKpGOEtZPqKE5/rDaPrRgS3PRi58xEibWWjAnnGQXCh63bR8xAjKybunnulFNh
gkIbWaUevpezP/fku9wz/6nR3qQHKy/wrtq509vLEVKs5mNnL3F/JSZ5bI4miqbn
eV11PTjuemaPtBXUB6/oQ9sr5VHjW3jfeVS0/SVKkb0B01k5D52scE80sGM0EhhB
Cq/AUrHitT1oLEA3oJOaNRYcyuhVsT/6KHLSK37IpdJxhiK66n52LrMJFwfzpqmS
n+RZduY1jtt78cUu4gejFNGQTP9pp7OB515nDS7I7SGODNPYeD4TkWY38hoOEPqT
MQoEbjZ9CERyRDLLHood18DDbKcmiGQLo9lquxdcg3D5PrtbbPnIglXOd+51D4+X
pSyR9R4X8FHRAfZHLyTosTyP1MYX5ZZ3bioFM2kdJ/ggFHHw2lP1pDmP5A0S3xLe
xvu9sFPtHZkaDyIeM7dwtIRBzd2nBFJDBbyHPfpbmVz1HaAQGyGJIkYqSeLGge3e
d4lrSe80CqCF9yBsDH1g3ud9geg7dksPliCOPQVN3GsWPqnlIWCz1ImciAte3Ek+
wzUrnZiZR40ZzuwOcT8h0FQVg0HLJggzDVRaLMFZSvG/ov1lxJBKbpKkp9y1Hyna
RlZY1IC6p4qJq0MfHYoXOjYmoCuIkqJnTOa698ypB6BvnqxELYDkghWz1FKX0fdu
+t3fR3L3dkLbePah3lXMtlBJgcJm2SBGqQN3j39s4qC6UHOlHwS/r/ZOaFgfULyh
YxALAzd0t5UTqzbv1IWWviZk4XedJXCNn6jNeamshV1MwJLDSfamwASJGJLla5dd
WmEi5d3woSLFQmQQdezdVDrtqgsz/c9pNbIFLnA3zIvrwM9nswDz6dAwt6zc9w0g
2JQ6f1Ezrod4UdV2UkTwiR2pver+w10ZAr0ul2EN39oUUUj6JlPgnqAZsxowkUUS
GuoK1ffipNbneEY38UI1lpOEtNC4NFD6LlX6txUelfbD2wdLMlY5qzI4UTNlN6Qb
CS8qej6tBgK51d4aE19YpWE4xcwJPSW88RRDuD6nQ3+wZhYj7mSqWBqmt+I1L+sw
hAKT9blHeZQQPsJj2MeJhYlIvb4x5RugpWhDHDoWXYNVuKCxcvawR4y7COAYSuDC
tYHbdzhqkQ0/ctGp1ziduVoKQH3Zfzvwps82CXZ5i6Y55ET+Xck9Zo3YQ5eEEtuB
snZvMe+OoiUf/uwE+TWPakT9lmA4tEYWvv8nx9lQSXfVkVB4tSv7jRqQ+r6KZbP6
Vy5id6wOBCGEYoNOgJ30LNamlohdKvi7RE8vuUhnNBgYLqdc1uTcVcxuej64HAG1
2MKCRm7MBuI2sLzjHnZQdhqkDjPE+uMqwGzAGClr3YQ2ol/u3btl4RKVsPN0HZdG
JESDS2n+sPm7+TUpSs0inrvyC7zjRHLhyequUfG3pwpPpytJoPkvX1kcHriheLaT
FAw0lkHL144CXAS1QxEtuXsG2tBw3YjbYaaAmGla9RtCsWf7NdA7JTKADFAgm6vs
VgcrjvzmZBAWteYNPU0qYmKaryZ9/Y8uHzPAdct4rjFx9edxjdG0hbOwAsYkj41O
ahHjbmWxl+khRJ0MB8Xkgnu8A6mnpQGi0PO0eZRTgK1eNeFmC12v6dKfUshLYtUt
WU11VTZ0V36IZlTpKyzgGCuln+JtDmjgPACA6hiALQCZa7Ju4D67uqw3I/Wm8KYZ
qDjc7xgoGm9r1MWjmeIXWOFbr6jPNvlK+ZCcBS5Gv4Blv0/NbTEk7eNrJeuDqVRY
OFMVZ8zpZRbAsPppS8L8sH6pbujfvdhzxnFdOKDw3j1hVuTrZ11eI7077BvfYOHk
7yjjdkrnaxv4COOw9KD6INETESriywLuqzterm8wraFUtnn1ZZP/YWSswElTnUJK
vdGSIQ5wFJfctrWPFyz11gS6w6Z8hMvvFKGlRW1FEIvn7anHC3Wpra/B150I7pJU
dLgZSmLaJ6Z3XndZCaO2YZDJBTZt3T01/4JKlGoDWPbKcXZkTjbnAeWZEHK2PuFp
LQMSW8GUzbJDQCGircCzntiKU/Tjivj+7YIFtJiNkR39zxKiWBCkAQakluxp2prD
EeyWc1CM5NGsgqxT6cZ8UFUUkB0tU5Mkah4osscFoMBti/swpLUFGxn9sbMjJ5Gu
WlbF1AAxqI7USOpFD2tL63OMkSFpESseUteIrXK9A6/84yj1Mt9nLoeqZIF8scvu
6rvmRoTZCNccZQ19JUPJ0VQ1qBMO9xSabTCIzNgbx601++g2QNVrrp2syt3r7d4d
Vxycy78FuGGEPeDSF+64iGu/WZdSo2tOWk2fH962MJ+Hkj9Sui8C8exHtRoWtu19
e8b0Kx85SrvdyC1zy0tDyAyjzTmUesVs1H1xDkkeyaFT7lxlXq90W4w9ZS4POV14
bMuGk1QN+soe1fxT1ryb4EF4YiFDey5TSTjc83ZpT02OVpVw4K2F8VkVFQOy5otS
iT/hpJEf5F1CZ7yBYvb2zyGveo7K1lxtgLCX+ALsB38yHwxlgBoBkSScVsKA3+Vy
z/25uJ5KsJeONd11QH58TiE0WOZqCZSYgfU8BNbYkuNwlGnYRj9dKPJVshnCwA4N
gnn2zXZki64l/6U9dpQU6imLWmrr8ZRA53Qdw/py0d9JjDHX1IqSy/+hhW9VTPCS
9DqcWpr4O/ke0qEkqGxZkHSgd4+WQAuGz60qHWUfxi7F6Qot2EsUxxEo6J36xrvk
LVXk28MG9ivaznBGVWvSfv1FnyhT2l1M5LxnadanFHXgmy5IZYOo570KpkK2gU4H
+sdjIWPidMT0Vlht3FggGTdCy0sDMsZ9zJ2sW55Eloo2uX4zuCYvH0Unn6CSewOB
OTXBZ61xvcJCSo+0MJC8nytAxi7qb4Ba2caU9ElMEy6huAKtvF6vSvj+74HSjZ2c
V7ksKFljbiUk6iZmB1gT0sIYTD9WWGk7tA0qJm9T+VBcGk2lMMjlEgH3hiTjGbuc
A4AM4tumYK+WV9IrwB2fJ9CPMXhlAEqibSCm7NYPsCf+csHkNkyAS2+fhLx+3nOS
XYbABDDZqDDJTY3knQYH7VnySHbEPOM3fR3CmVQG421xSbA+9TB42vQsKMalQ5GU
OXrpKkH2ivmfylmSGFoLXRiXFIHNnOpENURWNY0PZl162cRY9Z6R4WkmQh7wznnD
Scc115+OI+wgBk7SUN92R1jMEJy8QgPGPHjJoAvec8L5eLrRJuoFBpN4prmwkhRD
w8XOjj7bwCqD7qVX/LceyZ3bYyGgEtO1G2daMGEyU/vTfUr9apctzHZct2wLhAJv
fMs5ROHww0Znmr1zgOYR8vMUaeQ6IJdAgrU9OmotYZDUm3vZx6eBhyYwo4d2nwqJ
Ztu/EaP0uKHoe4+vS8oq29gi6hejQJXl2/6aCRo8q5UlQ5lO0387z000CO/1rV1L
FiCXekH9Fo1AAHMTJaKA/rIgRv2lhXBg5RxrZZuj1ww9sUE2Xdvhw2OCnQxUWvk6
vbpuzAnUelhWWvglMmGMOJGdWUrbPn83pLnS8mKyPjZhiswgTttZV8b0FHRiiaIB
bhF676EFpniMFFyAbq8me/A5Hg/4CbcXYeN6/tUD5f0299ieGR3qZctXenfkygCw
qp6caocn8QpdOyFcewKNnpbBeqCH8uOe0zJL10SwEw62QkiWkAXeLHiq7QMqx44D
GQPawlrdpg53nZ5EnTBAJNI3ULQXDG/017D4EC4hFyxqOU8yEEyHKJl6xnJYcoFS
W8Hhd6ttEcFC05j3jkhydATP2FERHj/4rKJTA3Ix65P0gcVdODbkDvaIObU9XXPq
PAtQPjMnNkt5rWQMK6mLJrQPXg9g53ENgF+mdddtPyp3a3tI2T1pdN3zTARijUbh
XyxnIrS+E0GMzGjQWgdjxzx8k+l4R5AWGeT85IgTqAaFeE6MloiQBtD9+RTQzaqR
Bn7B3vOCoHkbvApWNFF9/uR5F4QFhoyU/usmANsijTEvPcpBIb/FRnJ0rNCJv3B7
qoL8ok5z0YHFnh9sgSPHVvb+nXV52Fo/SGUg1ZyuO0sPr8Gvf53IpkxE5kXjb3d2
/MJHdMBJwFucrdZaykt1i2LRySFY7CuCT9iv8FYgvdeaSoEeNHmvG7LbM+5sc9r0
4GkrdsWerf7lXw4EdQUem8M2x18NgACBAfSd6YEHpoW+uZTF5SREQybroqqMhYT9
tyVRzJm3tBB/EggIx2NUIYIiOgbWGCNOh0HPxYIfwhxfPF331VUDO4enK+2U6+s4
nz/XMwEiBJKSw9MbJlqYRZKVyLWAbhjn0m9qONRQFV0A/TDw4xO+3nQlmIwm9RQy
2TLisjkwcL2oDF/trHgyG/EjKFWkbRrKMX17T4yxh8i4zu88V5+ZF/5PS9ugrVvC
GL2uC5fHGnZft7/G+KldqE13Sae4+KWxcIlNO7Qh0z/Pg6Ipyv6AoVvtXGzX7Ak9
naM9tleYKh0IjeBXs0bUzdYimJAy6mLF6NxShmV5ce4svOQfmTmdRcJdaBBKQEYE
rVRKh88NzUWPoWiuiGk2LPC1QYcc4h5cfnH6big+jdvpY3iUhYiCUg5fiEJwsYpd
3DZ6KbbeYAf9fiA14BC5YdVUl4Wm9SMey+YEfnY/ngcqIyrYCRZcUy9Hk7SMS+zy
FUx/REMDg/R7bKsZnjw2xk0AfuLCm1CTx16YKU4lecf49p+Yavh8MgIAlGSOI3nX
KdhuQOb/E6blVDmvCKLdp85xk6Q+AeFTbN45iXOeAbjjEYOUTFIeGOXKSpNhsxLU
fub9dK0ZFA2UnYyyQv2fRXfAaoa3bzPh043em+WZB9Qa489HyKALhXs20YhmK7cs
bQ3bPAp35NsXlu4JlokoWeX2ioc1fS8D6jEVWjqgsdD5VjNGKsrhPOFJCygVkGGK
3uBVXfMlz8RRlb0+pdSk01ziTP3eeTvTGugDyGdhnpxmyh9w8GeqbztF7nfz64XV
PBt5xpCvJeYxsJYhP4zUXTgYtRHTBMIY55xAUhUrwcmbOEXztLzE+aGbOEZQ6VG5
mtUs4il2KofjrCOQ3T+FUKvVaea1ii3VzDBhtQO4UK5ssOva/kFMTLZqplRu1H2v
6y/Luws5vOuGgkNuJPO6oTozoW6jtRXwZM93GMqmUrcZntyrfVecQi4ejzALPbSG
l+ABhgcUQ5W/w0+m3Zk7KsZZTMe12aIbYEAdXHRB4PXKIE6JEOErbbw2BKD1G94t
UEzJbHUSJoTNomKAFk9rzolgrYulforgjCa7Xg/J0A3wyW3mqChVby35Hws7IlHG
FhJbb/1ti+Ts+wRQDnRJZH+m1xHcFbe/ecWaL0+IxZxFBD598ppH1Mn3CrTQjaOf
7OTYILvWd7Vw4vgvBoMHNjxAs6Opo+NO2Kiz38n/8+HGngn7/UsZqgts8C6m7vQS
I7xMc+4dsPXX0tHxjyCAi4kx04Opi+6FUpNdFDApPNgbc/aoASDcZh9y8WAYcm9d
0lnlv62KarWODIkVFlJHwXwwARu+/AO2mArrodTJmKEdSwkrfleLSvwDBmge6M5D
5tXvQHIsdMi2fYO4cyUdnpYzgj8xzjPnIkuAnXkSuJ8+XZ83EyozACUeuWukE4EI
mpkyOMzzGM2CRLIR5CniTqO42YLesQ6n5emVHWMf0CDC8z9Ayl0KRc3JIKHKMmaM
d69JWGtHMQDwisAEwFF2G0y8Z5rbX3KlWCfirZ95gje8hFEh1zRIvcwJ5X2JzY6D
m6Dm9jYacmFOXUjWvEbNzJtM9k6XkjxivopII33QTqZFc8HY0aHZVOJM9fOzQ4P3
qcEEibbBFsI6b5yLiHzrbIJD18dij0nQ3CkWI/b6mIOx9WlFmjo9Nyw48eh0ouEI
Kvw4YQhy1QwFMdgE0tnA1LQFdAbhNLACzbw5Xd9HvjHbx94AWf9EBRewsrIqB9q4
luicszbb1TqIBTkxJWk4KgNuqchCqwAi7cukOkgz7t50FGET6GLjMkUetMzdDeYU
UTimLKb5Immz9sXxAC4OUyT1AUXVKEkPMyyxznnZmbDLEczR7AOBPD/yCfcxljh/
pYI3DVzZNbXQ8MaunmfVamXTjZQ+9p4jtmqdkEjAP4k7h0FUkzB5eRpXUmt7COVi
/Q2mVFfNlmfjiWtfdHAzH0N9w9fPl6iZjgQIexkwNvi3zcNEqz6W26uYqYVsY1Ol
JvrdjD6ET901FIFFARFqAIYWFILvlyfEuRBhLLYA3ssxCNIdSeDarUuF4zkmVZ5/
olKpeVrrkVUjZXoLME5lVwuWv7Uc7/2cdojNq+Mo9GLEVzGmlrjKXNaoj8Sapipc
31CChEep376igWa2oQ9wz3SKSPPjBS7Nld4+ARRdBbaj47jz/vMDq18IOInsYG+T
eRSvNmhgQqpXlbvdNb6Cx/G7KF8BzPwmlCi0ifeGkqX+GcFRa4T1kZtgm8qfnVf0
aLCAtr6KquicjNuAJ/6c1azB/PRiDoU+CtPAporac30DzC9C7YQFRzmn4TwKm7UL
j76zksHb0NJPvEN3A0+x/qvEH9fPsNPAUP7pTwA+SH3bqV+sezHFtywjP8CKFgoZ
uhuhER1CUmWPlXILdUO2cZBC8aro95NgzEzfesUDowofE14MvuN7ZzVIMnYOFR1E
T67ID920HD4XAk7Ex1E9UTtCzhbxPYjjQeaokSB6ZXyTJSplgRGKYr4RpexcQVzH
IPdxSFwTYHsi6w6Scystb8iv90kB7AI2USIO87z86xELuyF+X9o4drdJSG0DzoMd
OTNiXJVLVQ2sKXuiFziYNHi3PzGBzg+0HbWMN9yZq/GOqPEoJB9vEjcLp4e+wQRy
CpJdtoKaT6vFsJXMbWxpf4qMcqCj0ZY5s3PxQ0GkzQVovQ/9niKJEnORL0eYK+gx
Y6/z9aZffaIFWKOCJOzEUNIj6LuDCXztJXTw53ROBKP7rNXa1U7UUv8J48/z+G7I
s2QROdUioqPem6KkXDDZDL22KZETiRyT8L3GwXmNmUDpoIvWD2RuyIDKuEyv04ZX
7TuhUETwYeBTBTOdvZFCUN2CXb2B8vFkAabIKh57szay0sAutRKWd4LkwKKES520
TSn+d3rYO66reCv4UWQLFs8B0YIFUilVFr3zmuOLV6XXznqeh8E8+PgKc/XCoo9Y
j+999dfpfopC7gQBoDoOwjY12/Objy6RTOv+p5BauPitjO+4SOOC2mjbdn6sdNbB
tPGaaE/coRaoy1SKX18bn77AZF1DXr6+NpPp1Oa3Sem3XIs6HFLUYX9pPNag0nhb
+X6/D3w3cWgJ2OgMMT6LHIN15qRBylbsY9AkgSfgJh6A5CFWC+jyspJuRyQvVhIm
q/lmuYwtLHG3MGxszhVdz6YR3TYfdzDqV3S/s+nITg8mvl8Ix7OkFlfLW9vEZpbT
N8BZH2bP0P0QO4pCkvS2oeOMiBXpExraYvdtv5e2qrXQFfH0b+CdIYPNPy4mpohg
EjRXAZk4gH59nF8waKlojbjEmcLUINKEuRAqonZ25efFn4yuqXzS0Qrr7Q6KztEn
vpXCCjRprG9Hc/FqIBhURJyqtxv87O9wR4Ao6Q0OH/RLZlmaxHPvAkKCLomJvHPn
5Yk6Utooke7hK7znF+zI9CREGvrOkpudk6pBZy9Hy1B0LDGvUvzRdB9lwUJc4I50
GwQAlkyKwh8KsHdd68iuHUnuPjvvCDeR7Id/OgMwOPRLaxKtvaa4JPhlYq+GdHWg
SU+vKg44P4bZNFKAz51Yhhg+GNXluLbuuI0Hf1vkzTQ7H7Ivh8WYnlgx4h8sZPDC
IBjAyVJJlrLV34IJLH3MICTCLyDoNchu6FrCnTOVnZ3jrGsC6UZj6PpDZYUiVG+5
2xb9rd9p3H7hFJ5IUpWe16DO0+oG5vQ/avk9l7kjlKqb9M6sQpQKO77tdAavlk/z
6FTSfd5n+BrTrnbeTOU51bFiY8Kr1BOVImlaSad+/Cqye8Qp71OG0u1HX3ZEq6ol
e9ZItV/q49/1b+xq4jhH+X0JysNB7JQzQKHTBqhO62421H915tuvHAuUSquhZQ5M
dBfZUIc5pzvrl46EhRwreeVzumvTFJug6OVuI6cHwDNloLV79U70oItK4+Fd3yQH
0sDNNI2NmrIyofYsPe578GfFmTMgjSkgVUq3UEiCnbT+59Pr5ElwFFj7yQlDJvyd
gJrSKg2e4Te7yKCA3xk80XkHd0NiuVI/AkUIicczQvevafscT6SFPe0ylk2QrWtW
UUgm9zmfB4CM9yhCetJfV0LYjB6Uud7GMzPm6F+S1zwgqoHDqEuRurRljLaRvHf9
q+xWQhXV+BUr0UHSWFLD87Ivpsd2s50OARmAoysrS20t6+UwQAxESAJcRsicfZc4
hCh+17gdOV8KISKkO6eVXOcGB7vP5cVq4+PufuUD3lme1zDTolg5zYIiLLju1C9o
4Yj40ajPr73iKkyroKAKM7jMbju0AEQ6zLtHDslzz95f573Eb2aoDoiYW5fbl8+y
NtgsYs2rzeVJfUuxEQIZR7UB5LU3zMssWt3HBui9JKlVGar2QtL4WbI9ZkkI8C4A
Gly26YuK20U/Zcl4YWhlqAyx+Upcol3dx3WJfzBTcpGdER6p8wZilHFj4FURF4b4
iLB9+WrAM6XU7q7z+ZdWu/DnuQrTgc4qeD32fdS1AwbwJ3hjc1WUABa1nwTGciKx
kbsE4S3oKcONVo2KBfB6c9IDbf/FxkGR70iW0rhUdclzMk7gHL866Fu+kkPg7/Us
4yo88Mxi+bBRE3qqAuR9jWNMZ1smNz72oQADS+AlcoI0FIuLcf4iKvZ/fNYQQk8A
20aKXpVlrxz6e5XRhKvIDdjsLw56OGz6qrYzQIal+HFpE0hfDkjD40k5RAnAiNNb
NGLO1QEpD9X1g0eJjCVlU9wMaH5E/K0VG9A0BK+LuQ3L8OX86/WZIP10+5PcwGSx
pc8DCYa5Q9csxm388wn+PyBa/UPxzYy7JYD7LvwuNdO8Yiq94b749K4lBQ78RWhb
+U3WpWn4ElobJglcnqS4ebWU5Umpm5KGIYuILlon8b18N8Dn9osQaxaVNPa+nBAd
vB4r0x4PG2A4Gc7hnKYg9ukn+6Bdht3lEBvOjODIror3XxwogJmNdOulImS1qTlD
qodZBuJK40O1G9fPBAwbgS0lYW5Q4NMIiiuJU8qMoQWY0vwGKbJXtMxZPK/c6lIm
X4BpZmW0yT9z3OtVVMTluDndDhWZOkNb7ku1QNkgq/vqVaC3DnuGP6F5VFICfuel
n5nbQfcG6mQvb2/IuFmf6fhkfeFnLnPONlR3cq9LI8JGwEsjxUg4q9odcSPtu8dC
eR7elejIW7nUSORJy9qjlqfq43KXOBH0H1QwoV/JmN+mL3jGyaN7LQJ2BGm41QAs
IMbMtGZif4Y2M9oS0z0cV+KMdZrxtCAjOR7qqW6d7OIseejIWz15yyDtrN8BUW/J
bq51eTYYt5YgXZeEEwbUgotdkanZTrB1ctW+pyWaaaGK12Lb2O82HSBuwQgGPNII
nxfgLoZgcJqdqWm4Ipbg+cQQNh+heAIwp/kBbrnSuxuDKtSksOuHNq1FWndk6F6A
0yJouNSxtJk9MJhT2V53YmRbYMkDU4oe2PnA3KTACKZB7nV192IGUvi0W1E14NfX
Ss7zeGBxpljQ5M/qpFZCmRt2Hnk6LZQI0UGJWHsBevcC10+iIc6Y1/uC6/uEefkA
YeacWygK5lLMXDA8d/0h9Tc3KnMPaAJjlBLL2/aIowniZ6cz5iNkHFmtkrQk5KDL
+gHYcbqUzvIdEM5lOj2rtZnLIuzY9A1tpI400Lz0vCrhF9G3Aqg5YosG3ro1+sgQ
VjK3mcq4uYmq+BreIpSYmUvlyibOLjghavh7iAUwKFnThFrvOpuPH65vG0hVy0ik
skivj1peVHD0LLZ5igk8AM4CwYQH0ILsw8No6k9C4c25iPimFqcJ/+O7ES9lkwfW
Go6MZC2Fho7G5dqtK1ULWy497tuZ9bj5bedYsNLbSUTLLvVkC5DstTdkx+EAZY+4
v+kERK6Tfn/sJ5Nh3Nf5cuykIhBnRfn2I/Jqvza1PbajxrjLVLLaJzUKSKT9AQBI
aNGI6zSHsbvfCo4hQtwOsdnNPHm/lNgr3Mnm9RkrEt39ffoDQU/lV4bdLdCLn07I
HgbYl9IntCrYHIX0/o6iaI+w5+AkO04lWi1gg1o45xb36k49Sh8p6g5vtzmO6/hv
BKB6nO4bXLkbCtca1Rb8Aj3HEJPo90bLsXjJdC3ZMmXUKZC9Vrb2knQSKJYx0tWw
+VgREt3RpwhQhuYFEanYyUFiP3uWKcgQS0jvr7ggdCuoa9zcW1bz7aZJ9lXHoaaz
8vaRRKlbbD5l7HzTQuZtQ8sBga59NkuCe3CWt0boBMN74uUawfhuiaVG6TmdQDBr
O2lUapzpU/QN4YZduWI+C3ikChJDmouBIt2+3y2X3Eh6y/vRwaUatntAlfLkQsK6
4Tgn+A2MLVshYKmEGa0ddDK3+maQeyfjEz1AMrmMJO7EQUl2INcEm5F5s9wG5c/U
1X+qFHmH61WIu3ut29AmXGBotfJxtqe7Bc4w9cXJd7hoWfE0foPiZkjpU2bS/ZpU
APimQOyPjjHvuhlaOfhe/6zsc2FJ//jpXzkYzIhsDznSAbGUFCCWQWeYClKGc+lO
AauE5O7r+y0XTI0hrCDQ9Qt1Kl5dbJqWLiNwIe2DRp9hLjyZAwlnCs7Pl2t4qeQD
cIUUuJV6sMRbtaeGj6Cya1BcmPSdCgxJGICNFPeug4i76mcaNtRPQtU/lJnO5Gu1
8AiopXZe5Eph5twRJJneMvImtAcYYmILMM4fOuffATUyS7Om7B3bttfedSjPy9fD
eQGBbgzha733ChWp8Cqqqp6oNoC27XO05gVzYDBxulzUHukGwaBkUt2lgO2q7cbH
9ueQfpeXQghYDENXv0zw2tG2oF0rJlwoWjskkGxLvu6gixf0ki0swzPlfn4l4BzJ
DDPlXbjia2c7+Z+wa3v9sQKWe3Oh/yYljMpewm1sA31ezl7rzf7+SxBeMdXEbw1o
HD3sNZ50TLZi+HavNb8XxCIgMxZ8dGkfK+r6ewPZUF/ndBuwrapftLVzaF30IHqD
qMAE7PhXkD3DRWVzW+agPb9dUlT9Nkf3+LrbXVquMvPEvfkkWklMRjNSqMvlcsfS
EKRQpvVQBO8Id+5p6bebYMrQ+yLKTquZcxKpqRVephndcdAgTfTXJyCmJJh4PvD2
5dxvIpXYVTRqPsGZEmqBwKWQu6sDu4gsVNdBi+hy42ScmSoXHtyb7ynxHEHlAenA
2MtffEKBqYW+jEZR0Tjo+GhICPZHbtnaaSHIo10HQ5jdoMgygnJ9CvAvoNFl/fTa
Rhxb77b3GQlX9FSnC3+cPr6g/DOsTt7OuhERQtuhrnVYlmsSBAhc1iwL29FXUbTW
8X2aOWgLowlCwC1A+J3RWiSAks31g0FnqJaz62/odlJAkaitoDk1BKZpseDDERJZ
gvav1hPqVavmvnqt9nEUTO5qvcbuhxr2g6A7UMYEGhPGXXH+gOcdHL2uBNhYYY/i
1UjCO4doLHyG5hnOAvOE56QrFiQADKY9/DVXrQoXF593ybBTN37TyjfnfwyKpq2d
MLpyGghp86kD3Xb/wejGcTzUfUPEPOZG8G9Lg2oXzO63xFZav2XJPOGZ6B8MeJ98
FkECsOje46kLogETem2lM71AwWQHl8YXPhCZOs9QOTq/NER+WTfyFmTgk4yZ9BCX
x7JjMkB+c+G0vIcXh2CNLoru0fdpGRF/6ToZMt8RK7X7NyF+0XVPnNCoj/+LDJ40
K1l9mISd1hfPRhQ9s0qzZtGuTjeklgEId5pu+36FhbepprCW4Ux6CPlI1qWoJMMQ
Cf3ItyW1UWMRFT9ivLzrBZPFwe73QjceM0LBLihvII70FYYn0c28HltM46/X8IVd
aXcqUwXKN2anvhgRpZ5OWzRt5BLgsvU0yVqayd2EC5skHXZcpsg4c94GJoQhkvax
mIU81T0MnQsT7FQ6ulMjnXe2qqPIdeYjelXAzx42vHhm/QLPLsbv6zYC8ea8c7bq
70EPlXo298mgPeR+db40gSKTkprReXNssYx8jt0K0OYceKok7o5Bj5llNA59vLVl
eRUTHvkfFtOD8scBGvVNAvFUzUNN8joJ/lPVBuOROTW5JS6O2bLLyJOjuO3dkIeF
l/ho2kT2abvo6vFAAFAFopT+ww6zUFo4DacRpNUWAQzMbzvK7Rdo610dhYmNBgHR
Eeg/Cn1GjjLrB+idwBpsEMEoN6t7cPdhB7w5HkX68xF7JrCIULExcFV2kzZ/ye2V
G1and5wrRgKkF2l0zOFpPyyls2bODPPNxq88NQlX8qLCwsBvtfYpy3HvOf7sXNBr
bLZxyDp32x5Z0r3Am/huvSeI3VPIsdqQ5HfRtFFRKICBET+5EOTe87FdNuBsKFHT
MJhWPYahhlsbS/RwyYC13R4o8U1PyRswqgl2iSZlMe544syMzR5g4NM5aYxW1D7M
B3wwrPQqF4zwZgZW6DK0jNZv5CLoDzWzmuKc70lUr0S4cjb2EBHXUovvr7HP/roj
ibMc554Wv2WnlIQyRTPWqZj6Aa7xE720dP+WQ/kcjLvFuUgZj3ak27Qx+TL+eUjP
crnPnN4xJbOypHmmjU/hd+3C/Rpj5CVLnN0Mh3O0rh2sAoNS/YvGBdBMgQi6aJ4h
t2C7JsjbjfGOCWW3fEdzNW18IiqpFFwXNM1dpEdlYtDnnGFur8T3yCodjb/zUrfI
D4DhO85Ul93lMb5W9zre/rZp5J7oaI1AeeiAoSyv9lxQ8yjHgS71U/aHTiJqOpkc
MhaDQwl5LEHy6i8KqviJ1aYHccuHfKValnOFzgveJxhDOoDK25UD8vyw2Chc6SWc
pGbN1bx9FqJb/zfk6SWipLL/eQML/vP4P++JrNjKOdrIy9iHHMTUDF1Q3OrbnKA6
UIkCy57DPg6gg/T4cKOuOX/lOUi52rzDKvhycVaenPJztQgXogSS45ItlNVGbQBN
PHRDq38lw5u5xhOOhN+pz90xiyiCXeKixUFBP43GmzlWP7LdTeqKvpql1esWBEbL
8H4N4uylBcJ0VdOM48QwdOVJJJZjS1vym7LEKIIIMd2zrnPqrnkWww2IxlpCw2t+
bENTEnuJRoC/JhOgkTSrc9R5FOEu63eytQfsazfglBaaKUQsf0jEyPxDcoiFWqHx
XFI3oL67E2a8F1WCKfzgeMSxcxZSl1exoEML3uiC++Eb5D1+OZazraZYtrF9CMYG
eSpFTzK0Ov/5IyYypuQsaqu+wTewWubSXT0Z86G5fNLeYJaMpSUSP4yPBhK6RKFe
hLuq9gKwlgpUVZjohgAs5Evd4ykXoi+H3J9DihgGXSbbzbHWrMm8is/MMAHOoZLz
t1WviautqfYiQ8ijL3Sop74VSgTtRa8YCFEcrFHUKhwPtzEJqvxARoEWQZiAGQhP
xdkAYnITkHPbmcBOuELIyDuHM+3XVqCJBRZR41rr2xcBBkUKw5c4vJBrtWcBp64A
ayDA/0AyTSnCjmv0qJUgDhW7nw3jxncUl9SVCmM5v4nshTsMSzeSbktZlNz8oRD+
I3ofJhjaRm4xqStookfVWZmrZ/oSVjs7UaXCNtZ1VMV7semXtULkApO8HnnKXS3/
x7sVYpxBa7mIRyLtbcAEa7KxRooA2y23b3tyz5SBNEDE5FZhaYA7uPkegAIP7Tl6
S4VN7EjHePNFkNWanXTDaDFmusyMQoLQ4parmPzR5hEh5w8fXaMtj3zRpPkB2uwp
C3OSMu2rHucHlTAjpx895AOzB2kes1mdllEUq0fcJgjVdWiIccbLVBXQFTMyTt1D
SZV5SCI2ph3AhHUJQDMicKxezHuily64DVk5TVBrtUXolKLmX7jn2t8TEehgqpaY
HWWEyUjEPQLHp/4SuRtEOc2/W4N+MLtTk/3HO6TuJNR3TzdWJWJmMe2hCvaRylte
JMHPvNNnqkhzXfss0Zd3C0AAk0EUcsYOu0lnpupqT0X3pCJhmVe4hasAGlN+eL2q
7tjREJZoLFyjnSPZTl8e4/nOS0v5B4sr9C2o32D/n4nwRdvPthEkDiBL9zE85RNz
dml3/h1Vo8Yy1zZ+gDo89WJt9k0Tqs69Uced+QDa2G9gMnCXVa1VcHZiZ9W+wdQt
qc9NQ5D1pOWleMYTo9sToaJ+DewKHdr6of8JbULaKaU+lQR6PtdSq6kYBOx9tUIw
NdfKcv5Dpzjp67xq9wxt7aYSfmeO0y/5zmMY7G1HkQSl8HWkP31IkHJiwEGFc9PB
aEtCCEaljwJ/FyQcWE9WtESrJMDmJqHQGWRCaOceJs/5Fhm+4w3gaL/n4U3IL0wq
i4shnXw265SEbMRMki6mAZDKMu/zYzOZEatdl9wMThsSg+DKNqnarYI1ZT7pf1EW
C87JULLl/vkITkharEGFcr38mKNxuV4IaDt6Oy7b3vEMbe/bunsZhUEaykD95saw
FRuVO0CSJhSg4YmcWX7AX2jOQMNJQGy7KgxCLM7UeyEx2X6btv/YpI71uugdcAEa
4X9BjWTYPMJpG3TXz5+cgEeH4ciB1Dv0+Pv6K9EBYzqP7AKl2UPtJ6w/Ofx2QsnK
va4yETTd4ETot8xCSzbfv0SRM4M3O7KvHsOHeKeL+nV2s8jxxa7dTdV02flro29M
MmTBHrS7IxsPMu6litfdWdfP98zF+dESV92xyzxw0oj2OfQCX6b0VipcKg5QUqG5
ltICSxHzLgQvXGsCyAruEdfXBCfN+SG/n4WpDK3saIA/iEjwRzdm/OOUqWwkmjjf
2ADmzPH69HBgs3a1Pr8hDQ9dAa3oB4TKZJJJLyKtnRVZaKthwNCy4U0JqD3uIYBf
szZQKcPEFrP8FurkzuKUEBsMvDudGWc+UTQxcUYhQ86+osync/ak4uQV+pKGhBUe
UPr1HZy23AJ00wwHHwHzYsDzBTEScNwtZ6chOKFwl1PZ27ySXO8ygePR3Th9ivNn
QuPX3p8xXOAwgt9S49bbAKKig42ZnL0j+KG8qlXO5O0OesxtkGYD9d0z59bLOnDF
o3LnCke8IzC+oQS7sosvU5FIpwVLb25TibxUZz61trYOemQkQfaHAtIZ0JRIoqWK
z80djHeJJ0jvMumNCh6KcmIYcjUiGG22dkxwtURXLzM//OQ7RtlJKjcMHxtlLrvQ
q4Ln2w4fvRY6BCo8XuC/U4IUVAEFbl8Bva4/Fm2KEYzAjYxgc/6itKtvSwgwuJTy
cvoNkgCDMxEl/BYoWL0TeM/DFoTK6uTDhyvOoyJzWIsAdfLSU9lHjPkMRy1JxBy+
Cwg9+14EL9A8ryoUtNP+hhswOC1cR5j408h1ExaFVmtUnYBJNqcvf/IotvW/aS89
V0KGy6uGfGR0ls+V3CwoOJhLFpXYZKVpS7q+a/+pnATkowVpAMufq1zjG9htbmbo
akLUxjng2m8Gl9QnfgpeSvbfJ7zlcW+PUCDrq7p/aTal5fdxZIeQjq9T9b9MJF5G
O2al2XBc4oRpLwubQArCcaBM93eWcIQXLVP/Q4JZfKOS9FGOnX4cIdzUZ4JKnvzP
eMqdYgK7khrFrpgNJejrUymYvBfCmnBxHeK7OlQug/3AjNTJRsgDyTmCRaLXeTvO
z+lchJRpMDIYUFj3NTgnZPocKN9K3vQI0pIeelXmMIsrgmf+VZhhttQkJ6hG5i7P
iZWuXw/vjX51+zNqUwTQlWzs/G8rL0pY/IZFFN3iVfy2EVQpQvjLoteN48h4Xu5f
csk4gePbcQ6RBhB9u05n00zu8PBD9MD+01QD07ZCsePhalyqKapID9LpOtywbdfi
mQbPO+53YRDksj0puvS0qjz9TbfPrn9C5RdKsh1QtxDUdplwOqx+DU/b+ilfJ+O+
4iqu6rkdlcNZV2a8fUFz57X9wiuGFRcWgPrtTGO1MnQD6xWIKjh0PFDAUqUio12y
O6bioSxpQJ5qQd9RteKPT7jPcJTBe6SIGaOHj7gh7/Fdakl2dUkHiP9kxMrfZK2T
5K0U+dZmM0TOOfj70t0mqDVxrNjoENYppctJqnCWyAjPESnl322CoRVJA9tP8Pgx
Kzu6uHCGF9AxJyOOMm+5CQtZ8vxixGjyaKCm+FbqiRwjs+sx8H0a1UebUz3/wb+6
M2He2737gWSSLY/5CJGIPk5fJwWgSUSJ/Mp7JyoLmgrYFsJpye6k0aDfeGz92KvD
msX+T8T6tPIbXhT7PMQmzWo+XQ317Aai3rfuomuojvRGsRyxDWrMDumOQtebhME5
wm5ltXwWpUvprec7RnAXUwiQnpUCSDhoIvQgQDfcLh6rrzelCvNf/vDUbGjl+Dhn
rKW6xPU9ojNRHkrhHhP3s24IE/jF5iUSEi+6NPfxs8C7O5nq+l3v17NdWASiLOcc
2U/khNUaxejmckloPvoVYbGpdY5PhELeT5VzQUAf5/9ljiJVi7YaUo9ihoJvNghN
vlyP001Z8p2p08BObFplrbQmwKkoSk6BcMBrtobJwLe9Y8jlkZrrjZdS9mwsN0I9
Q/zXlorgv5NsfMRECzyYyt/B+HHtG20zQyYKXN+tqCAzakZxTqqAs7Aj/ViPUbRo
+UYraVanqPk511YuBhoAOU+wzMdH6SYfFsmRsjkClOgRGD998p4qr+SsoIevKvQd
fOPU50VtW0Trybm1xdl824FFwhFuBvqpaVS9O1L2A8pCN7ekWl22RqqvTIk5Ty3w
otbq7KLLpLEklMXDOtJ1QyEGkxqipkHTxwRbCA3okjNt9/Saq7wxSN5qR39rYp5/
WgIKS1dIkLn10rYo2Hc6ofTSq2EdYJ99C5euZaj/D5ZZz9Gr0F1e7+uOPaswu8Vl
b2OpgO+blBzy/1B38nAsJwUzh7J32vTKXcrFdFJQg62U5OF4ZJe7xuBP4VpMUu1p
KiZvJH4zpEFiXlL/LYFZLJU23Z1SNlofDQVsiaQkPEVnS0r6Sse0hYn1sWsyOtwn
oriKK7wPG7rJssgaCVzCwnNpsl/aZebBUVQd/aeNHwSrVAD1spOR/zFO+SkutoEI
0N/zYny0Xj9BkNVFsv/sKF3ziLGV7yhmswHaC0iIqycoBkCgJ6R8Jl/elG+Lmv8T
Cftuwo957BCL0kZH2fkMrg6uHUoxlMEqENnoCwLLJQLAvVGZDyr44oJ8GC5ooZug
EHdtxbDas12hBUxzknISCeYbbZf1En94OgPgahLJBgdlNnXjkvI5MpaCeiWU0Htx
7JYKotAXhF5aBGpsz+cNVP/DOldSWq2rPlbBGNr6992Sg/rb57/0LWIRKodqAs7V
gMV4YUbagvBoaB24BvtW5RZPfrlSRF2upN1SoKEeT7u7G4FaQsX/umhhH59l/Tnu
zLk3RKeSPgVFrRd1gPKCdjio8RWxR745NMJ1asuDR7rNzWb699Ue0wUuYK/TZCIt
W3RBfKwtXbWRtoDn4Q20Hx3+mO1ev2Q2TGZgbjiQ7rzh92PZQYfgmSjsovlLjbqN
yBHdOci4+ah+OVW0yixXYsbissXOLkQNZa0r+Ga/chh3czKRYbrVxASdYVB2PdvJ
xdyyxLSLQ/cyfGlG7myiu18QL4hghqWjWIwYQDgQie0kj5ICvbk2nwB6HDVAV6EZ
Ix+ItNnSwUU3k1QRZrbRkSpJcmab5Ire4XaqdP9D4u1d5gUeSg0W2e03DLJ/55p8
94hZYBWnkJgHlyuG9OrYHHYpu6m8uzZ5xOjGMK9CvwbEGfIqHrlJqSOstbYCL8Th
ZuIOeIrP91wfHGRwbsczOWPQ8RCBSzm2oko4JUVGBMdUZpYIBXYIW1cjeLhL98O6
OViEKGiC7iJ1fwmPdR0ZLDwjusQgyU46CKTBrlXUuFQYCWCA7DbrFZ7QPE2DPhNV
sF91w0DiLIlBOGiZHb5RMNlqd81oqJELHkg/SH//pfRUVnaGxY9sOy8DgRDSvmIW
NLjp3i6cjlmWWJjqvNYpz22G2p7Zl4rAd8Ai2hF0DAN1jgn04J1P+AYocwooUeiW
8Bbt7EInDyT0icxikZH4H9hG5tssZpf6hIYiClHIZ6dBMaY85BvCbvGuQQx2Ii2G
lCpaOn5QJeMR+3pu3POfCk54sPxWqVM13X3v5tDccNTYoi5f/WaSzatDe9W+cggP
zB5bRG5iIyotjmvpoOn+PeD4T+mi/9eQaqdiqH7kXXUr8ueyEazs/mr6P98FDOG0
uDlRAjlSsZMMp73WMmtHW6QZTKdfpbPoPYPeyP6o/kWrrebFn1jm6PTCgB3F+42g
NfNxHmO1RI0B0zA3eyegZERGowvGy4TTtVuSLhVUv8VFb+/ZN7ZLEmNIjA7cS3ut
QttzFCLqv5YtLdCMCRY4bab01X6rs3XuK704SAC84FQeSnBEA+yghLfVbQv8/e6F
UT5koAae7+sOrOEumL4UOGEJpxy0buPwNJgGI9p+uo/Zf2dpkU4WuS5Wve3OBe36
n2xHhCV/mjD05CkhRqVlEdgggHHZ4FAx7WDUgFcKf5v5S9xSBWM2tf8uep/cUjK7
zauAGIQAcQ7w6XURThK3czWqcf8Ffm/G7INSCzGTT9cmixuob2zghISaE3cpAkS+
CmDp5Qqm0c51yHUq84WBdXj9bTe1CjhdHNc0MK/h74TTs6+yQf8kmycpK+zYqYr9
jCRUdt3qEIHbvUaqIXKx3ZMcvk5QFr30TyJtrsBHuH8kE0SrkQ+Br8wboSlDIDIt
MdLdlPKXUYfS4lGgeW2547bBRVwgDbPCJ6ethac+9d5Q+0Hmlsl9l5Z+y3pkwTxG
yq/6Ui7N99U00zj/cDS2eHlJyVJHL5awP7zfCM/DBPplGSbgHzSD62T0FGCX2aE8
pCCPrMKHTeJZEtq7jGH5KchIkzV58azLrbogKVowa9ZM742pbQVLPEaIWbb5Nmer
uPGbWRsxSaR1JsRVDET3Ft8ROUysweoPijoB/R8Nb6/Ba7KIorx2Abo6Rak4EPgd
boJGwRJKXNyvbLX0QWgSV9tvr2TV7ENzz7QCQWAoLcXhxXiV0WNAr4WW/4XxatvO
TDW8A+OG/Yl/Bnkp8R+ofApw9kZOlCHft3eH+/kWgyaRxjLvSbI/cm32OQbs1K8Q
8BNGqOGXj5LgQ3PjbdAMRlTJyxCdrJxEbqsrlYtgOtY4HJMwzn8NucIVInDcZgWM
Zg5zalK4d0SIKX0A85FGnsf5VFSQhsLHJpqQO1WLweCOHOGY+dgSKTfLgAnRGozf
Vibp+WpUI0WkeZ75tEH+jto5Nj3g7YC3aLmzrEBbCpY3Y+Px1cs99YAe3p9OA8UU
U2mms6S3w+uQdhDjk0EFo/TtQkev8+IyjM2XwnMTrsphai5OPzHRMoKQhsXS09Db
V/1Q3HylI0Yzl8yY8XQgnWnSmsoYL2POs+MuigIVYXWxEaCvqJg/AK1qRkqaMU9W
xec8MW7wpU50phAp5q7MGGg5rrZ88v9jxSg2t5n+Cb1IoPaYMzz45kr/491GJQWE
DwtAwRP7n2H8cMpvrp2LBOvKxnCXYgHogb4wT+wXfEAwrY7D0eoFhEmdJr8KphPx
Js/06tkefrc9TEqYyi5qEWoPNJJNpvq29L2PvWjR7SIcoPrOxjOQQtU9FpQMKMhX
N68PRcpeJDPWnynWq/xSJbehjO9MmRshnM3sbQ4/qORUXn5+oAdykuuKGDSzPAFP
MW+WgXwm9pLZHxCVRy4O8GlA2G5aukIAzyXF4Ct1Kir5HZoromt44moU3uBwuM6+
+korx+5fDih9T7bcUg9Ie4WiK/TwLLUZnHoALuE52ikBlXjsjRZXjks0sCtdkcuL
+WVHKCoGIEZc9NLMmQ/1Z9cKNXCe78oau3kLET4dkYquEu10+I5Mp1KfQM3SrS//
VHH3+uWKsmnN3mLPqnMWQvhDi7XsE9gwT6dSoI6bthcJkUPPygJqwiCayXbT++pr
jBQ85X/8+qXaca7gGWkjrr58ivXRsbWmJfoe/ZLKVwFjhgy0a8tJTRyptwmeYLUf
8+uC7ZO2RZpfVFLYv+52zDDwpGfa0SmOc/Rhm46gtW7LfQ25KemGWeZof/FrRmi9
q9u0oeY2jZu/SbZFjaLExR63iPbP0P3HHWN15bX28/HnP4bLm/x2xYB8dHKGDzE8
1XKzclrhOdxAtLz3jAsx+cZABJUgTwgtJfyW2UWM6h5XAO9oFqd+/Q+GCSNBn8Mr
iIvixfraUTU8UMp4CZXNcgC6hmWk1b720gYcKBUEZJ+qZDDJ93c/OhF+UGjPiKs5
4hxc6FvmsRDphu1jgs41ztqQstuV2flKxr6EO9GJc6ROd72i9TuyD7PhDrKl8V6k
UZhYrBm7tgmZz6XF8ksInrJ8aIqJmrld0DE4X/GkMSyDqREoGAj2Il5WzpwJzEaS
mFrFSz+l0rwVs7VwzoX8X0Io4ioGxteDTeF/GpTNGGetYDquJvr3GfjS4e7sAUIe
GCEpjUXwRjHyBq58KlIZsVZ7cgB+6hlK61cRvgCtH9YJKaBafJbQR2uUvUouv7Oy
0xtZRSl5h/6Y1L9bqL5u/I7tPvHr0XqJjxm+VEcn/CIWsoc6qAo+LCSiagM5K/F6
G9Yq0kG+QpdcD5f/G91TRi7D2HBaTRZvCGFL+CObqlvir74EM5GPArb8sVG6CUJA
0q4Nf/COxxEycuSod0eV+zq47jb/BSBDercBiAQ8l4xCvJU+SRYJdjtYduZO6v8t
us11TDKZBkqOD4yfGBWNQ3UoJtDG7+dck4W8Y8psEZ2vI0h+SJRd+GbDl4/qFg3i
J5mIzsiB4hU8F29bvHJ4j4VoiuvIZqzSeHRRs/7vGBQoQxDDM9db/SnqRZCaXcEl
me6p+6w+h9bKOQB7cyUtXYF1tlM7f2zxF6GF+vYeXXv5LUJAZkHyUzt1mHCHmMfE
AlL3YSKUtlgiQTeupYx61wWxeQFCrAf9THMkkz7fyvf3kuDZ6+ThKD0u14WcwvCR
prOsVyPLPqToWzP35k4e+LKOnofxXxohzOoC1f1YPl0zwB+EkIe8+67n1tAykhp2
42mMsmKaNwjLGZ4yFo448G43ou5K9R2DqCpufU4ZvegSLi4MCkXIxtX5nZhId0fa
cRqRqQbo43+fVtcjQ+imZlCGGyGZ7K/ZiSRmBoDYprwK1+jfYUZ0x8eiMqj+4wre
yvhkplJDgWpVLXnUVARuT3ykb1oIaG3M/Z9FJHOnowgn+9BnsAM4JWGGeO0awJoJ
qMPgYD+BjKRraC87MBqVXljz5WiOgok60JdDvuQ6+j5PvMgHywDMMkd1Y59ZY+kd
SYqJaBFsjy7DWKD+DgG//5j4XEdhAYn9Xi1rBo6Pj0MsJPvck+et0n61wnZvho4g
Twq0TWeDYq5oN3P1Fv9ct+0AFXu99vLjtYP+wf7rr4Sa7oF/G0qquQ1TbYSIkLZ3
eGetTCN3Pnn46YryD62l3bi6cyo2yWq5R/C0+E4hPc7S5O02Ak8z6hTlzjOx8heO
HyjJBOtU5ehYNkVKCoXj8PwZn5I5WIrjRWNW4x0V5FVYQiUMwPPe9rRIq35SwBo/
Y33lSoTcdY7WXtSdn9/r728Csc9RhIk/YAILKzVAeNLlUPfU6O1gicHgCgQE7eA+
+NfnXBalprQESxazPedB8wYpxifArbQdVQWuxQk1WVqblTX/w3FXfRqkiWTHyl9y
uFu3D2/c8zZCQf9Ruh6lm0YDjmtT1ZJvesKWLRgx53yATErIVBgmvweUVaw6vdA0
dqXwocmuR+14829oJezO/uszSkQrxRVWfq0J0Y1KAOD0uphYVRt8r3aqM7yaSnaQ
Rux812cLRp2F6PmYxZpmti8HXlTMSKZgoHxK/JqqXaDbznnAXvYPRT4+6LQObNWO
wO6VzLPmyoEW/J/B3xCHy13pamX51XBZaq2hdEyh6N3kuMKjXKyziJauXDM1nNV/
e07YLSW/Y5xVpPvo8FMgYiTeths27GbnjomPU1wGxDunyy8qkrnLjKUTSww5X03z
J7YjsfuEkIt5PiAPlBTKddgeq5OvMcHsLwzOmz2BiH/8m5HWCx3hOa8CmG5hwRYJ
xYZ00n26JaJwZj9JLHbwHiuZmw0AHuqmFXKLo9m9HSb+/Hn0512zfHYTxPtuuHkz
82ogzKiHyBbY9qPJW8lZNmFlMZ5r5zLDWR/zQKN37FpO90czsV9iI6+CP1DmAptr
WwPTpwV/ZrKJ6hgvG5KIGBb1nUj1/lF6pbgi6ScjcQJ7OHesUrT1FQpazMm3bsNM
xazAdLnZ1T3AUVJUyShGTsPo1Tj5sN5U2CaPT2XPRjHVVFMUmNj4eJImonstF6pv
HkCfIuDWJF3xF91Fv0v2EXyGBMO4NCCIMOWiprca6zrtP09s4JmnKCBKHRd3wGHO
/BjhBEjkOaNJp9lV8kZweMgH5jIpD/qjZkbTTwcyIu2/i4LNtPXWNCT2PB4oGod0
6BX2l11pC7CyJfduijt9qpm/9EsTtmn50M37JjY4OT6TKkVlVCl3xpzyvRCxouEU
x1a6QDfHSKCEdqeRER6Kc+gXOyoX2KFiDCO/8AYUzJ/YxFsrM4aZOw/beNZLIMzM
RRaLP/FR+7HucjhjHv3su2ar2OrNOkZTiSs0ZBx2RANA+Zw67V9vydAYg35D0Zvk
M8N4wxg4IeJCDjXu7aF4Gs790gA2HwFxCGgy5rXx/G6t+dy7f5dwocXv9i8qGNjG
bb/QDn89AMuGUfyeBMaHOHHUSVdVtWEsb6KO+zgaDa2v6cij+HBAUuXQ+KVHMIIp
z8/TyEP6gFjXu1NFiG7w4GNA4y+Qnx6lknfpChGx13JSqjdfAsvepA3M44jRDgJM
0xzmACaVqWmfkfv+Noup4EdMS2VB2UWJ39z0DKSSyJ+PrtpNPYl24dtkrdHDD3WS
UGevK4zva/pToYNN26AwERfFP6oI0Xxr/NU0/bPlPtABtsI9g3nReg2Xo/IKCplo
BojovQEcDjgOmF8pFgpo+Oe8/sxEYRWnUzQpvOFSe1Q2WqT0N9SP5QX58ndGDMUP
lvL00xp83NGfgSMwx+/4T8+jbXpiz8LJKMZyBZajrvSyEf23ycMtZxteKDVwVilP
Xpya5j3/oVVpRB6J8oKuI8vZg1jxkU7HCIPBb97qK8e6t66DCoxf4ob+uA8Hz/qI
RUcwWnUxuuuHbEIUK6jjVef2VgRG+e77P1j61WdTyaRcrbe450OaQlgk6hsRJ98t
uAa8uSJZ5SasmKzkkntSh6YZJBpMOQszLSMWvUrNH9etxO6xGJRYAoKUdL+FhmQ4
FulTfEE5LHvkqXP8SVJw93bPk+sOYtgkf2vQToSJpKVSzLNiqIBdRyUi0Ct974jk
scmgHNFDsQbfEZmwD18bafLd/tfSWqkCLomxDB3H4kofG/TP9iuZ2X1oHeGUbIDx
AT7spgjkn2FSOtvDOWSvbGOinVLAbJuAIzOpS6HC++XDSJ9FtmxNTXeYR0OniMOR
AgFlqT9bLSi0gcnFkcVWAiJ6luLL/UBDkZ+5GtS42twuA5gXu1RsVPMSr469CQKz
yHvEpX5RtCd5BN3KN1aa9Ejjwm4IePcynxoHKxGwLBp0eyOHfAv7mSoXwyoYrNq4
HfCUx4Y+PlBrgcnbp7ssy07URKI1xnNI94Qg3E++rUniFwdKKahJxLMH7GsNItaF
pgQZ9oOpIBuRpq+Sa+ldx5KRF4364EovaHv/UO1F8kXYnRGRMhm2lPQkvQyBcBoi
ZE0IZbU/DgSs1NKjlQ4EFlw/r+ZD0cMAoX54+EznilFAt/wFMDhZ9wW8MRTKYRlE
WeGzK6rzBRN7eDX7x1Mocuwtnch0NU7XtDL2RHobNfRrbI9a+KA4ZwKgB3NmFbk0
uFdhYO855uTL413CcEx/L/Gw05CeFb5AhfvC36JVidp3Fv2AfdEmgVVCvtqFbkh2
JbLE9ZXk+DAXp/jp5ovCCtc2u+A8dtprhQNAFRyEdrLIC7HROslPtSmsuymBJUPf
bJaeS1U8wl8D+oBsbj//bbjSnNDA8hqezgLV21oVnVizMlYX3wVleysmnd35nlW6
5PGhjAqbF5NsZeiMB99tI3SlDbMQZbeCZb0IKj4AxhWITPvDIJZ60Qz3QTDf78Wf
nE7JTpnscK6DSlW7YB4cn0jN7NCFvChiLdNf6S6Mj3dd3LRx4+bmX2qfNUcwQzCU
mTQ1l6G7yqnj7hmsOY+Q/7ZYOU5boZRbB3d81nYi3xRJasNZHVtYD8Gl8WI3h3sJ
BOKeN9aLyc7MGwFE3LSPFcH3CQVVaMYwq475MLPYdW4Z4UlcK5wpKeoSgJegg/YO
yEa4GlKFZkULJ3XQ6fkUbkiy33AF6I3abkbhY2LFINrrHkkHUtjiJ0Ei4W8W5cyg
eB9Dtq561i9jmlCN24JdLkBoma9IS717HMRROTsb0f1qVjut1YHYa1FeN3MxyO1/
LR+ucx8yuDVVqJ6/y5B6ESXM7kBOQ4NxxT+QrBDJHWNPqn40aAOCBbYm2aB7voqh
BajcFwtn3XQYuMIJKgSoWvmyvIu/tTFIGV5JH0/i768ts72R4XjY3zaN6cr+0mxe
aug5dBwbwMS07vRiolr7UVpo+wq89ZTQoxYRoHlSSobce6naDpVGWCGgOZBmRPis
IhJjDNmZg0tck4Hobuz4sBsfsy+XV3JJjSmOoFyedypulX4GL+X3pUGWzOgpw16j
9r9plooiIIJyhkChjSytfNH65xsTGR453kfJt2wb7cWc8bdQCWjmp3acS83aC9vb
oj8IV9PlqiWkeTgpXRKg6nYdGzHeDZaJXeqn8ocGb6Q+M5RT+lps54MGzv7f9P0y
nQKJX+dgm32hacPkZFZ0JP61jduciPBuJZLgUFvtxfe6nPh/5z9cwoRCuLGl97KM
IOvdEjqoJnJL75UxmZNirPPREIsSeRT1Mhi0zFsxtrYAvWtmKXv8ZkwXOHIv/VJz
29Vq0sWw/wPnrUYHn88BYz2dl+IzDaBR8IoqMkTrDKpC5wNjgs7ekMbes1PR29Sg
f0zTfxaYUxQDxOTWxAqYKwRz7skX5ou0aqpCLJJUz9sqmd3Y/2kRDIVCjJFPuGFN
rT8HMGrDEWmv/blIRod3w++PY+S4skqQKKimp5Fc7UyyaUWqXfr6e3DozsOtHc5K
5Atq6k3KCx7CfK1Mgvn9DMyFBOL7HyCm8BLHJ2IR2tb96b1bRDhKeCp7Mq7JsAWE
AXnV6z5q81MFEhi91wcO1GS/+jqu9aUnLMQBVk/2TiOUtaJ8XtRihBBMBOSwF7WE
lpOlni+6C5A6A3wQUtKB+id8m0hXWLPjjFi9A+MX6dh6/PYUP1C2J5E+MrDjlJEB
8m2Oe1KPelf2s8Z+t7pff6kkie/rmfRGgv72IgK88cyXLVTKDcepo2qFRFN7VYsc
2SGHTJyu2bLSM0H6uQnALDKX/td1RFGRq/00KPV+hoWZJd2XDEZnJTNpv0yUhCHG
wp0ktDsVxPd+Fy1flBYeDDLmAYxyVm6i0+AcLxvsgC4MCesoNfNZntKi7r7x11N7
h0uwG4LbQiyYB4Bb7z/tUyo5RJk+UHPh1A2BLwTKXUU2rvkvLg491wdTytFYBDX+
GEaahS4UaibpX2pE/7ODwaH+JZmB+oaPqFeF++ebFpUkPQCDbxxLjJgKvBMbT1nw
cWhNW72GXNgrfbJPUpoYaTDoGWoK0bericRLb0bmIYkhuo/fsy+D+E1vfA9cnOr2
9TXH3DIHpR4Ttbi+YK/KUrBaDdEdg/Zv0xYPkhsEy702q1DtxND0BOOYadqB7mdk
Um0GzEcmzDJuk0dNFORbxjhqYtsdQiHgE33fbtsJR7ZxDS/4N5m/ZSKah7XCsNMZ
Nvv9R6pOnDqm4s4nH2BhVS8K56KBLC2eR7fVCP1gqGbhdC0SCsKVsvV5iQo7LpeX
dJLRLGz0yXwoOvsrDNAVvUavyU89S7AejohB0iCi4Lwjr02/pk6HPrVnciASVsL3
Z6mfki1lUgqG6aGOU9GMMdbmOj0r3oEGFeel7H/6VwWoQe//5WFGr0rlhwjsUn+Z
afdXB8FyHIQQkrpmMYSFDIit1e/fPJFaZX8IGSl6kEE9cwBuRiRZ3hsnkmRx8UAF
3zh4+kxCNeco/FoJ0NIlHALOU6H7ZOe+IaoMQZHSbvDjv9APLXzlHXsY1OoOKLHu
SMrr0RHnzu5Zd/DQ6tnjvF5NZpnZeVZVB2EpUiY/UVaKG2y7QEaiuiyS7H0m4SJl
vmMUQDntconadjpMZ11OYA4n2P3EIOakPxUfdknIrTQVFSci8/AwIKFWq6AR6P4T
BLLuggwX36TZUapXhxr7hKoO7tViHXBdInaBRav5yad5rc1GjJIYkO1Y7PvWEphf
XWSl0aKbRZW+2RpJtBnEfTcwS026qn11Ncell55469y5E4wTZXSHfDiLNSz9Q5vi
vxvSXJddUbUk25tlM7PWJlgshncjU43P0doq8GUnI/K8LTpFWjrt6C7kBVrbD/1K
f+fYP9OP4aDeRyq9VzH1KbAVeyS1VJK+7by1cWRBoPDPK94Aebnjl0tCWHGtv5Oi
ALq3r+cxxq/okxsUnKnKsgXxczdZf7IMP17Jw8vtmvfpQw8q8IJp9Dvig2WzzmtF
5lTHH4zwAshuEN9P4oFPQ/+STVbhIWzwswZYMXTe5y4QijU18VwMsleOAKX3JCVi
Ukm6ugC5gi0LgL7O82hRlAuaUpvLJ/6I2lCMnFxR+PVVd3XZYt25yHHUnleWWXHM
9C8R3LEKOEuA9TKR6DurOcruSRGkxCFstlasrOZnHnk=
`pragma protect end_protected
