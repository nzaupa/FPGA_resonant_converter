// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
V9ceV2dfnzYjrd2equZi/bKgsMYE9rZJ5s/K35W7k1DtDquIPBvWVBXmJA3VQMCQRgLXeit6sm2G
0lt/0ABJiU5mNncpCleOW4RHZGwg6lvwFKeySOk7ktbnCSdnCxf2aQnCM1P1ebiTRW6G90qV7m+b
aRd+0p+IEb3SdoCithXbOIr3FXdlYo01O2xwMRxQ8CWMiNXBJKdNwRJeq7b8dntwL8gy5043MXyI
AR/GiIvYyo8bvCAR3wbgfDx7HhwH2tSpkj+RZB0AXH2H5JGQnMbMwADZfgKoLmrESCalbcF0iWef
CxRL25BPdIOBizKMpZqFF7GUowIOqr7Pf6aG7w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 21216)
sRRinFhk7lBNmzlK4A/uYG/nmXlxDBpNcg5BqdoEyAZSgcw585HiwzX2EoITztlFbsP8GRa0djAk
yZLGoOzWBoGjLQ8GQ2WoafToqOcTF2+hlKh3Be6X0/WezWjSmv09ZshsnEV7QCZT/2MIYIwyfAgE
aNMpQDQgS6bvZwgyGc5tM7SLIxNbWVcm9XymFhWt6HLupN5DxskmJxQpjFWiV8ETCMQXSBRMKSTT
jwbshm6wjabzizSTzASjyf5gNJJ30th2WO/sVX+HNTbL1JzbMBnOswMhPh/rfytSzQKA0gaCoxpb
oCnJYIauA5tl/C9aTHbK3j38VFhBjFSPOr2ac5T4pbuDsiBMN3kBGabkuGRa83bxBTeJ69XFuDzO
bMnugdP2nZdU3+cshxTawVR3uhMfcxF8OyVNER3O2VI2iT2QvSSOU9RJzSb3FXcnwJ+GWM4R5ZMm
9Nd//UeyiBroWkyZ8DbJxWFk24aDS5MTX4D+PofY/iS57ETg7GAWri770DIfQ4z61mwnVP2A2g1q
LUOgUTJOvkihjUPWlVdLUz+8QHH9XG6C/mVBGPnzOdgLMhjIpVtAxUfbrPyOtZjNrYmdhke8iAtO
UBFNk27nV+btTIUIt5CAflqKxWVhV7AxcncD3Q68Gijphc/+nJXkSltCOc8LaWuRevi2LHAM5KsI
m3OMM1NLkyBGKq/cmolKEQyFQD57u6Z4gtOJqg36Nff4eSLyXmIo9AP0wbrgtCyfLyhRToJ9Y/tp
aAz6jkwN7F7bQMRj74N+IM+YFG2r0LLll/tjQPzFNGQ4XOtNiBzfOs/9y/N70bGim8mjHIqHpmxE
0mfMA/mpjkDOLbrqeP5nMVSKYLMTAYAGkkgi0QSSv2vJ3F37qs7Dse4uLdQokFeqOGuhaBd7zxgl
fASnf4dGLXNtx31yzfUAWLVYJVxG4VgGrfV0Eoj1320rEBw8hzCg0vqcQmGV51eJq2jMFoPRNQ0y
X0+3S6WfAvsuiOS97qjNq0sZtxdK7Wiro2Qj1DweL3uFoHIzKFTYfZppSDQZ0BbX10ruAFE2GgZO
l3zfWDID3Q5/IfPTHplZZkFS+38+sGyVHMtPXqDtXYGp6h0TSTYsOFaFm9+8L2/AWaXXentAqx4m
H9pHpfBpMdbY9EDOeDo2Opgy+HEelXxoQs9TTyM64cBwkfzrnh200XQsk8UV0lGfCFKEeLtR1ei5
QG7GPP4z0O+AdaHbGjvF893hemgPXX1IP+9pGGw9jmAOxK7wqfAHeYOctzit26m9mFRJYjmejNj3
SzGxTINAhAaM5njDCylfyBpQlJOmcADBJSzt+er4jjhFAsgTg+kJ32EJTIzkCjvVYRAoD65Nm1b9
KKFwsJIIKbgH5m7KNYZpeinOj28kU4g+Ew62a2XAnRSjtOu882ynTGAftEJUqcgvgOpbW54Dgi/N
/swrQwuQyFW2DAf80XQqz3UlmYecZib1R7IBKEibH9Eob+nCGdD8YJgvYuSIeXNs5gHAsACxuS39
a2OfT5wpMo6MmH6CyKeUN2l/mGHEfMdV/49Zldj7zhyppo+L2RF72vuzwLvDys77t1qDF5FjWKzY
+Vk1zmHxDe43bPhrd2Z/ZRztPklFLtZDuUK1Bv8aV8A8N/DHGiQnbCW4TfP5amcDGKfrjEbMo9nX
i2BCIFG/EJEhbpdPB2wIFjE3n3YHOw9uXbjO9YGuXUI8Nz+dhj2KKaalaTwYL3/vB+cu1hQNGhV6
fnjgymos82M0kgwrJE+I882B5RI0hm9KzwRrM0RQpJE0RnRHkMo5A0PMm+c2cfPXnPCwKxq6xjM1
bf9KoheMbruOHqtjEjhICCUQ671PtFa17KIsYPjRwWAB5blcJJIxSFmkXcXkD6kHTgLbyR7LdEOI
BZmDrvGQnu9pPi0nY7zZjH2b1g7LX0TUOKtm4uBIq9R5PVQ2p4A/Dw1dIo184NNYGYoKK9srlq5V
MDBGtpYsSEthG/3/S2AtZUUoGj8YSj8oaZalO/BCBecCxR+qXrlq1/krAsL4/YJ72lbDTJZP+Wvg
JWk2EYItChK+a097+yeKmwLB9xg3/mbiIVS+yKafibx37gZWn2+IziRBQRBH2zwkiqYd7ssfZgCU
wGiFjriEiwDq2HGJAeWkV951SPhpzagglvJ4JV/EHaPbvUQ+gkblKj6LazPIXUliDn/tdgrwiprQ
os+OAQAJTbb3fvCfViN/n3TUO7sbKu1Jv0dXcnWFL+utjSl8Mlm3FKxyLr6vdNI7iECaXdCte/gW
rJOM6Un2Cd8NRbIoq7MeFhxrLOoFwu3sRCGgaWvDIhRZy5437GjkdxIp+tHFSSm/CY301ncV9Flc
9DMCcvnYn3zmhddMqFxcNxH6IEOLm+h4dfDcUUmRH7fa1JzOUEFdQK1Smfgf0abn52dEvWfYMHeR
vICTw5wJ9olfFiAUTNnpB4T0kFZe9wo435vs6kQK+i3nxjABj1Q/o1CbahTzhXhHFfdYMIdYchVF
vxm+yF+r8otr24K67dB7GMc3fQhUn1jS/hiZEmjWESpvmPb2+2TTHmYf3okqwB1JvajPFEqW4dGF
XVLAJ8BG3EZK+JBfN3OCAFHPDT8q4qYBMhunyWZShHwSY7wDLg6quTUjIXcy/ZkV6jwPYV+jG4s2
czwc/RZE5UL+tg4h7Lrt2mKTMc/NuwPRNi+34rDuG/NIdKX58wEK5T7DyP2WyFGBgyYdmI2oklEz
bF2Pz5CSB/Q5KTEkMBtyADy/QARfevfp1yqVOOh7iBxFHDp37JNprgguw3e3kXflGVztgWTS8BqY
pY/fOd+oZ+ywABmhfrcrXvqvDUWxcxxEr4BP9iUEnVfgwrADg2l46VBiUcOceIDEtdxLHOOr11go
ppfYvJ/8aTAXAFLFKR9Uj8JpGGoY9LxMx3c3G6XugYEekaMytmkLyU1zVG53v7vNeBj/E2RSheRx
F0V0VjugNxSEJ6PJTAmKWBMAcRgJ5zsRInfodAsR2ZPXYRFcg3waMvgOqUOIL/SoZErwWvM8TlsX
L/7vdAlAJsl8Iy3F2fnoJsQWFEUUSQ/sepkayF1Bcz6uHLylVTpMe8UpdrU72aIOrC3H7EfIedGb
HL3v1tjx0v3356rRoyIudie2YChzAiFEa6einU1xhT9PrqMZNEfLq+Ssll7pFFg1pUkoHPbYU/s6
9URC1h5NSW1b5572zGsfwnu3Ragd4nbnaP1r/6ybo+Uid2BW/D+tGZ+WLtm7LAQ7e8mjiySHgMx1
Wp5cVb63dRuaVUULYkPfxJ2LODgWy5O3I0jnGclKGnzPIkT5SIYrTmNGiDq2aZ4cRzE7l0dzsqoi
dKq1W8gNhke3SrY2QQHv+fKAt3H7nlBguXHocbLUz36D52WjVCkq1f5OCBlrsNzEdOmge6q8wFs3
P5BBrQMSyfVO9PTQnCqqOkU8eEIfCVest2CA/78jA3h17alpm3Ku9xedHv2ItRkm/arbzr9MAdRX
1JbyF+jL3G+LBCvcgGZExrm3Itw3/diFotw3p4b33aVgq9kOmMPUay8/H6SsaqPk6Qr67y5uKkyM
RzErEFgUH/wKF+ZAz5VVi7BpaYhKPYDNXKrGvr7aO+cRW0whO2KwLdet00hHZKXTkm4DIYRvkM5e
rWnK6IOubvstooo9Nsk4j3gfTTAshReO3hr7hT1a7vfgq2WnKwOra41cnFpBDV0XttCfcDxGU1PH
J+pO8m2VTvYdPki+JrxdUJuXYNbSMXb9qALJ3bHnyAMVqveJDPRcr/IqXU0qdRgO7QnWS/YABEd4
JvS+vnmx6i7cWX1Z+z3P1G8u5rKOJm1ytEpch+igBc4asZ+W83D5WnmmNjZ2YxFqKQCsGRxYZcH0
Ec6dIx3E4ctWb9yJtWvMQ7X3f9m17DCQGKlDfbWrtFv/ULeokxuWHAkFCerdsPkJHBNRcOZz9uFU
QW0MCZGdb1qgXCobnOg+02LzD58/EgmzBbFcUPTdduhdR0umdfZQHfZlFUeRGJnbUA5BAfqIBhTg
UcCrj3Kpd7qgduEfI0/FfDn2gJ8UiFoB3sd2vjNEJNql9jm/hC0/frQFeM2p2jIsK2fxZ2Y2g1cS
viZnYvo5wtAZZNOtPTSIak/DzYoh5Jmurf12gcd0yz8RVjry0cWlsl81coDN0nUSG3H/+5v/eToq
JobmQblDZIbxFq+k3tbOG+WQtc3M+8szu1ny/oDgldi3gQzGHuokswB+5VPSZSEznHzEvDgxA4E6
1zb3SQTb2y85KN80DXDlUKWe9K5besIT+L0Bn+wZvmEP4upFDxFsDG3d3+TXi9zrpq+gJnWa6pba
P7liFdno8ZEVtVrcoH+f9F5XTwaYUbXEiXn+vc0Ki2MgKKNRykJH32XYB96i2sJ7x17efzxYGPp0
zGWPI4M0iJ350FEBCh/Tp5LUuelrNfK6TRXqGo93amZIobjV0u9CWiexrw3m0KxJ+MrqyHtCVLaW
s7kxZFCBjaJgBPHThMB7kDet2hjtSrNy0KV/NaRTIwbdNiXACXnWa3C2lnFJ9ZdZrOCAt0S4hqy7
EZz/3zn+ECH5pCcIvPOs2iSbz83yDp3LeMgwO2so8r3MUKbb9p7UUiLmvfj5Qt24lQMldDnSJpu2
5E+t2/kr6tQo10slmkxJq80En8vN+X0WjrDt/MENgUFMLCx/zA+IZATqP/gIcgFl9Z9xPCPAPtXf
KCQP8+i7gB4wuuKmBHcpdfJ5zniJhpsLuq2RqRtEi1t+Vl460gG6ec9NXuFtKSUlKTT64mpt9sTD
xQ3VeB8S6ZzYAbZKAAuVb7+GGmRqKQHgLX5OaJUt1xE0N9Glq7NF7a98NQW6nbrrT3/DzzQXbnnW
QTOC4XQvrlBSAmjfY2OBRw+xdvodRi87DBwlAzTTlyud9CEwpKmJc79sqRVr1GDxj8r9ljvCHJcr
ssNymd2mScbw0MnD76RW/D72yu2GjMwgRGV0pE18QQpakdv6wJ6MJIOM5GCNls8WYWyEtbU7KlCv
QwyE8Izqc0efSnljRwkQmbnVSzOsA5MMvR28Xo6VLZBdmHa1+GTK5aVtTtQcI+KvYzQUPKqdWmq4
bfCnxHwUIcnN2RDdBwTkFy786p9fXX4nHMpVpQZIXw5Z6vg6wqENMQlZjMz/3zdarr69sE3GVbOT
exysd3xWgdsaR+J86mYy+11fsGzGB8dxyDzKlLZ1o53uCL9oLU7Dz/ANH88sMtrDcLsFLwqYmr1d
W5irteVqxS/gNlyQPLsnOUQQT1/9NW/lVtxntY/BnLjdrGkbE5jYKwIQ01m9Y6MMvzWo08hBBrQi
n3MQM4vnKfVg1o+78I4BE/yaxzwoDwbERkk4Iy5GC4qwJQcEw86XCNzVbdtRZ4CFjFVYGEVznJ/y
1lX4xpLnKj5C4VCyNb3M8LS/VY/Fq/CdtV2qxH0ctb2PG7vxiFF0FLAfG7tVF+3xsYRzADifwzPW
epmuFJSAbOOOIfVy4H6K+0aaGgt+aaUeFrVXL2+d3v53EI/Mz8ql+AhQkHbiC5RB8ojGmOxifyDD
hNkHRFTzDLsFPj2bTGUsMcdyXFMzYAi4xybl89pyOi6ib0fFFnC4aURXcdlj4pSF5bvkU6MEA0CV
ZefgKpsbmn8rb3EqdrHsvMwW2MK/eJEQwsF04D1efuzR1VTovgcTw/WT2ZKy2IchP3f/hLQDuWVY
ESB2NimM9NKgH92A+iTOajfAtxgHdJYWxBFJbnQSg3l9xnU3Lp9/hrXjV+EhqSZ7qfjNG8gbnjBn
TzhDbrfTQ1sNrcgVE6vM+Js1nKFBTggBhXdBaNyq0DSYunxp8qcrQJHp7kAoDMgrQXDbOs5KcGzg
gLadI0xmTSWvhS6Dvd9GnZHRRxqcVHES92oQf9H/3R3ZqeHCt9+1yTPeyPGxqZ0iDexQsmhABFJt
9gu2iPPPbAQewNY4ssRrCG0SLqccVVGXEseql7goTQATJ+lIs3mqy56Hj2+1SqjmzYtC/PirgEly
0CtKwS7mssbYVPBDgYQV1Mg8UGx0yY/gPPtDPcxZ/1oopCogeT1a0cViSGE1Drxw3s3Do+chBdM5
H9UijRB8yoRcbFzmdPF+BD/hEo6RaJYz4sJB3tksC2YN9PGZOOLQWL8gApLhjQizxW9gDhnk6zxV
ojiwM8a7LjEiz81bDdFybbwZhz+JL2bpmurC0mopV+bio/dyCBkmpABQ7iJL4wRhXlL4MD6xPGNb
z6nK6bUawTakidJFvt2Chnoi7GPr6iJ9Ps+ttJJmQtOlfQWCSaSDp6zIeqVQbuhUDRfYocN+llbK
GvxKdniDJWlXvn6VnY8QIXdhJ0lgIuy5LLcD+ftVICyOQKR7z5dbpO08Z5NXDdg0Rk4lBis/6nZq
0AFALaxapn+F2tQCTTQbvdEUIGCkLfhhj2zZVgAgAg+iyz8erk9izgfsDS3A44L5fSZv7+5uDFGv
0HNoKMyRYUHCBeyRzm2+yFqZoDeMQkyATaHpnr5uVKiKZhR5MA7EBst8fhOAy1msabecENN+QDoA
dTMf43fK4r25072HB024Gjl/5ZeRIgGaVHCM5f5iRxtGSBrr05EVbyPSBePurVx4AcQ1GROfSKtV
llvUM9to/Eweadl+mhD0+iuHKCq8F8BcnO2JZpn5XZPWNvd2QE+xUlPG8jrv+vzRjaD8wpWjKvsp
tpEZGiq70LvLzswK9112zOLKeV9y+1bVAkCGujoLHHWojp3DXVRt85xfSqXCLoCYE+9dCoCP0MGj
Pb1HjkAmVltUoNkW8kRHKArlXr21qs6VM60gBjYSJ9QmuvpUZb0oJnCvca2953Ip1aVo3t18STeQ
roVE0uxelS/tt+27O5IwCcXdYZxNkZ/X9IYTYt+OLnveB8d+RfJOEnSG//dCM6PpymCA1CLqWl4T
jsn7ehkibVyfPDPKieInScL5sPELmAq6U4jonNzr872f3jGDI1rPxI3ep5tcbu0eH2t8ghDqHq/0
v/v25zwZ7h2BqYQfDL1Duz9pbUuqGc63AowW2LdoxWh790Ki8dC9T93H47vSgspK2gEEdsi8iIvW
pYDF2H7WfAIQ/8GhyBuccKYpAcmomEnQNYv4wBcsB/WgIp0tlg5OFlP6rTc6t0J3VrpzAMQlz95U
XGtSn3/w3sVIwP47EMXiRKacaFFA/poz9zBnyfLqYn1pTJshyqvyHupJeoQK7v3vRmkAPUqG85wu
qibbMJ9njYLv3lCFOn2y0CTA1g39/Tjztu/A+9PgC5os4KV7806+rtTbJ9BJVP0t1XsNFOUuGDoE
nza840FNmYEw9oDbRBR229OFbasGbvzh6L8SkjgUC0wUPa3TYUi3yXwZVUJMOyRxeBBhKs+H5LSc
nK9ZyagIoUMX1dCGRFv0+y2KeH9kZgmIJFgmXL0Y9LZw+8e4shfyXfDqRg+HZ5hFlPA/W1EWjDSv
vsFHSYYrv9bKMXrJ9jgulw0PAohNesUNim9rHowHe/0u39Coe4m65yvzsVCmcMRLK8S/yLWnL+KB
IRT0ubK9tttpn+UzI3Shc3wYnp3eLy1hoHokhafJII1eRzMAW4Uv3qnRAmd2410qH8yY0c9XNTPe
6J7+snqqvegsoPqWBWDtMeqGX6FEvRV7crWIkNkmVq28krWiS3zg44n4Ji4ce+Lzf1VYPHYZo+Ld
xQycaOB2X0cnaGD36Fa/EMo819FSRsVc+gLS/J+++9rXoewqwl76TWv2fNkpPxxgmTQEBEHcAMEZ
2LPKVSntpNlnUF5Sm6Wub4v/jp59YEerdAAy6KfAUKbfdWFc4dL1xFWjY44Zh/VlJw+XdAc+u8DC
HCZjJeMn2+VnOca6HbgNOoJayosfYHyPAWzo7WFL9v44OqQsGMx5rag7nIfXX3vDGJ5AyBeHL7ER
+1apnie90IobTlDSsP+WRlHyPMzVucr3Hd+uE6KwPbOO6ImAhNzlOKRYQyus9GBeDnsI/MPhdetM
pH3sHbvffRKkOBTAW7X1TphrCVgsmi63zdRQXywyymGXhK6AzJebSpTtfcHy+egFJWyyDrZicKmh
oy6YVWAdz+JDk0Cd+37ge5jFbdeT5Re7oaZW8akfK3DK1BfYzyU7D16MZLvkHJW4TO2jEkYRsdM3
9dU8nJb6mfdJo0C02qy8Qgkq3YnKNg1M/Q1OcxqqnxNIoas8Ca+Cb+FaF5jeeLrk1RcaQ+EhAO6W
Nhnj2y2nmPM56ml0cAQS+q0k/MiuRYfEx65HeIqohboQplPxKI0U3j7ghUTNCUTDyF+250KiJtT7
8KmaS64BPiH/uC+SzlQlH4PKHl7LeCUNPAhEVnGAjUcWNvtxxoWnzKwXn2kxbi5IThq0BrKfaPA0
DfioyMnTe9imT1+5pi20eQ5kp63lpct/jI1h5NwYgseGmxelu3JIYu6dfYOYMVx0k/bc6MVLJ2kK
ZKBZACBXQQnBCd1unRgkvT3yIWI0JNxBwLRBJ3MU19+ZQTC/KrSOTlnEGfwpkO9Qyri4m/ZXR7X+
U0jbi49Z43eON2qw+0F35ECE68Zavh6uSesCLUF4t2EQ1URQ/XJLqarqCSPjeVLWT23cpLWiRrQ6
yXTqQkR6lsfYt/0zCW/ACof5C5401mNl2LZtAIuciJ0ByJ+rqF7WEaIgG24Mz8RTrTXSkOL5/Aeq
qy0luvmzol3y3qRfzjJtvZ5HTOorTkVBtfW23CmQ5U8ICu2rmuVm+v9BgGOQoKjj0HeGBO6A1GpW
EOs0wj1nDnW68cvxpZlfCJgui9yPDmvnwc17MzRFLn29Mzi+Fwfb3p+ORh6Hylz+QS2n0/cQYTy/
piCpq69zpMI+PII0SCXoACto+dHRb4Wag7CBBXYkDbhYjIB9CL/MMrwHYMaWIU+8JyxoHM3uq8RO
Qlzpje8gKHm5Sk9l0W6NFsdp716ObjsAqNxjW29tr28oQSNy/9Q1dzKMWP6YWvZbLhobrHqZ3BFC
uLOiRL1/wttMImCMiq56vPxLckQHohJManq+BxEE8NhykcU3bI8KerTOUJVWfTm+REcxRfQ18RUN
b9M/msCXUj5yUnVxJlByvliOhc9g2ZreNHsT5p8Y+fROwlIzwwvbxlo/41y+y6U405FTeh5YZcmn
1MrSPeIdtjbffJmoAZ2uEZ6QCrbmPQ1ZVl15G0pqjVzmynF4BuWK/qwwKEiy00bioT3lCJu9DK2w
090kxeFHp2Dq2GtMcBXzY4pB+8kSHK2zBqQyA2pvWjYTzzd0ZArZ8q2QWQ9txRQEUx8GPzqyy/s5
Vp0rPB6MKzwF+NM8qNFFfdIK++OjhEFK+1bQEHbITUrQmpDCe5TZCLIrTG67dTzYC32+jGtQXS8Z
pD632hA/Ewt4QyepLyV0garL/mJynJWrsVSwLO7Qtz0iHgeSy2NFKb/jxEVA6NX4vUkhEhzMzFPi
yg8iPuys21r5DczCYpYsG2JRi0apOoKJlU8UhTxuBwAVUkIBb4eAe5lHjgA1a9sUiBVvqMwSwar8
ZRFfdi65GXIkzgrI7RyfS4kt+Tz4B5CKGgoG3tv0itqv8DUWoj/8NIUJ1UGKJAgL0nn22513ZtWL
y3eiWxZ36vEgsby25X7+MBqmWu3yVkz/Uo56w587zwrHhvZznZiWi67hwkARrSNzuGZrxv7vkQnd
zeL23NGcf0AmSdZT9hRNXFxSfWLx3jTFtQ9Lh7UWntPO/EHvhUvYmiAEgskiGqC+d8nCDyyWuv5/
Qv5tLW+Y2LXjaYR5qgcrRhQ3Dgq/UnYcqlQVfAIzOsWhESBYds6jtc2vstVC/Fkuhi04qYNVK3lw
V8yzGQ9u1G7BW/xx+Y0Yng4Xzg8tzsfTC3l9wQTrlo7uuIRQd2u1sYD3hUGJNgtWVvD3OS44cnC/
7egBfbRgUtMcdWcJC9LSp2J3UDYuFgExRbLS6dG5JhihlU9EPt4iKhy30R0P+WmwiWHfWGcYDnCs
KBUVFjboEwIuVV49ej36OCLimUEz33sXkmLqWhAXIPVMkYwbClNnRfnXuOB/lYaY7iuZH8Sodxag
wfxAvk3dPVT0fGlj2x+i73NarCrb3SVuN1T2CtCMNuWoSJeB/Yb2F0GhPIEW9+tnVshCJdTW9JQ6
bzbRgXfBU/KE8nhuVqmuCQSwHhaejB3/w75S/9rp7N1VF8DG1Vu+rlCFxNzWi+YX14XH9kqs//nU
2/Wsb4Q143OTSsRF4vCw4bDNgUL6u/Go6fIG8teTNqeeBZqzJ1W1yfwUnPycKoFMGOpdvZpE/CI5
4I7S6D7iNWYl+4Ble/AMEZwoxWXIAxifWqodmQE/570KBl+Ip6pkZ4AIvhS6Xv2cOsztLFHLYupp
uUjBsfloNxcwTFw+tiYJ7L6Udrd+BlW+6sKORuu2pX80aYlwBLGNXjgogUFwBzJ39RePLxh2E6tv
Qk/VO8/njhwHKLvsDXXHxq1LyM7IMpUBwXy9xEGhN4bRJDs0Z8CvIkx2qG4ArFbmuXOMRmbi8pU3
1e8cbTVioB5KPDVB6KIcAN8fXbOee1MMJO73EgHFKRF4VLTu77IMGYL9TEzK0brST8i9645bJO6k
Dqa9WTTad3u6XNLyvnfMocCB7OJfR4HEfMvrGhjKtliF8mNmTPi0esZa7UfXOZ5k/LX7mqYSc+pB
UymibaVTUE64GUt+eohj8TtYnyz0Ehr88FpobymXd/f0/w5uCXyx/C6GpMb9CwvBmxwEzYrkvFRq
leNy8Y2YF439y+YBZKcFlqBHPezE+39EK3d5KvCSZAF32UvCfOvLlHezRU/gX8UPojiiwb8DYXMS
82IdO6lCkx/SGIj+a04iR80uRPXby+BS7SbMjt1vKOMqiKfiTRrGbJ4Bt1OnWle8WAFVybLwOIl1
HcBCVo2JLdN7+hYIiWPe8SZKS3G3NyGRcaBR9buFbWIfcdceRt3fC9Ab5gMP4oGtrk88fp70YzHo
rR/nj9vNaALLhpg4Cl9amt0CUsRW13ss/GHuXqraIh4x3ZnvSv1xybNhyMCQYz0zJbcnxGrIyDuu
4DIp+KEqY1R+D2O2DxLTAgqTzKlXx3Wriz2QVbaEYuWx7GKMuHIGgSt1PnfUXZVt+ayI1qyX7u2N
/gYNl9zLAztYBUMHcFdBT85s2jeecNgHngzBsyuEYEw+E5qQMXzaemB5HjBIHjkHmk5ksuL/65Ei
cMhzJFqbwLVH1B/nag/7KICQ39ozUT6zAPyRKLSOwElyL5HncQTvzDjVaNsbsc0lirXlHUaLbj8e
vijRNaZcfn074nvInyXs5AijVl4B9xmO8q3r5ECs2uRgVz2EJUDUrHEXaeiSaMcku+hLnmQ17ph+
arTmj9PTHZ5nFT++PnJ9dNc3pEc/sZuKOo0H+qjAX4taWS1gj29zASzoYYXFkEmWHg+ETxmUuw+Y
cRergA1wgWn9AgHpLbw91ZNTCUyuFUMxYm1jn2xQ3otTALWkoWo5YivFP6EemCtA79Z4P3OrinNH
BDYIFYFa1CXai4XgGZ6W6lSNkUkF++W4HPWPqa9TztfB7YdPTHdvOdWf4jRZ+82gdHKlL0xFKI9b
GS3+pYMZkm1B5P5/kc7bqE1IvPJWYegMzoQvi7bGGVlg/FZL9JvuRsze2I8cOAwsit++Wr6I//Bk
BCCFZwW8/CBhS+PM9bY6Tows5EtCMWkvS/RDae1AE00Rj9HltblCrzgsUfxcVaZWkOQzwQkpJ9im
3gzDgkeXINRiHm2IJtH9RIcT6+Kux97LxA7rgDYHunoQhH3NikIsi5UP0n2BsvzDX/Jpgye18YYX
yCdZz6S2JoUsGCMrX5NV610yOCVZ9n+k3oVkF8kbhOHvs5iNW5Gdv1BnIjZFNG+Den9F6onUNF7P
EtB3+PmYWOdVzgPQ+9XIH9iKcrF04C6abCOMv64uJUdtkxsP65q2Y9ysBxKzwfdJgrQTkpEmD5hC
PKtIlwvm9yf09BmRw74CrT+8YOTcWrGycGgfnqsGk10h7g6ePugE3En4Mcv49sckfBI/qvu0PaVW
C+DyyszJjMUjkI8yF3RfKrVvtFI0E3Cabllw7Q45Ylm4JXuHYXCOEfnXBu6h4o8l6q2KddSoRkFQ
5JYBSLFxpB70aE1CPCkoVdIOXd3DDT/uAnBg4ta+q/7IeC7vYErFdytZHK2apvifvyrCyYJbfbOR
XSJwFbVPlGM6IycbKSDwwIfMueNp9LnF0azjvBOZVS9wJVLoAlHvLRkK+MKPQ2V3mCTNnAKfzo1k
erAsYX3RaPb7xFQCJVRzKggf0gtilSiRSRs2lSGgKJNLRoEHPh4IFsY1DFze8/6jAgn8qjPEAg8h
WI3VYd465v6C1rYX+t260kwJd7YcJMnlKndUq9KNvUah8FVNVlFfOjs9K7/iCEKYGLuBs4UZ9/XE
vdrUp1Y0NMwKK3emKH0juYy3pgNMhVc57nMxEZp9VzRsW9fCqViflUShYsknAQFCZACxz6N6RPbM
xNpgnOkiRjnTIbFXzKv3DNREj0V3qMEyUJww3mfiCohoNWAdmrZTRYSzEoj/bWcmBalH1WkEp5iy
WpjUgZ38tUGtloq9P5a/j7PQqCYqQQUS/ry3oPpxi+J9C/FqYZYggBI3sV0Ib84LH6pvo8tWLCH2
p9NnA+EZRGPTIybTzADb9AalCmj6vMESBapC+Rnd8v4RvU9eqna0lzI/wNeGXjzxVkS9Rit3pzNr
0mr/4bE+qt925YLaFIwlOIvix3877leGfk6yGbgo9apUlo1KiDMUcw4BCVD7UuhfythLDdLhu0Xs
FRjmIjkVKOUWYO4IVpLxt8ffc3AERQAo3z5myq9V3zKSnlLDsoXhk/zrr+DFfuzO7jFD+xQtMMkx
0ahCj2U0rQGM/D7mCbQAIWf7vA9V6B2SNByQ7VRWIIurFtah2aHNZ65KUIgj73tF715KKKH89Ryj
5IKTTuMYNFXMX7WUSQszjC6AuCkdTw7pegVJ+Xq6AhCuyW3Iz81GyuxowMyJBPKtMj9NBeUx7oyC
ZJEh17y8HdJwtioElYbCTKW76watkgr58PhNTU+YsVTefWek89Ox4tT/YyA2J9vv5nIZX+/Ef+WY
LrFBtlapPj+H6dcpJIQYpLcR2AKkPydhN8t4vKyZhWvul2KllKYl1IS+7lWicXlVaGslC3BBWZxN
/PO2+hpD7XSh7Xga8D340O0ox6kJ/Mw+FIZbqb2rPDACRDyZ/aBuOPOGUWodcswMDs9sIN/mt1Y4
U5l5rAfi0nSBbKvBuEux/LnAYGODvR9dbbkErgc6ja1f0vbeD7D2aHidNUwwDOfWVc5zAPXj/Daw
kb/+4fis64n8Eue73wqwzG8kBJq00m2Ri6T0LzdfBK68KWlPB81WsfLjc+Tnyz8IULc9vwUI3t1U
YAx5zzDgD56KkKade1w6kEbefKaJ3S/T8PGcvq1ULNVA7kxQVPzPLdtVTLnJDuCUce4dOE6IJAI0
UQwJiIzCEmiRyasvsruv2O8G9sIg0UTxNdlafumw0A+7h/EI+jfKJZJXdRIYR84xXUgzijXPWLGY
0SCTmj8a9PaDWg70DsOfv2nbPlr6d5OUs6k+BFdSVEN0VEU2UD71WfuixHOcXylH1AzPKKVvjxE1
TJ/1cek+QKLSqs5vDeo0iS8A6Ptm3Z2Fz5esivtlpHH1NSBSfe7AbdmK3+bKnYp34gIcHjqgoPO6
VFD1jhUKjmrCaTKBg5mEbsshxINqr0RWXM/0IvunsQQR10AlIo6v04FRxroCXba94oZQPqYEZjT7
179cg0JXx6P2WAY3dCp5wp0cKqulK/K9NZvK0g226YtVFsrgeccNENPjul5oxJwxdHTADmuF2iBJ
zIl3wZucI+aheBTNs407Y71yoAlH6ccgh1oTPJNwYmLO4Lego2DMKKSjcmmtgaa0pL85rRqrsent
AKfTpHUf6dOUjI4poYgnNIE+QDtrH54su8VpVI6H/rP92FXeBpD8ZEVm10zqIk++S+b5r4CoZB1k
syN3Hx4zpG4H7DMFOJw7DrUTgCVzXysSpJmDp9zSIQdADidXP7CxASqz9qqBWd/4sV2obYd/avWV
HFqKdIERv8yMkLvDm+mqv5u3tJP7lk15HjFTJQPp68ltcRwlF5y+/LHofrTofvoWogl9M3STnuH3
pqEVnxjAqZhjapWMiH0IpO4PtQd2UlxK+y/2tn1v7c/nAup/3iSHW4mxnTWQtghyj5emHb2ireTy
K7+AmOO5QB0oaUhyvhj4cZYQvxnktRFgqSctI+5lIB7wilyfHuBJEkyw8LjECrZ51LOO7XxSoThv
o2mLrQ0OifTKiBO+GLeJx3y+MvxSNVZT9BsMiwO7/x8UQZz1vcgeQfIRNQ0+7QYiLVyJqje73QFA
VlQPX6Ay2B3IMif8woN2dwXvJoE0kzfRN3Un1pVLSeDIAsYnCWR/i4aqmMrjxmqp8l9ns8MTwK5N
1ge4GIkvTy+u4mDQbMwXp3Lcyk2h+0t45fVD7+CmBwmKBocf06xSb4gCWYEqOiF+2ZJ7Fa9E8YRJ
OIll0WpgHqmKX+GqGrULtEqwSx7n/+iYwacFp/Z/mmaY2ZHduU5YXARrtbX6THIcY4ICJmb218kj
vPVW3uG2zcWikYE56kNhDJfsSVqbBUEumWfOsoWx7a/pB6yxlaKlALssGcBoHnDWGcxWpgM7ZRfT
2JfMU3B5OBd0s3+Rb+fHgr3dcc/uHP/I6N3FQOch7ZxSQb4Jt4GPj9nMFcax11WIxpse0G7wofjV
z7MXHoYKy21zSadO0Y4EfTNgWkciZxdPJ8HH8MX7Y0CM2mLlh20mGNHN5tb2eoWrd7fEV+lRbovX
KSXy8b41xq3B9yk5hI+OTGMmdj8x3i6eTdsXXQ3aLuhchjZPBBRrqb1maggwvhnaxRROm6dGW5CP
KAXIQ36knubDMdH14HO3b9Jg4fDvjpfU/CQ/bLIdbsVd+WhBI1jHsK4nxwwaesgzgg2ZoW65po4P
fatDKVrd0TN2zuiWkhBEYIlLXywsirDkC0030wkwQkyihXweXnlK8WA1cd+3ltiHibJQ4DQgFbPC
6rcJ9EL3a2eLtVqIc6Q+mdXQRqptOCBHSJXZXBr+G1WsbI6KKzsSfR6ysDoRScof8eMolnpLMWPC
FtCvEBHNH3oe6I7hMtTwQ9hbvu9OZwQb6ciBk5V2Of9r+hrrbte+Qn+AUCxSCIq72X+S2kahfbV6
SytrYh2IoLjsGR8rp0rAQggOoYYdNRAn6aYJP3Y+9xaG6HrdFUJxTmOitBANMAfNt0d8lmlPJFwR
4OZdEeQuj72J4bpRG5SGrIgczg6YEA+nqBJV2bSpqd1V40pPi2itKQgN/StJu7fFTJVED0hcOZmT
sQ/YYJFbhceyckMNeOk9L7qjuzgH9Z1F+8PtoSxZS20SxyrZ5xeo8Ln7hmlDAnd2BCrOpFs8rzOk
cTqMfMMqTaxM8JPqkrRqBozn8Uc2vv5J7Q9F2TgJc/Pj1b6yL7IE0wsim5AWva23EcZEWc0l++oj
zic1BeUjzmHbRwunNbc9Y8KE97eMYv/5l7V27bmWiNN8UAzriRui9RjBty8Bh/Ohx1RmQ4PclJxz
KaC9hIE6oiwuuNcGWckVVX0ggZogli9MBhO2wvCPtLItKvR1kminEXqFa1BdJLxhzJZICdOc878m
Urw8LY1s1YWZ+cCLA4urR1tl5arvtRv/l9bg7bxMKA5Hp2gbUac/yW8RloMWg3Ce6pQCnp3Jne9F
VUk/PM26FNeAZbcH1cYLq9RoNr34xQ6yMEqNEsVMDPjpOs43/vlo7odD5HnBOKC1jTHNhypzxjAv
yr0JrX2e30Jk8u9qUqSvtdOOMnKyUXd3P+SyLyygvLoAygnroneoGnh5ips7fuzzkIpTZvyieqsg
7Yh7s98GmTDRKVxsNrCjXwq0tZFofK3tXpriNcovIQwU4Okopfh8aPySgJbeOMoFZbwgOwXQhZpo
w8K9xTiKRlurZKzrcq3P2QpQcIFMT3sHE2J+EDAHinCnpY3OGwtWvKHDMnPKhieSLCsBO4DVZEi+
BWhVlER5uwWVAijx5HOZ85DGyak0RbbdsO/rPuyUpUMo9yw19/RJqiEuu3vMYdUA07/Nrw+Nu3or
GGryKlw+DzFf3lQY6WE+JPQaSYed9p7enwW7k6GHg26GARrqRckUx/f905bmxgFBSzYE1LFGCg/9
VIa/hdx6gp6GqBZyH4wFowOPykNZKho2UTogEX9Gh+Gg0JIrsSADFPAVYW7mFuVpflUW4iH3gQJp
ayuHf1sS/wafy5GgqnmKEpv/m+Kd6p+RJJRPy1KJbbNbZJtunktD87IL+eIm4NMGgC4OljPJrKEp
3YnmHORNOBiF1yHXZCraG79vbWzMUnSvwlQsBF3tqvESkFvZy2gSixRT5YFyhYNnMRUDTarTgP9Q
8PJ+OyZJFS2InOljryvN7ELgJ1y2MJv7YNVJCLgDjd8wLZxLmLnFPThzw8HanADxOB12sKbTDGqj
QC+Oda19YcN/3f3fHxRyQO49PTgRGBSxoDJABfWSX9mLOG6Tbl9hViWMrbA0/AjCg1NuNb4EMiII
/rmF4FlyXuhp5pq9jaEDze9IBjRVgdi4goF7iXUaJqyXPG1absq0Sne3TESI7xNSXD28LLjuJNCi
zFxYvbvaXDZoektnm8gkEPQF9fDzf/Nd18jgRjCfsB4jXwJWqs74cOo28t95A32XG/TekTQQPa9U
H9bimOG55mCZSICQdUPGP5TNXVlZ0uMv15c4Eq26S+UmX9J/UqYfQmNGxyYsVzvqt7LC5x6uJwzH
t50dCAM8NpPysdXM2qoHgWERw+wyd3w9bGkZSq15QDGjlExyCQErAPcQ9QBR90t4iRQpMjEk6Sd2
Nq5V3Eb7QLQ+8Guk61wPawL6qo0Kll+6HbW3FSkZBNkXqo+1KD68bEMFfVkd3T7DarGajmv1xPq8
tIQbX4V1c2IQOaWfSdKkElsTyR3zgxW6vVuUE5tH+tlj1smHTFH7+nGHUxdJ94Y9z5F2hPut6Fmb
fVz7eUIXO+omvPkS/9Bu/NEe9ryHK52QeVz9O2F3xAiGaaL24H7qtkfoGZq1Fj5rYzvk/dzjcvrI
HIN9XfDQZxBlwaJkdvgqxmnze1cXBLH/wcz3ioa3Q3L+KybjrpUteotOX62S5jlW+F80QAyTE9Df
ONCl73jgSOl2O9eaelDHLr8pMGpcS4F3pUYRifUSPUk1nEANzh5QP+Ncm7CoampbSigs71fuq1D/
Sxr47xvr5tBYzAOW+vdqcPnH1SaH/EpNsE3FULS5+1z034YmDHk0GlA6M+UdMJljEGIl1kQ4VV39
KcCau8YMOzm/Pr8VSeVVhPGU9SmyFvwfEVc7h3A6i5fUxPheTm/75MnOVAzYhpemsFFE9ZT3W6g/
YpaHMOR4QibGOudsTrPw385aoTETZJcuByX6xLxgmK6YP//yiFDeGQb9WUTgCFB/Vh7J5NF+8H9x
iPTToMTqM/mw2n3ox2SldakUMfDBuBEbktEpMpGcWiwjmg6hkn7fxiYJF+5SWBg8IGqJzBkka4Aa
veR/2ZypiiHm0MqBp8BIqQ+YDHM96Atw6ZD76Y1zB3jvDAgqRlLIr1z5q4zNGO2Teuf77p8akfEE
2lDexvJEwuCF1u6xpkuiB6Pnm8sFlN8HF4t4y3E5a77+Z6nTXStEIE9R0SUDV+0z2gnzvhrC8kd9
PMv6SsKosJJn+gz3mhiDTyS1h0Ww/SO1nRLJemWYcjZ0TZEKslCICepbSuU/gJFb2wtEd60dlJm0
GxiO69ouTXjXZShZbq7YUMqtsFytQ9s3tRgsD4QfSvakhfrxtnJ47tWAsbeIrLwYemYr+bAFhGwm
pLgRHElD4tkpDKOMYDT1eE8mAkGb2VXHwCRofQNt8vv5xMyiDyyFqLX4MmeO61E9XELUEdGGIFA/
6AeAZvqcyibrhu3apgKEaIQHP0n91XxYbe8beXgZ+VMUEkO4QY8p6HTxVO7oKVi/oJbI5MSPVfcJ
NzM2Ys0E1p6kcghQRNutoN7fxmjRaW0sn1W2qqJc/G8NfihEBLi76N+Kl5K2TNBi/XKuEeBUBDFE
UHx8UKvrh4g2Q2usdCVKzn/LEuEPDdkr0zAhF6IEsxi4f72rxCTDmCA9Yz20fauXnFuqIQdUItmi
+xkR18eERYtkui+OrzvUsxoTlKx+wXSweJ+GsNqPSrqlNAXr3rF8GYt52I2nXxs5/ZshT64Ydlnx
G+N/1SDxu1YgkF32aFVsdGuzUTXyYzxVOVDqGvGhlUvcLZb13EIt1I1Broof7VTQtpRScUxqElQJ
8cq4rWirb9y59K8Hhw2dVxML8OTPKanAeOoVZKqqV3Q9errzlyi/fU+Kqb78m9aCUmlx/hsZpP0L
ul1NYbidFWmkgXz6QVWz71tqfzJFmD9B3fRwi8mhRFbA4T74IQ6horuRezQ8WraYNGp6qWNM0DgX
/rp4tfYAantX8coU/wlbA1RZaqEbQgR6d61YZvjZbPhEcJBnlTygcIWlmzudPyjf7gLR7ebU1jZg
w02mxyfAKcfnTt9z8tF5klRH1bHiIzQkOa1N8URey6Bpwe/8dJtiSuGT15dPVokM+zWpglqAh1Mh
db8/jl7XjXPVxH4r0ESICBIl7MfJJwpSJl1mVHDj/L8I35A7dNSW16PayA/cxWT7J2MDDd97k1yk
v6xV7FtK7QeNFzHeoL2mO1ODO0VcqGMDjV4N6Y9VSqVBDj+syXvQJKudZL48FAi1/XanSCqOVOg6
m6zwWiF5fKUrcflQP8iJpx+Kc7mR8ys2gYq8u0jRcoI1naXzifrHXebkSK1babGyFinBnG4SUl8l
7C+vJFf/WCdVIftZjcs2Y/NMgsWYO7ueZ1i4HK+7Sja+7A0pP6C94LiXi1T8j9i6/q9YPQ4zyiVl
Ldcv9cPRZiyPDoQaPAQW+j8oAOfbGnfnc7t2UWlBkfBaaseGoxguz4NZjBa5gfo4kwHyH4024qTs
C17secLYZV5FZgR30B2BHdytUhBfsgen0w3FGSoXIWyBecp1SOIG5gymUsV1MvABUga1bWRaU+b2
v8duT9Me2wGsOS6J/oKrVJc8PdBCKcil3MYpzjHFocdR6uHbsMktSj+SRZjCxIkyq+zoId5Z/uoh
/F+lhsVjJ7k5TY35XTd/QNQFZeVq8uYNqQmn8SMAxm9XJuSNMpAYCdYBT0jMsrN9eNv/HuGhswIz
aGW+BIEMrlpLFbBmQP6u0JmVzZtjv+G7vLBR1KNTaRPN13vQ8H4PqFLarMrTjc2aOR3dVW9xcAnn
l1zKqDbF7lnZBegZ14GpPZdZ4O5XVqyKTXK7S5NvwHqTp4RqmocckDU5h7FFSGdMG6eVgNunlbE5
flhVEX8AIFyyitvvD1f9ezhWJD2xmFvhzoRRjTjDiDoTog69u9ovgXk4haORorfC9tFUDMrvNj04
+vOTCE9+mrGfgv3WMT3QzQ5iN9MWel1U2rlvQ8DD1zJC/KYBmeoB4fKngKNTewpAcKFdrnGloJ71
cgqMWOZVL9Fwd+KY6pZBagvT1RS5c0tjXsWhDiPPxLfS1YmYSj56vnjnRFox/Hv7RRgivDI2AX5h
/oJma8r2fIyhH/u76t0261eyn27lmZWpPEuzTJOX/lNQMa3ECUHx77ixd7nF9cw/VkXT8yyaUhAx
Z+YYwV9KkNB+856Bqg2vnAz+iA4mdB2aq/ueKyjjm15HkD0gSNSf/Owwi2GISv12lSJwH0kUUYkW
0vm2VIQfYlfA83Yu2DlJmf5ZkVZ5lB6VlGbKWPUKWNwWBjdlu1i30X/Mc0vlewd3AuXAAmHjZO4I
281aliHglwlr77bG3u8/ezhkMDxeZEdoSYQe0QMORjjkxtTdVPfZxOBJeoW7AdijG9INsfLoPX5I
WAKuc009EWvEeokvtQFl5KCAJhcT+SBuSpVKofwDA7wDiAF7laSI4iKd+ntM8Byjz3RTsrdhMgeq
PLwdf0myPcO5uPBXyC7ynE4yojoliZQ1llm4J0GA+IXVaYdj8z5upiYz35TV754ibKf0wmX7JMhC
N2pZswMbRYXthlyG85IQURHew++R7/La2ZoU2Mt9Sme/Rcn++CVpBTNMNC5urz5tVrFERlqgr6c+
N4fYAV7a7x8i5ZdsIsl1OBXetqWVQlyOdfFjnwWTU7IC3/NfZWoiSMKmSwyCSiLRC6tx/MFvwt5M
7HPtAdF96yNUlXciyO1I1W5fCsON1UdSHjkzMtBUbK+THNebXUbkVIUmxNvHHaSw8RRrVw32Ancd
EzkPByna8dbWf/2lp3lXznJOfkul2ecQ5n/MQCajhzQ3cFUwYSd32nCd+VCEkg9odSCjqR+xeztN
3bAS0u9j5NT+mqhlaz6mqwEITlti3Y70aof319CAB06vcwxSNCfyK+O+zffveXPRhDqF3kk2rWs1
zmNYIF0Vtyr4j4jIHUknn+N5YR/VmjH3ADihQ356+G8jkhCTKklCkOM2ESpHMRkFUefSyzgVk7Yc
rba+NvQujuq6j9Gqstp+mBL6JLFYjzC+tm2sLd4kqLK5qhlnX3YsuBdPTz4YVluIBvDYw/1UZCtR
JwktaFC5cfPzuzXOuXtgdB87e6nXmef7UZv5kGftAtbYzW+dd8ej+dN5BNvJTsiZLFVyzMXEoQja
8CEuiHxIomVKMYPKw2I8FHq7a8CnLegcwrQZj7+zQfFnGXew0Kv4CfXo6GB2o44Fw1m4htdRALFk
6Ra1jlqbuhL3PLk//6SKEr7yePpnwORfKnup+5PcePegefrcBHmf3DTMHtKYT0UsGJeoccMM6PI2
rS6+WqL7Gwryulhc0L5NwwAsdhoYFNGNXCgmQe81ecBX9yPwhUbkYEBhh9ouUlV5Gzf25Cv5ESfU
KhmG1i32Vk75MnNu96V9wMBY0XGqarpV3mPrOw3lxE+UUfPW1qfRbGf1W4R6Ufla7aWPMN2GzuLb
vY6ukSdqLcyj6/1XXhX3M/3Wk5pe+p4lE31+SbqPn0CgmOUsRl71CuTgI+edaEYlB/5KVIGpPqx6
089wIggW0xAvJrlDlpChJ0BPUDCLvTNvPGwHM12xjDGVyGKlio7fY3qDBOt5BX1DX6jDFLyhn6az
18df/+Sn4Id4lhFICqjh6eDfVMEJEVhW1Krk3qz3qQ3Sp0zb+IXk6xwsfcabshTRvc7GZ4d3hnaf
xH8MBh2IO6afQwAYzJjfWSHIQkvhpEuYSv8nD9OF09/temgOvK5dZdyVkc0Dbvyy8PSNJTpav6h3
2qgyiu3pWMei3q4CNYS8DwhwQgod8tdaAeQrweAUNdAu2ItQo2egX1kzKN24joP8SGRYzFiQF3np
eCeO/9DxbK37gRWlpbZgK04bU3ZrjtrkyMQkdWKsP5Y3Rs4vyKzvDMfgZ7/EJLWaaimlQz03kp7A
BtYzW4gMn1cF8q9RqNWOAsX4EyyaJ2S9YZeMWbxRzuXylY17G9zgwPOzdNQhD9nf8MPHg5vwxzaw
pbkYYcZFyeYnSj0DHt+ZIve3aFe09EpFNPlAtK06WireaIIHhr0RoZSWvqQpZHs9joFj8uQt3h9j
NjEwDTdYuBvGEFMabjgI1mM9fLIxw1eBuIBZGbJT1iDoBIC4ek2CWx1ke0UAwBgxEaH1qOn0Qk1q
X3um/NkmLJWYAhltxLPqqBaIFfVG3SVpxEbqdJ83apO8zAHqEmSxSB+/BfXKuToMDmYGc9+tg2hN
wEIB7NsYMgbpNmU/fFpeM2p30f6O6k5ov83eWcYilQLG01N6XTRPrCdZ2PSr2EyzntPYYb8TfvHg
E5wv20z4ayeDmp2/CzchxxiltYMLU6TQ3VCLaLt/wf5PKnhafX9Ai0KpoB0acIdU1StmTs8/VqqJ
b7jqvX3B89ifwGrU7BA+gUpD/2CJYZ06ou1W/PxEkuzTM4hEwo8Oi5vTjWCd2MLSOVSI3Ft6FnLY
Md1YvngFW8W476tj391vMAySvkywqpAZ0QflRv2Cz3+Wwamqi3qNikIP8k6S9/QF32wRLaQ+NYlm
exQH8m6nEUCPC7Z/zFz4Vvy6/Nl9hm1EmaAVTw4Wp37NhgtnhdTCXh6peX31WpcrDnxtK+yjRGFi
mH4h5otGCHMhU7uC3XNDC6ia0gu0IhJVHYQnT5aov6YZkGSp7Fw7r8kPjxeuPzjw8/6N0IY22ClL
m9ckIZENFxN6R20b2fe/+ihTVhvXLHCZm6K9GQhjBuaskKlEjFgJkFUVSMZrmooCiqtdnTBHsaPO
UskTtn+qO7gYdCQWckDkOA9EnVKJ+hAOvF5ZKVp2sbxD7CM9T4GSyHfhiphchYNcSPR5T7TvallL
/19zOLDLEVMxKplW5rOao/HEsB+PcvZmIpQsKWVp4uB72Uurxfr4afHsJ+7DmHV5D+4OYbSXKL1x
XafVH34mUZtygrpl/5Akb/NcMserjNZRZzXDj1U7omjCdzw1Ki1Lk6cJXnGGptjUPiQlKgbJEhOL
rp7+WIQuRNgDBEZyb+890ivaiEyzZAUniHWisFfXBaHoVSNP7HOhBQuiamff2TnU3+IIEokSb1ag
oiMlEYNconU4xYYhdzjcwLlECDT9jXZFiOHvl9X03KNKx9FGzuQGUcEE8YqA4Bi7nWoPZz2qMgUj
/NAonaC8FbadNmRLF4XXa1fstBEQ8Czgief/lMCEbYLrJiFidkUMK4i9M9v45dkYaMjGmrnOXSBH
lNN23BENLmrJ8aT1FbPFtwzRPwzPcXpgzurE6l4WUoQw19WUbgG/Yx5Zv85LgWFl5zR0uKxw561c
1+LBUPFMZtoN8H6oQ1HV4EhiQhINmfr/iHBMnbxfaUXS6hHD4LnW1AWnYUyjxaFAQkFAcDEEK5CO
2g2nQivr2oYBrLGGxomFA12w+v8he+k78/GlXwG+tpHCFhPFowEAMCL7bbHLO5PtiilAjO/FUdi3
OVQWebluG0BVs41d2GR4iVc47dmalx2jq1AQvrvFMPVrhEAlWpX7s5+CFO6MtWi80CqkXukb5e/R
9n0Y4T2Bphe3eC6bwF4YFPRwuW5E1wjg87k3S691UKNGlWVVjCq5R0YKbG9OJPH8ajQd2xDZZSc8
6isU3cn9h1L9h4s0+Pqt+RZf5TMmGV9DLR7kQClLkWeP57WhNdV+mLLEBFB4X/mykqtp7wdIoWDJ
qk6iW+eyBqSADn635fIM++XwjxTGMmBgV6HYrGtc2rVQB7/UakODtr9nWRQUoTpZ5nILr9UqLlaI
1dVO4++bRYM50pbzPGulixi7GOWXs+cUboaJ4lqTlh+Yx59Mrl3GGyYrYsa3oJy2qjJnkuurBlyK
yRvpyu6+wZP6X0A2yXOV3NBlSYHKT60JZl+RMMmCx9ZMyjb0IB+tNvGcJJu6SiDfjrQJWFWxNlSZ
MVUcCXg5shJslgsLIDdNk7i4zkCZ5eK/5eQ9ZBOgPrS7k2CCblztybhMvratzAHy9QG9RSZHGf43
0wolkvbAd8+Zjg3XzPsavIsJwUh0sWW4/sqKdQpOB1gM4JPGLfIdPbYXMhQ0YC8yDPeC5o02UUHx
3uikiNuKAau0C33MN1uOkyzBfDYwR5O8iV6Ss3KRJ7KduQSm1CoK6w0WcIheWRSRmgoD7BG7321K
pTcp6E7paySe6kji7b2Emp4qM8dyC4i/Wio36pUC8Ii1POt73Uz3oxl2Wsy1s7HO2OmU5ZtnrnnZ
/JB5cwWIjx38V6mEyuvblmy2ht4+FffPK1IKb5qzg0Qy1eIcLuSVKt/1dqcFkrgVVAhIaURWqZSF
bVQF0OutNzhXIsAOnAniIvoo+dlpnP9Q0kLzf370aB2zCr6lzJevc+SSSQU7CQKE2UckdDCyPBeS
6sJ9RUurMYwlXTmhYA3UALtUDdHQiO5PbKahkePA73GGrrrqRjTuB8bCHJCP/XXYO62C46hGLvFM
Ky3h3xULLVsJeJ/IfSvcvP/hNend0AevOtfcdbgc/JDAFD6NtEVkl55FXihUZH5C/2DUAmsdMbB5
ElW6W6JYycBlf/BBa8sOtdRGWdSNcFYgqJUROu4bYUAoDCNm8rKZGavP2mNwSJCTwmblWHHNAl6D
qYBqjkCubjGP+/fci6rgGj0uDYz61H7G5IlERuUtvTiVk3WCl+6uFfE2IEJI3WpW/6vfB7V1NLTo
y1pXABZUs/EnlDdxnaQvEbIGk62zOyyVjhG2ehopywQJdJ0fUhRDKzMEQpR5av01vSTKql1Me4d3
G2CE+zLZoLp43KHD6PvsGxJxc5h/+Jm9Fdrel5XTQPqBX8r/c9i3vBskaHflBOET68E0NQEd/J4g
lOnPPSauNQ6vVsnHgEzDwc0dSAhGFp8y0u3ZI6lG+zFu7NyxNgmBvz4L9bVof+P93DoewqkGgDVy
CxakXDf2ExpM60YMFa1StSNoCLyaYW0rcgLOxk3nCjE8+mRypfvSqub6mmPJvaiqjHrY+9dkFsSi
kjkRPWZqjaYAAarDgepHgUvjseL443xxzQoSEWO34aA3ELnlDVcy9UwVfwhEU3QEi+MHGlk3Pmok
+z8rtt37HTNXnmtenFMgj1r8BNcOB9RYP0mJS6J46j5HMuoKcfaUWpyNWC5ZRMoLfafI5swwzpOQ
mbaGvu+1MubOnhkoLlL/XdRxseh3CmTDt0yi8nosW2WisJHyCO/pvEEAXVibxzA1KzAjOjLK2gNv
P5WvHnolDwIVsZmQOQs+2tBsnSWMucnlkb+CWY6i5M46GHwWA4caeNM4hVeRaEtFo1s1McnQRtYx
cgiJKQI6uOcBHFr9tiyPgE74Q7ucDLAGPqMTQTUqVoBWCa4G4DOdopNfcUbh51Yijp3keFvkTLWh
WKUHqNmN+UJdSApnx4v6grVgcVb5Pn6x3sR1R/78rmbQPBLNmjZDg4PmtOwQeGRmsnoGxzLY/Ra1
r8UF70KRcl7QIDKEWLtjW/4Jk/ChUsE1/CqTTHINxSOWdSkC084PjYbj7TvDQjNLOdZa/o2M5us2
5krkQ1052mWuiBl7HQK3z2Kw86DwzA/hPp1QQRsyh+zcLIkG1hjeqiqo/M2KOMEwppxKKI9G6jKj
X8OHn0gYEvH1kYuORWasrSggXNUAGSnfKu4eVF8aTv2mEy38bcZpRBNh365nZL3YseQDs7aYPipE
AEjYIMhXEefsNKoPawBQLhvfZ66KWsN0kfF1x3ag9HFibXzRxGozOl2J3ltzGIWAFst+4yJ2brOG
vJsrdwkjrS0ZzgKhfLQWBqMeXKqIfeXj2Ie2h8sl+Dq0kWM+3fdcWbQutiQOv+Wcu1oiwBcT3616
JJl/oQcnBeOwJg2NjQ3G2+g3J42EnoM+Vm2xalWQ2TvXT9e07av1re7bI3aMgGjnWgBdoF4ogIFa
M/K7mds9WtA95UiRSzp3h8B2ExQVKY+628P7PXTsbFf7XAwNp+w97bYCVj8vv1CEqrtiEhdjdH0Q
kCl0TP6oZobAKTpeRmvhfyeGHH44jtqVN6Q5yw6q84UUTbdMHCql+o8iYBy28dI5Xys5+jcAgduj
7rJMp5YnsuXBFPNUvAQNQNO+Nx1937h3PSRHROenwkviGlY/1ep5ZkSCxJRzoFNItDnoy+fg510H
U1NCnzKwSR2t0vKB85TttUvP0Hmz0apCFPaSam7sdjeLbELvici/drkrF7XWbjs7sTJcfYJXAS61
3DQPQwwcHxXkpm/WwJgiECVrN8Q9Jq83khv3gJSrpgUIjkr2AE8xBLvC/hct14CynQJcMjgqW5Wa
+uFg6YkGxRkke4RLypWfkZsIzRxdEnYJyXVsAMweSRUl+7ASN98gzAAW04OXklbm3WWYlt7EsY35
wj3BEY2CN34vNJirjyDVoN+IJztZ2v7fmriga7TuCl0SmPiZFX5PFdj0Kl6SWEQY6hVpSSC2xPbD
6xJvtcfhYYqyNlo83o8DoDwKmsj3d6EwevT7pfKPeCUBFw4V3oOu036AweEqQqf5fUY+jfmK3jA1
ILaDt91xrcN7vgjD7/UKxWicsiNWmfplXRTSnxFQvqjraMfULqsBZzxv8hsU7svSFDkx2X/UzDIm
YN/tfDOjSx1CDE5agkP/IH8FIJ+Ds0GZXKWl/tUcgZ8BowabKTNr7ho/jrrqdwGFc3gEQZ/2YPnv
XCpzjriJWm9UMIDImFK2Yt4NE32ka0N5qXUBijxxv7VnmspHLJvoIWs7IpfQK2EuWuTEYf7RiC1b
04BX4a0wX03IZD6IKCpwSPr5V9xhNSsl1KdPIO61c9Z8oAnRb6BLxCXbsjlkU/QEDnTsikd0x5We
syuw01SqVCXVns599Hm8JBSBPFAYyY+uMYKSfE1jcuJ9bF0vuwUvmwdONguaX+FKPYxUtkOsXOV+
HiNTLJZxFQMkPUAnZQyq6203kTkde0oZVHI5cRcIqVzWv4juEEC3fH0zYYAtCMDmJTSvpeJJ88OF
q9mk8Cjbkba8JbgNIuEwKXkfcibwBmnUlfWDzMkXhpOJrzIwQzUwjc/Cl+hh5Ttxl3xknkzJNbbv
hupNJhQxBBWv6BFe1q0u0W/InYIwdHUHD8hGfZ7Jylwm2QU0xVBJxx0QtF+BizcESSbCtfBuCasd
bZUdx/At1TjFUrjxEAkM+UKMKhbHo53vjB94iW9se4tqwQmIKcQrH9LPj652pjmRwrtUhqDyZoVn
rne4aY5O6sStJs68kJMuYIwU/qZZBOpYjTVbuGkj8+EvkF0JZcNe+YYMrUYgWNKss24FIib4KBLc
ORE3QdLd0hcHiSdVbUFmkYVX3asIM5JrE+8k0FgzKGoIRiZbeXlMLFOTFPvXJoz+hSwZQYves1/n
B0JNlw/qxJjbZoWonnPzS0XEoUuvmIKgD7t09ZEi4f5EQ0yYtfJ/E90waZ5z+YZIQZOQRFG99mI+
8A/htVDlbHNWL82s4jyeQ19/WrevQ5FpKRTBjnWqPjM4LTzgE72rjFQ8D16R7F0b4HQk0S2zxBBg
dIFQ/VOdk3/HeQAac5sc70NmM2T5JZB5Jy+USF4xasjIXyRAVcWg1YYEqw7kTysC6DCucPwXEh4H
d2iwdwZrpiRks8RahNpIOOmDjd45mavX6VWW/rAkOiGhy6KWXABFOPNsDPBl0Xeg84PMqZB6LeAw
KOWhccJcj/9unU/uL+8g0/8SWo8Yy1d3QqmWzap7yxexmVl/eJAP1SnBnw4mk3HmUpisoOjxddhl
TGBymQMU0UH9ix6gIVqPazkNTsQZklndsFcrUM6Tqk+xksnxrKt2zSCDzptSCsL8dU6sbPcu+Bt0
Bw/L6/uQwidxNrW3hHaPtyfRCWzjUiiwn1SGLaUXuEdpARiW6DEJ6sN4l7yFDPo3QjqrRoyNpEy+
jAPRMq21pQFmAUEcwJz0+eII6tiGH+nqQukR+px7S0qicQnr60XKm2hRg2umvGOpDQ7+NY1/rCqI
FPdXhlnh0ndGfCB+pIJiWRX769nN+gQ6UC7/PX7PKte/TnMGAsKWXgEqlBBhELoWZYYc9EDU9ahr
ToBwvlnihy8yNsi0qQIOULLxleCID/uP3VHXLxEVoXivtHadymuUuzTpaW31eOtqRcXUFwrD8TxH
iYZfjdFfXHGdGMpGY1339CmXVQE3RVwYMJobqICF8UWV0sI4j3jUQI9ZpGh0+UZW4WD4noTcbWWm
oEUB751JK46NCTHDEvhkI7thwXAXWFnLblgOz4s0KlgX8K1+NHQ6jbC8viiHZIJ7337BTawALPPz
0/4AAyMu9uiWBtq0Df7QcuCRiQloow2ZVq0uu/Z9A3KDwVzpw5fSHeAFZbSjNkkXusjXlFZQOetc
vxUAyeOxPK3k/9fXHaXKAhc+7kJ2cds4OpoGjeCyR142O0fYbs/aJps+wiDXLMZLFXKyGE2mkssG
V6+pGOKxHxZyHeTyRvhTNQk+juN7Z8E8lZGAnqSNBXYhMo4f6Wq+mVaq5+rDEyYZHPqknslLujbz
k4gyuk0pvwwBiBahL3Ll0hXYc4og10RIFrsIICavNgNpNE3MrXU04secInk6i/tN9x6YpwNKRXNb
EB6MeAb86XJcLJFcCT74caSg1ISay7htlQZhQCzu2HL5VbSS+E7NlCASzlBcEzuxsjQng1LKVWIn
2rKdA0Zp/x1arFLfCkQ0nfqgtWeUPb/QBst9FfAj1WKG2utxRt2xYwtoL2IMcNwfMymdjBChSKaU
KS5PNuewXS0T4+BybGCGvjuRBn3WaNfbwLrre/DqlS7Z6V7tGgS8vSUalO6+9BcpKdrWTMYUAP6y
8seoHXVAD6k6l3VE
`pragma protect end_protected
