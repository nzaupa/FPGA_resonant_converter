��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_��^pDR]&��>xJWB���<�ןh-����s��/ze�nri��rT��<�6�uEmV�y
L�nqR΀G�;|��u�(�L�Go�[�C���m�L�@y�e�瞢|pN��v�7C:p�O~�����G�/HįҸ�&ə���L������R�O]t�*�s���&B�0k;z���We����
���#2�ԍ}�<1|����iQ�8Q�:�\E���|o;�%Y㷪��f�_�ׅ���B�-W��d�h���7:EKF1�t=I��hQ��%�� �h��kA=y︕���u,�/�څ9q�k�i-�y	U'0��Ģ�y��ܽ�pU��'�b>m��K7��$�&�k�t�~M���f��ni�Y���j�pVI8-f_np� W�F,�%@��b�"�v
�V���nl�%ϟ�%��Hv(�.@Ag�K��ڻ��� �����E}�o=��.���v�@��`�ߐ �f@��u�Z��L׫9E��Yۍ�a<NTp�3;M��sX�
�i��M��m\�;W��{�Z��m��\-r�"W)�R
-�N	��P �\��d_�[�ǯǬyS���'�����T������Th���@pxO"x	h�7V:n���wŎ�{x��J_�k��p)�c��]j��O��M>L�wO����܀T`�?��������������q��&�	uH>�V����&6bW1���uzX�g�"6�c��g5�U�'rSR6�qE2[�V�9�gA�\)�>���J5��ɉ�h�z�JE�݈ޟ���u���4��>y�8��h��S����T�/�?E�?����M�>���N.����H�pߕ;�$�ŧ��d�ϋ���zW#�^^}U�����'[�_�`!��R���V�m�PsrX�/nWA��l�h�*��*γ6��.��Cq��:�=Rr�NT2#���Ȋ�-4DΈ��(����	������WFJ�^l&�/�3i;A�d�q��5ٹ)�B��6�ѥT��|��#y�C�/���y���bօ��\Sݢs�gI(������\���2���x�Ȱ�\�Ql�$�(��w.��uЃ�B�=#Y���=��}K9W���DZ�����m����U4��ĮG��ܑ�����4��_~�?�~yo 6��l��f�"�$}���T^W����TJM[�=s��C�zU����O�:�t��aP�DK�0�c�.Y-��|5����S�d�T�D���"V�	���ƉC������G�;'e����r�G�i3��8��A�:�r���~����lث�.LEo����fp���eT�0-4NH��^wtuHB�ݓ�0�).�����T?��x��;z5�C���뭪 �6#x~��ܴ�h������[���@=':����BX���,Q���c��|[Y���)��R�[s��̟ܵ@I��Ŝ���>bOs�n.zC��Y��cvF�s��z�[/0.V�J�Շ���X.���@l_�ν�nZ�g�.���J�\����p��&�ۉ�%[kb�4��{)B����M��R8y�r���y,���@�IDD�lRc�q)�i-�
o��2�Z�R�+�s+�3��x�_Z��B��*p�u��v���8R�x�N(3O���E9ݳr�}\����3���� ��l�:�vKI*#C0���X��a���9�i^yZ����wjxo�� �*d:�۟��GAdtR��܄҄������{���quf��Nf����j!R��1Y\uUu�&�=�����A�r�G1�f������>�c̃����-}����sB��B���n��ߥB%2�Py=���N���FRMu<R���-�s�%� �1,!���c�)�?)!ͨ�N�p��hSa�1�|��m��?x`�ƱQf�l���z+�Sz�֘)*yՏ���hess2�%�)9�%�"��0}��h(��v��GV�ʌ�S���Kp�c��]	���đ�+3"y�Q��^O��ݑa�~.π$%�L�X=qV+�J���r/���i���1�#m��ߏ.T�����u<�I�6��D��Pėz�H�s|�#���;�R����8�<�и�իQ�ij�1o�ç�
Ic����}բ����H�ON�Q���;��pUe�F۽��7�u�p;�a�a��Fi�������[(�Nq3qIQ�T:�ɾ��|�ꆵG�<��7|yS��yY�|~�Lk@��4k���3��!�]��
f3�6>�����+8�̤��x��}
�BluX�K����e���ߧ�T����=#A��PJ�7s摎���(�S�)��$�P��ji?ZZ_�_G�@8���>M��;��%�ތ�G���-��t�����<�	��N�w����ݻ�nɒ��B����e���NUS�LQ�Fh�	�����vd�y8ag�� �N��/B7��y=~ X�SE��r� UZ�c��m���97��^�x�oMZ:z���Y������,� Ov�j8��re��~M��pE����ɩn���lK�ٽXy�����*Lڍ�)����>��c�T�t��,<iJi>�5~�������i���Q1y[V�C�);�SYQ/�I��&�+���󕓱�[�F)k��Ǒ�,�'�%[曕:��� `������6����6�	W��b}�<�HI��{���o�&�HDd��s�D�0��"YZ�}������l 8ؚ[�.���6�ߵ�np���U�w�ߧ�&��/��@A�G��<��4S�b����G�t�+�2�g%˟C�T���:fQ=7�D�ڲ�w��څa�$���$�+�l�&}�P���Χ��w�l��~rq��e~�Ɠ3�׭�؏�u�9w�aʂ��,8g�S�`���������|b|��Yt��)��Z:�N�+���)��".�g� :4}jD`��cyJA� �le��*&#�eMk���a�/�?;Ǎ��Kt�ϭx>"/䵐ΐ<��� 5����\<�!Hh�S��`HW����PS|����\�{����P�^�:âW�T�'G;�*\���2�ߛ���"0h:\]���)������j�x��pƊ�_�P*0 J�=Ѧ�6�i�1�6�o���	�YhCx���o
j�&�_\�#�w�+5�]DG]^��ȗo�r����I�{�T��%c���� ���>k��Zx�����R�e!Ȃ馔{�U�$*�F������e��#���p�˧1Hδ���_2bs%	:�
ϸy.�>��(�s�HY6 '�w���A�d=j6* �D�#ݚG��Xn�������Ր�!Ўh�

���x0C�uu )@l3FX�u\~��T��N���;Eb�Kp��s�Νd!��ȵ*�v ���ߗ|J\O��:V� JJ[/o����I�ZHv�m�X_[0�]�覚6m����m_w�-�1�E~���m-z��G��c��Mՠ�`x�MUm�x#0"dH�,�}��lbb����s�w�.��j06Y�u����o�{]6y�}���:~��%��|ts�W���+[vI�,PQ���23���5����M����V��j^.rB�
�*'j$��^�3��}�����_ic+�� �ƈ�u�rmC/S7���sUX[:5��g��m�N�]=�w)��0թR�$�*>3O.O����JY%�ŗж����D�Ǽ�6�3:_[�,ˋhM)i��D��v�۱(e:~���&�x,�N�l�Oa5�����W�a>%��Ŏ�����>��(�)�%"T@�͓��5]�1-�J� fx�,�vh�'ߪ�m�.���L���#�c�Kw�r/xx�,b�c�}.���7�*��z��t�o��N�?]�yx�������~pѤ	��?�_O�m*�}�?c̥/ۛ�Ut�)�P�Rd��'W#'��֗�BX��ɀ?NdX��Г��9|�_TZ�|�k!�x��ɇ�m'����]zOkT͓���K.k@}�a!���4�ߎ8�_ca���;���T����0$d}U�nF�{��>BI�ð�j+$:�����M��ۨV%C�f����-΢�6E/�����Ry��K�}t�Ȭ�^�_����u�	5"X�t[����.<H�+��������ٽk^�L���ռ�a_���Ss����G�X��T"���=�r�D����l �4hd�0::>�R
H�j>�Ȑ�]a�6����j2�<��[e��)�W�#��}�4>!��c�-5�v�zc�b�%�*J.�6�g��mbQ��'v ��1J���ڵ���������h���m��w�;�),������v��lQA"�I$�!9��8���v�e���q�HhȰ)���,ے�q��� ���4���A���Va����'fW>Q��
[T���*G�����x��|���	`�d�X~��M�<��"���]f���y�d^e)u��7�a~�h��-�1j�6�j��������|3a����B�t�Z���ȴ9��T3�p��b/�`�&������`�b����wƝ,�)���.��ޥPzN�N�; ��Pi��z�b��� i LJ��	?0a�ZMT�a�zfW=�L�Z��eFP�v]����+Ѐ�Qj��鲡�.|�C�Ç��RX�U��\xo�h=��ZY)
g�+���Y��ڨ��=���L��oQ3�lW:�ɵ�����¸�+0���&��I'���е��4Rr����a�4�<�|��I�- ���2�u4{ݽF��W�"�Ʃ@�OV�D�B&T�_���@!<���׉���s�
 @�����E�J�,���x���a�)��}x�%�� �i�plv降�[,������d%��V���i!��`�#�o�7�!����wD*���\�������	�Ҩ�O_p�u�mK_�]EE�	)\��%�qf���+���[�-E$�>�e���y�;v��˸}��!�N�A4�<4.�&��9��V�N5��g���i]����["�"�j��hY��`H�<��/-ޱw�b2�-����N�c�+�Ǿ�֡�t�v�3*5�u0P�|���w�Hk�KW=8P_Ah��JY7���Ej����>� \��0"9x�9�B�R����NLmш��S�*���� @�NX�H����3W��u��1{h
����U-��Hǉ��g`�W���$� �5F-�o0��I�w�p��Л��x��lVV�f}f�����.<� �[<!.�:�y|F��y]�b�#O�\�ʥTn��J��RW�HX�š8�S��#R���ǹ�#��.�:k|�����Ǎ#�0U��dC�.�����6��Ǧ<����J-+���,���2�Q+�D�H_t������.����!�X m�_�K��
cg��r^�:�Fd����Y4��3�\c����`������/瞒��ϖU�9� #!f���d�M��l�o+6�s)T�����{Ӆ�)^��sSƌє�����|_�z���1���<���.�|��#�]~�H���Z��M�x>�� q��+���{w.���S~|2	@+�f��a��2���sn��֞��	X%.CǓ+�g}|�r���\P"|6���z�,QS+}[eh��Au���ζ�Y�5տ[X�8A#~���ʉb��%��C��L^�Z7��<8��s�I,�]q���DQ7�"�|�>�����Nu%TG�m����o�c������2����T?���2�3�EJU�;n�R�;:��'�)R���4�������ָ�a�A����v��� �������i�O���;U�5�~�YS�xR{����s�ChL��5�^���d����8^X�(Xa���@���D�Qr�?0����T�J�)s6�U�G���w�H��3Yx�-�o4��5���t��6z���ϼ��V�w�� �X�vpr���'iӖ��2��@�u{���λ=�u]���&�Q�W}JN��U�R��\�_5���1����!��IUc�I�t�E_]�a.�����g�	-	��{�����y�"bMۆ�%x��Y	1�'��+�l�ԧ��HH��6��i���
�.D.�TFID����;B��foW#�~��Z����x�+n���UU �G�s�6�{������9����L�����-+0����L�a��3��5ʟ%�_�+��/�>�	"��S|ߡ�(���`����K���T)רm_F�mF����1X��;�F�.������C��2�S/��O�PϷT6�^ǝk�	���izRfE<���䙗�%��:��cFA�8$-1�GӉ�\����%!��%B�6oaJ�B�v�c�Za�t�����߰FqTZ���lD���L��7s�LoȓhTC�ϯ�6<�Q4to9�&{zI|^����!J(�F4�U�3+���nV�vnf�p6Z����C]�!V�j�N|L������z'�	�p�f��JY���3�MO����_��ϵ�@Z��f��e�����VC�E�~'ZΌӭ��Zm�6����F^@�K��U\�ӓA��mֱ�t-Ց��U�][H��A�X���9���a|ep�`<}�����ژ�J �c��q��M�җ0�}5b�z��ЧQ��nǖ���L���������^8_� �B�a�c+?>�@���'�Z�l}�.�S}eHoVm������8�I��6v8��s�9,�k��b�L�&/.���-�"�eb � ����E��Z9N��/K'��!M��#�.�f�Я�^���&/a�P2	
{�r�mE��+�J�$n�_�C]뛺���4�G��@���~{A�6 &��.�Ro�]0�:i��U�	v#��'���|��N���)�F�R��u=�S���0�@���1�9���C?'�`�CRy����qg�O���deŭ������e �]J��X1��D�{
�=�:�zn]VZO�ŤL�S,;�������A��ն�I�y7�`��:��N2.�w����(�V�m�Mw
�]h^n/���lE�K�p�������l��%X�)�-C�����~���rP�n����ΰ���7 ں��4Xv�c��.�� ^��:!������ᷠ��\1tq��m�Ӥ� z](�}fvb^��\\\�؆D<P��|.Y��y�$m�.N�zY�Ҁ^Ν����?�P��k��LKMo��pAI*j�� �2�wD>���e��'Ը�9��ݍf$A�e�%e�T�×�\�����"�z�R��n��'i�:��UK���
W]��l
ұؙ����l;}�9�u��٧����K�]�(�w��������1���m�R?/
�r˴D�+y9Y�B��6�η��JFY��H�m�Š*�U��4��&B��D���.�����. �wP���K��s)�B���� y��L[�����O��=3�㸷�orƴ@ 4b�sS
e���r�P]*r�[Bo�m�=Z����pZF�z{�R�"z��N�I�T���v�3Vnt�U�����NRs�KX��ܛ��?���Y�m�#�Uz@���PM��:�K��N`�o��f'�ҷ�=3L�)]`A���=��G��"���a*�^�=<�l����t?Tm�zL�8�0`a��h�m4�닖�
�M{K��a�����z�M�ۂ�����_j��Tzˑ�i�>��\_���ŢְWC�����I׹����r���:0�k�,�2�AoI�~����dU��\^c��I��]{��bƣk�0G��0|�S�;JLQ"0�$��
�)��D���^���� F7�r.��X�z�[��1��D��\>�lS����O ���=U::�n7�R0�O��1[�T�̷Ra+�����TL��i�F��Vz%�F�Zκ�d�9{�6�ߡ�<i� �.ۥd�I��̵[9�xj��>���ҲNL�u�7}ȅw��vءW�9�A	�!���}�n�/9{��r^��]J��ɀ/�2=�)s ��2|�!k�ګ��&x����"�J��=��77�=��N�Ѐ��d�� yNnK]�ޫ��"�
SI�a"*|*,6�2��,�ʓ3��"Z!�v�/�nx�a
��Ĳ�ƶRN�R��~�n��E�p�-�0þ'�E����� ���(O#>/v�b� ��.Ke�^@՟���L��`�F�aΗ_�8�z�� y�҅}E�DT�ާ�WU>�f�v��Σ��6yC]�PZw,���; ���"9/��"�-|���r0= D���O���v�HϏ��jM=tͭhez>Ww�-���F�d����T`��q�"Mtp�%�qu����%������hs��rlcve�L�e�r��H7��~�|g:ҿ惤a���]�i�2��m��OW�+���3�
Ԏ�W�g� #�;j�%����k	����.RT�4��?��Y�]�0@/`=�1P�+�x�B%�< �pb�t��y�Y�]�a|����#�S�g�c����	�:���/0c�~���67�Cxg�Pf�E|�ı7�k9E�m��f*�RۙI�"�s�� ����]3m�25H0���Y��"���l��+#�k������Q�e��m�tM���"�*��7���o���h�1u����}��ʰ�b� �R3b[G����"F�2�pd|�D\���4k�*�z�3�:�A�#M����>%�;�x�X�����a���N�O��~�!�������B�Y�*���{l�+�I5��@����œ ���h��Ά�����=��Y�����~x0��2�)<��]u~�����Fy1��ɰʅ�+���:L��턧��`�<4�֮۠[�L#e3q�J8GQ����Va�V�Uk=s=~���X��"Y��K��%P�
�Շ�hV�>�V7��8�[_� �����m1F^���ţ�;���֌|����|]�:��В��n��/��F����'�q�7�#D>���A�{��aX7��D/Oc����^�� ��Ǐ2�h���6�nP�3V�ޛn������&]�'J���u��?��C�E�?��Z�Y��<y8֖w4���H>8A��1�H�b��kk&���%|�S�J/�/��6��&�B�H2�3���0Dk�*����t+���5��pl*�p�Qۈo���h����s����|�%��a��6X���vϜ%V�7Iy'� 1�F�VI}�dZW�E��A��D2��і��8}�q�=%��hl�n=ɢ?����#���JÔٙ�����YpDa�5�eK���X:|���|IY"q�����9�)��`ѓ��,�麨�t`�S�U�QrIO�#wU�ҟ�]T��f_�ܔ��ׄῚ�J^�����n���t�H�Q�&�0?9������֕�|�,@G�\#B[�l��r0��S����x������$����ح���n�KN�P�!�S`9_(���ЪaO<���x��}��@���*�*ݰ���j��	��
�ӫ�4��-��۪���#0�騜�� .a2Kt�`+�ģl�"�D5���Qgp8�e*[��i����N�~���*+!�m,�Kv���ȵ�����4g���� .׆�D倆;)q�W�yz<�"�v� bmz�K`)˝=@�RN����x��ZO�CK���)1
d7�f�eȾ���-�fעbO����Do\/�8�M���)��R�CO���0 Eؒ�Z#�f-�0��Oҧ)��CxJC��ަ�Wz?ٛI��e���(�EyY����R�����5נػ�U^�Z|�S��l��_�q��b5a�*n}�ᮢ�b'�L,]چ�.��tݾ`(���;���ӭ�	O�w����E[�f��-掉��z�8�Zc]7=��"��{���[P}�L����I[���u���� ��},�j; �c�;��r�?�����w<x�Q?����ɖ�8RŞ�|��Lyt��+'鐏l���8�Ax^�i��_K��^�jeQ��S�M�Vū�h�]*j��æ�4Q��;2���:�!uN�t��0���H�����+Cb�<]�O�#�!������b>�.GB�����5��u�Q��*���~~�w�^��q@��0�滚������=�4�+c�5��&d�w7��=Fd��B�,��)a��?DlL9���3gB���}�ƚ�1�R6/���"��d�g��rf��;�3@�΃��� ��n�`ꚃ��XT���^��Ch�{v�^F�B㊗|~c��#�uO3��ʅ���t� _�af,��15󪥷k�J�+`�%i\�-֦ϸ,=��k�MÄ��uY9���z��=Q��m�	j�T������)�/�W@(�~4�K�R9���ɬd�c����t�˒�R��nۃ}!&7��*Ͳ��&^�(�OC�f(�N�d�<�Z�����D�3��ש �a����T��/����l��=mef�������w���P�c�yE���kUԵ����w����(>̰���p;�`��������]��0����~���������H���W�ؿ���🇣d������[U�ck$bɾ�v����p��W�,.XcD��A��QYVG2d�bh}�yƱ��� ��CF�Qa)@�	~��|В(G�D-�,S�öv�F�!)�WE��8��Hwl��[0�]"��נY�v#&�иé/���а0��8x@��߂%��9L��
��>o⚗�r0/����!�db����5��KY��%����Vw�ҭ��o�w�یx �*��3��Ddګo��3���S�>�'�^�\s��fǸ%?C�ۼ�w�8d�k���ZZș���ۈ3���s����!��-��ŢT���$�����.c@=r!Hx���Ht��b��a��J�M�J�4_���f`G-.�K��ECS����ய��F�Z"�j�l��Q=C���<m2n	�3���+��f�%9����
�)���ܮ�H(g�P�i�]�_i����B�>A24�9~y+{��.���9��D�F�F
.*&��2[c���g|�99�p,A�J��Ռ�o�����`��^|FH�vŊ�.�We�Ayy�n���vZ2���
n�v	���Q��>y�_-j���܇��K���6?n`��s���մ�X��pF(1���^��K�e�<������(�j���Èٮ���ph�Vr\��w��U��jnnM�.a�Ä�ñ����%�����S�]�TR$��՛��1�P1:;$o�R�x�`�[��R���]���8%aȘ�2M�W���͝�X��C��V [�����'����5q�*�1�:�:*~0n!OYZ��a-di|mӤ���؝ho`8iu�<�<��%��_Cc���C����W%�v��������-
��m��2�
J�b;Bܻى@W6gx�1^N7��5�%�*&��%&���[��g�`�{�T�숵�k�� Cl�y>U2 ����H8�������(���C��2���O��u�ޓ%�u.酭�dײ�KX���Oˤ;��/����Z!}��J���;�`�F��[,�����o�	��1�/>� L��x|��1�h|�m�V�잚C�
���iQ�U��I$�#�$����#� �?��,������#����͕yN��&��k�@]�h�����u����08�BW�	NŪѯi��6K%���.C�E,]%P?�ā\)TB��)j�~��鲛k�/�c,��X�A��b���΄k@�m&�m�;;������ģF��_��l�<e/�;�}v�Q66�LDi���'�h��m��]�^s�1���g��E�ܼ�#�x�<N�P99!܂ Q�c � DZtF���*?� ^\�BǊ]W?l��֣���!�ݒ�)�z��VY��ҰX��mWDo��@��R��<?�=�<�����:+��C� ��4��{|��I�{�����1��`nQ�Ƹ����n�������ފfѺ���k[��9Q�F@�ҏ��,[j�,�Pl]��=�u�]���ݯ�E����Ө�A�_�yYP�.駥���VY�߳�)�p62`�PX�Re��3�1���x��(	u��^ؼlJaۄ���<s������Z�q�o�1cc�Iy�떚;�#������Q�����;~����v��ǼbU|���ˑ��3�j�D�W�}�Ji�H�~���~�=�sc�Z1�aGpgu���5�r��ɞT#��Lt���)7`���^�=�Y������&�+	l�-F��8>Eu�ӌ��9� �۵~�}�i�Zq�����X`�p�FN�8�2z�LcLȨ����`�)6l�7����W��_`�M�i��&��N	�4L!�&=��3�+uǄ�P�ڎ|��d!s�Aҵ<���VT���u3��UEv
5����YY���i��^����/����d��)~%��yW$��3�eIs��*�����A��m�Ӱ���,<c��;4���`���z�y�S�|�xp0|�n	��<�(��=�4y��:0˞���21g�V)�cvb���D�%��g_��'�I�#SI��~�nbԶ��=�V�p����H.�F�{�E��3z<�λ�O�a��2��e9u�t�Z�;nd��7⬇�6
�ڹ��o�;Td*t��!��Q��I�l�U�k�����W) �"ө��ȯ��ʫ}���L1B>;���!阦QoQS�B����{��j?�I�t[^]�yY�쁊��id�.h�����^ӫ�w���8�d�I](^@�+mI@3:�;���ae��-��̼��s�Ժg�;��B%2L��|1�&Y�}����X3i��U�y�Opr]@���:]1�~eW���~{���<=n���V���SL�#tf����=��KN���Ϟ�G} ���e�ș�#�O�?{��	4�����Y��.�|�39�F(�g?c����S*��UL;����3<�i&��0��C{P�����N�p�=��E�Z�Ϩ��_�j�dCR?q��SS�_�l �"�X�k�o�vT�i&z���� �͞�,�����C�d1F��s���n,����h/pnd^�Vb��J���Ɖp���oC�W����b�����
S�,O��#�������u]46��-����Mu?�P"�C)�8����x�]�?T?�Ož���������a�z�EU��YBd>vV;jI�_k��Whe���`��Ұ��`�(%�~�@,��G���|�������X�S�\�eLlj�x��e��r����['�0�ar'f�˱!�򜳛�g�
8�#@�_Z̆Κ�H(�\p�?��c%"M;��	���E)�ON��q��ۥhHo-hS���W�|�5��D짼��m�p~e������qtY�o��ɂ���w2��G#I _�O��Sh���rp4�k-gޱ_|��/��:J��ϻo�ꟂL�ga[��i�X��� ſ+���'K�R�"&Y�~7�_K>˲�^���1et�yv�(˾���Y���R;a��f�hY����z/����^<�-��a���Z���n|�~d 鋟$L-Jmi̕���O���9LΥ_D��*|ccނB}�{���Q��My��
��L���Yg�f� ��y�Xe��O�r�qm�u�|J�I(��r�N�u��m��]]����7����8b�K�Gr��%�|>;e ���8PB�	�� ᚘs�_����Y,[O�ȄJ�
��V����A�Dіu3���?BU#�w�;�i�v�B�3.���)�c'_g��d���\*�K�.� �ZȪrl���@|Z���z�Zf:�C��>���" �b69� .@�n��y? t��S�����&���E��@BC�?ȭ���}7M�dr<�#'�������@CP��Q�~*��x.��O����@�8��E����F	x�Y ���E"�;4AbvO�xD����됋Nb]��"0��t�~P�b���b`��Q����u(���oa�ޤ���LK�<�f����,�%���`�
��'�׬��_���C�?��~���G�ΟMzH<.B�N4��%�%O���$�TI����akI���\W�!º�r�����tr�T��{�G�$��}rg��
�����\F��}K`��O�nÂ����$S����R����z����l����;�W�>G���Њ �M��s��F�F��Lf�OGu��<0N^O0��E@ ��t&:��h��qm�{4K;�Qv���3�V����E�~����?��`�|϶��i���^�%`}�`كfx����;�ڕ*�͎�_���=���V��5B���w���
�#P��|��^�-��0���:^�_0��6�`�Q]��zc
�*�?vw�*ۯp}�+}Y��QU����#L���/@Lw!yA����E3u���S�{0��`f���zxp���$�n��]둼v�����àt�%~9���.����Ϭ�@�2��?��mHd��L~����K�'��L-��\��	M��#,/p�/O:]���'��?T���y��A��iXQu��Qa��Qb	����h~�t��"���`2m�2�-���<P�пz�Uc��� ��є���C�#���As����M���e\h!��c۟X?Oc�3P�{��Y؏ģ�R3Wth� ��ö_���B`0 � �7�Q������Y�9B��,㰥�(��$��v��1��o�"�󥗄h�;�L3?��1���$},��k'���cf�$X��TU6t�(%貚���G �������� c!<��g�p�
�&Rl�Tп�1�߂w_�Xk���;k��B͠�������Z/ð�)�n��d �2MFkR����-��T��.͸R[d�Y�k��"(:R�t��a�u���N�*���D����1��Ԍ<-	���ZA~����(	�K��8���>b��|�x�iӽ�g+�Y�v�%�}��:Xw�^!N��.)���jj��o�Azv#u�{�\,?#��.1����Ow?M��*U_�)ؽzN���5���]�89E��1X�:k��W��Vϰ�#Zu�����T���,ط�Լ�Ӻ/��K��\@ I��
������\���tv�K��8��(P������+����g���W�?�'�kz����6���	�k�ޓZH��D:h�Kӆ
��
�?����n�>{u�	蜮�XXU�O2]؟�M+"L�� Ue3a�'�$�t�Ԥ�n��a�%�t"�_�)����"}��w��(��ל3DXkq~ղIC����#Eji�;�!&Vr{r$ya�-�I�*�/��_��ݪ���ڪ�R
2D�,;LI�rǨS[�]%��(�m�]����A�@�3��&4���������z�ߡ����6p�:8��}v�,$(:�n��󒼓�\�E��������p�$���5����0���(B�XZ�n�~-�PVe1��/�.���?{���<�ѡJ��g���B�*�
�(o��x{� �'�����}����#�t0�k�8����2��_#aL��s%
��|�p��IX�tN:+�*�.��Q4��i�z.�A{��>)�J�%���rYX�5�����hF ��ȶ~uv� ��=<�o�:Y��w��q(Ǵ��t�F9m����(��^�È���n��x�P.�=�����`�&{�����g�D ���a{��:����O|Y��E�N0`��.8\�H�H�<�u�bٵ�},8��ǉ]~��01a�tLf���`�����h��~Vg���:2v`�<��b�nT�Y'K���3$T{���iSٳb�1~5 �v-���L��n
Aȹ�{�I6���\��-�g�BE�`��#�(لL�Y��k<��П��1��@7�#*���rj�[���GG �}�ˣ�k3[5>RZ��V 6!$��� ��4�V�R��D�������B�}-Ș��l`s���SI�%�4�7AL�0��-�	U��ZH��m����N��Iƿ�Xy��s��\�<���@�|߸Ïa��Ѓ��ue�	�08}�D}�<��*�dM�bA�cLm�{ڞ&����K>,��\^K8��@�!�<�T, U��`=��e�PN�(̮�xU���Ra���#B#$!_t�B�����c��h#�Z�{g�0å� ��9�1�N��}���j�>�	5�Y�.�F�h�A��v�g�y=Q�m�'�&�x"Cy�o�fǉx)��xK�W���=X����'�Q�w�?��Db�lb�n���;�V���[{��
���W]��MeX�L���c��7�oTd�t��l�5��3�#��;�Y�os�£{B��G��l;~Crm�=����u�ʞ 9���0�q�EO2�,���o'�R��⢭?u��ES�F;
D�}e��T¨����*��0!����/i�.%͵��%��a��Bza�uP�K��%o)sЩ��F�
���2�&��g;�G�p-.T��I|e�a-�:�:wlBLL��W�
��.���#sppj�t�CA5ǣ������P����V�J�>T�\�T�����m������vn�arI�L��u~�-ˮ��ક�pkb
��nٯ����h���A}��O4��og)Ҥh��������^�q���az]@6��ǫB�~�R�nv�R֕S�H��-���	�����I^Ye �H#:�Y�s��鹹�+�@�4;t3��D!S��g%��gOa��W�Ғ�����JJ<1-
L
���%+weH�f�V��-�p�	��N����F�����ٰ�~��ޫ���?�`\*G�F�.��h�M��ٸ���I#9ٝ�O0�t�og���J.�m�g�V<rQ��8*έw�'Sc���RyYI�=y�3&�>(�{}J)��ޏ��?4T�"�ޡ/����.������?g�X2Uh�se|+|�"ўem�V�>;c�Xr�D��3B��߲@�i��gw���:��jæ�����W�K�~��\ 
8f���~7����Ʊi�	>}Ο��(Z�4/���%{����9!�3�Mz����G��otr�uL&��F����H0rEH�NZ���mc����u �J�I��_�	f	5�2��c�~^���;�7�xIww
V��Y7~�Y<����z�	/������̘�/����ٱ�Z���5������@�5�Ő2��D���Q+Lzda�̢0�w#�`�h��8�R7:��G�����Ãr-|�m�ӵ/�|s��x�:��9�񞠻e�5���z�@n�c3��h���=+���/k�8��5�$��I
�'��ɲ�+���l��o�p�Jgr.��w���y�a��]M���^3YtoO�Ug=����-�D�ٞ��4��B#��������F�ή��q�\͔�+l�BQR�`C�C���&�H��k��EF�y)��(��̲YuOb|�*y�x��Ӓ���������XH�T�5�d�d�@��ݝ�`�wWϿ=�)�,��|��o(��\�Go�����E����f���ۚF�HY!�:R��\ �s�ȟ�Q
�d����/��?�t��]n��{.�Y8���`r3��#���_�5�B�<���]@od�u�#��u��ݥ����<?��ވk��*�vu�|�����a�iʤ��L�P�����BM�v	a!8��0%�ƦI�=�e��"+�	ў�Enk�N�p���eT;��7�8&�o@�h0zeH�G����*��ŖJ�3�
�Y��'����J Ӏ�<�h�/���3Zha�c�O\�)
��U�t���y�Ry`���y�5*��B���L��9������:9t�� n�� )��C:�����-�k���_���o��bZz�U�݆O��D!z���n�;�y6�����Ϯ��F,�D�f:��)�{,���h�R)F�+��5D���7ҧe[��6��99��ϝ)d���_ie�C�?����I�`)�ܑ�����w[�����/(�W����%n��������G[�����C�!�X�@ą�y�Ul��[0)�q7��X11>J�b2�:Q.;��~6-���z�KMN�ŗ����_�7�d�����P��w�	� ��&a���7�@B\:I�'���m|]�ɞ��w�rƖN�Q��^n�z�*h2_���3�↉�Л���t3"TF�
,۰3Κ,' ��<9�6�,N�(Ȳ�~���F`Zd�I��fO��X��� ����ͺ!���><�C^N��i{i2d� �o��R#�3��q��#�r�~�^�[�uQ}�[N��5��wo���"(��A�o�1�49w}~��y��i搿r��ݝ(��x�3�=�n�+��(.�!���"�OJ)WGq��J�*��mF�а�:Tp�����G���J6rp�Q�-g* �] ��t'�Č	l�Vb�[2.N�@�)�H�n(}�e�?8p������r�[���ѡM���^��R������V�u�/NP�m�\�`�t���<�\�j�Az�����U�Ga����ӊ5>6��ɘnL?
RH��u[	��
��%�A��p�\4}���&����[�`�n1M��£����PZ'��]F��+����(e}�G���$�}\��]@�a&Z/5��ϰ�?�>��5	��N�޶ş�B�
;�� `����w#�o��j��ʧ�O�ު�W������:HKg���$4�p"0�8�􈽀����_>_p����Z_�gY�;��A�4�*���sr��m�� �p��j�rj���>8pZs��}�k`ou��\lTRd�#�oJ��Os����0���O�T��˅B�n��A{�c�%�P�}�dl��ґ\(>�ο�~�v���-��Xpa\%�g'�,b�yc�g�Y4^@�hQe+n!�"�H�jl�Ѝ�&|���c�.L��!�����_�9�tz�9e�¸�)8�z���� �B�s넞���1=#)sT�s���ba3xC���&ly�RH�r�2�^�̯��C����8͔���tf�v����P~Ի�/�aW87���I��H��63�K��9i����m�\f�݌̌m�7o�P躈!;�:����o���oI��0^��詭���Z88�����H��׆�0�1�� ���?�i�JS�o;C#K�x��5g8������V�$sY>��!��Dm��&��3Qy]�jaD���-�y(rrJ8)�{&J%
8��	��67�tl��m5��?%���������_'�4m��� C�Հ��������Y3X�2d��K��@4�^����e��0�az6�M° ��@&���g��g��,��q�m��}�^�r4��#$�e;�(L�D�(�؍��M��ê[*0�Dge�-8s��x���v�L�֫,����vn�$�_9jEP\��j ��W�pnPtx��D��@�|0�IA�� %��t�v֬����?Ȗ�b�����W[�n�I'��衦��|c�:���!��J�$av"�6��4+��&����v�zu��T��$���=0�*$���\o��$��vugȨ��09%3�`uT��UVn/����OҢc����<} :luA�.�u}��Y����:�YJ��:3Ns;n���bR������RG9�Ya��q��-eE�'�.?F���"��1?���k�ml��*(�4�A�ZF:]=4́�Z����R����U�BO�>Z�S��S��CUx����Kbr6j�|v�I1C>��w�Izߠ���,d�ԇ��Y��R9�>L�`��R��1�:_�d����]B>m�3봗cG���W�K��S���t�R;�ފ8B}nBN �X�]��ٲ�J ��o\���^ި?���	������A�4�v��˴:t�#KD��<v�5����Ŀ�M��ΆT���%�i=����h*�l/z�S+�J�.��c>#d+�7�Ok{��Mۃ��_b@gZ]��w�H������(� �T����a���A�.��*$Kyr9;4]F"Ъ���i�=�j'R�Q��)��os埮��*C��fQ��8�-I��:�[@GD�C�\�"�;�_"ui͉u���|n��3���+"=�Iֽ�4Ι����^$l��;��^c�W��q�BOd3��^eU�l�>o�
�j)D�m$t6����
��_&Lm@��2Lb�<���[(t�D��iJ��BF���v��i�y_�&�M�����ʨ���ҏ���R��z!ѷi�O����g�sB��?B8nGQ�_|�J��ҫt蓼G����:9j���Rr���U10�G`ޮ����I���Pdʺ��-���)��c)ԥ�/���Xp��Ƴ$09��V�g��{�FyVȕ�T6�&����ksB�<��\qV�[��%_���/~�a���Jcu��f^㝒ӂ}?	�� �7E�1�zCj|��ŴUz�
��Ao�_�͋��g�[��l�J���|�b��{��Pg�/R�i��N��Ґ�(5o�tF��M�H�UW�|u��~m�y/�3ՙ�߱��o��륗a�䅗�m%Nk���2`X^5��sG���9�D\�[��hp��{��1ArX����K�9�����R��&�m�,o��R_>ǽ�l��}7�����������;� fy��>���(���06^��MA�p:>5[/�����'�̄m�-:	�8ѱ�i�8�^$Ʒ1��#R
��9O�/Þ$�X���A��?毧��Xv�<r��s����bE�w�V�=vcxNT�O3PfT�*)�f0�� a�ou���]�3⥹�R����{}P�%���W�fP4� fx�U\��V�.b��J���]2��Ъ���h�d�\�¦����#4I����i�4a �[z�����:1�(�D��Ul��>��%��x���;��Y�A��'�:�	B��fj��SX�I1���mC����}?,�9A���F|�a��Z�"$ �Χ�SK�f�/�1³< #���.
�h�{_�?�on�_8�x�آ�I[FNIm#�1%����iA8/���	�v����3!������5,�܏'6�+9��)DW 3_{bu!��>�#!��^I���w���DY���Ө�&U�v
8��9e�����x�9�����!4k�~S��g�}���
�����b2���V�����r���X��9�!A�4���4P���  5Yfܴ�x���ߞ�G������K n�q��ɋ0ʛN~��#����Q�g� �WJ�,=HL4�٦N�|�5�*�6�[�ƅܶ6 {����\�f��Q��C��h� ~~��5GtR�+��0�K��$�4��I��-�le?V�����]Җ�
5���p#�PmZ�X��FQ�l~�:�6�N�IH) VMn������aR�(�~9i�U��A=�׌�����ᨱv�|3���y�A����Ϧ�v��̮
�q_��"
Q� c:c��v�=p}�ZAB0�#��F0�.u2J��Tˡ3��)�����=7�fkpz���u��;���=S�L>��ۓF��-���n�h�jk�Y��"�@w�;vy���Q�����C�J��=�9�P���΋���Ŷ��Id�({s��u	o-�!� l����Y�}LQDƃ;b�#Ӫ����'��&3�ɡ�@�����?����]�UAR�����1%��x��`��"��ٶ��󙱊w�^��6F݄J��<�3�	}��l*����tbl�#���wh �e�k�A=��u����s�e��=��;0��Υ��'2R�|�V'��}�>�T�3�%�BUKV=��#QN8�8稗���l�A��#S��RV�7ܔ2�a@�Z�~�N�>���T�Xr'+���J���5��$�Pn�2F���U_x+�@���̙�����P��s�TV�]2{T�U�� �s=q��2���1���PǕ�v�i��i�b�n���{�~�>?!���N���JO��[�0��^�h�{�	�%Y�D1����c`
���9.�ŌY�3kr{��C�PA٤wB��J�<�����q�t5� �H	���w�z���~��wW��;Md����b�A��ą���8\i���u_���l�P�ĉ��)#�1^=3">���̧f�{�O:��T8�3-�H\
����4�X����12�xp[z�;�u��`���`�>@�Z���;8�LC�^�J�i�k:��%�\���p�x$�C�^
O5p�����c�D+���C�u\����	��P�G�)p,��|�2!�nSj���O2���� 	U��4Q�(���ۦ���qk�"���uA!�M� �8z繢��Oasm�-ɒ�\d��_{+��鈘&N6  i�����	SM͉����9�F��	6�����aq�G�+�wb@�	�c U H��4�����M*�ݥ���D������"�����h���PRy-d�<")�6�F���1՜����9o�m��3~˶�N-�)��݋(���0..p��(m̉���	aTZ[���D��~�k
