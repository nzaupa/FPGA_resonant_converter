// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 15:05:48 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CUH1xs9MYBSpu1WODehU7XBs8xA7MgR6b9fUA2R6UxdiMWWatQ4UOHCJVaWNVydX
jqClsSdMq+fe2g6ERWsbIjLI9b9M0byYWbpGxwv/pXZCK9rAXOmJ4j+q+za1/Skv
1A03E3bO5Jiw3okS38N5kuisMDghz/ooDJIaryjEzvk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
7A8uM1Pn3oBUT1umMxXNYhSQMxLr+cUXr8VPm8nmdfQTe2KGGHvXtAr5+zJp0xfe
x+r9YTkZfo0p912Wz21B6Zi/B/VcsEpA8GtWebdk5SeO/vZbc0Cul78ky78ZHniW
Q++782K2twnBw4rhCwaUjazeZDj1p5FuXwh6wDWbEXUSpxkXUbZdzGLECEGOuBma
uYE0fM+VzLtfCd7UhfYDfzNXHCeSNot5rPY9hePDz6hJwGlg58UUle+92dvdyMw1
I5WSOrGlRLKj84kNj/x4zfmoV94HN5SJlL7qL2yk1Zvv2MP7t/8YRApeqze8a7l8
p+c1GSx+DtbVYaggZa6aM16lugXmD76IeCg8i0c6idJG2kHocU+2M38hrcDJy0Lv
Yh0RoyVQAQore/ap2Bm4Nd8h9REODpnmezVtPtM2FiOgtRkBrsvnH4b312T5Rn5m
nfzNeDXCI8s/AcenhPx6KMTaJavlQQ7a7uTy1/Hcuk65iFyINhVtrKkIC49uP/qL
UcmRhVKN/pA+DQprRXFcYOme6km7v817EhJrs97xXfph5hGxFnyGCnGJqY8aKYQw
EfHxO+AwmD1vR+QCU58dKotfDm+64FHohnksV/aNo+htdSqLtnJLP62p88EejJ8g
q5DUNiNPYirsmrRmQKnqN8b+ZpF9hShSDNyKWfQKj1ig/arVHTmCXTLCTy2k/dUl
VNHxdnSYZv1cdxUkO4tzKIZc2IjVb5ivpTrpGjcGhEWvgnbx3yt9RqphRNpcbIpP
7/U1Tl2/928p72+amCIrvXCZQIEEZN8ZAcWuqv4EvMI7Oyz9u8RROkGAOtkfUjZ7
J94Xn8e3uoF37hSP6qzPFTkW0nwtHEF6QTUL3N3zIrtQBmzZYSehwunnOmop2A2W
WuEAzIpHpb2eAfRclMkvdVHkgEmg0vh7SJJXIw3S8+Dk2FFKrj9mgCVLXItSfqfi
JY8EKfyytJViE6vYtaGgLEGZywh9G05wiVM73szrmIgp2JnhgxNmLdU1Q2xT3Czw
idmNiGr7UWiNTXmZawaC93bb6xz+d211cNQbvQ5QjiiT+ECR9MTncJ+3QXlZuH6/
kWchAOYsULZhRtO3FOvNXjKoaO9a/J7Gaev/YpJ2GE34nUO0OHe4F4v3yI92z095
H2FXN80NxtaPXthHOx7w5/RqUm+im2+4kc578h2e0M9uPrJRFPhbJBm9wN/OCYXt
7cCfnI4PA3aXuR7fh2DhWkN3Y7H2zmf0c24HxwCXCtZ0yE2Z7tgVB74sL/iBZHuo
DXbQEuRp7iqVWTtWwaA8UZfCFUlB2BTyz6bRUQOkn0xFEcDgpvEQAah5fZXIH/q5
b8eSgTttqo4gBlISy41al+mQkRxWJPmvO62R5LulVKX2uRp0gEafPa/2j5ttbcMX
ipoBlafcAEaTsVwL3izVWQ1m3eOpaA4I6rfOxZmimgimdCnWq2loVdNJAIB7G8Jy
t0UR+Kbh6ngaLautyBfBwNXlhESszgIe3WH6SUG6dlFtazRFNXjYeiH8+JFoyaJ0
e5FgDxOwZ5RUE76FdkAwhjbdkFwCwicoxqa5XftqP4ymqcFn++Pk9rNi39r7P2FC
gpvRONzBTa0enejBD4acQcSqUyOqIBG36keMY/iNt3qL+ROGfE8wj9i2UKSsKqLi
tVW+lHQws6Xu8vFIm4j4CSriclf3w9mjX5OiBnOQdhEo62Oxng8CzMs3OvPCN2Ql
Dp06odoRjDlJxrQVzM0gBv2gW4a8buA8Aqc6in4/nJaIp/neAzvWmHhv5H9ZZ2wO
MDndhn4K4a5nXFV5+Ft7F1KClg60h8iybyaLcMV0nkgBkXXh9AlU5vhnsU23v9LW
V/WKo8Be+VuRnkyqzZbpCfoorj15NIT7SN6TDifZyBoLpVKExcQ/SzNsthmye1z4
fdbDPsobLdlQf8SPZih0/TtpCbgijZVQGBy6M81Xilu8cgZXjuJP/GvlSMgwXfLI
FOlY73Rw9TByMnqYa6a+e3Y1O9E1b+wM9J8i1pN3COml7hqXlPFYfGk2OK+636qK
2Jzz/9aOOkLoIhtV/i7YekkDmr1f94wxewyb/r9lAau10OJYd6Qd3Z2p5lET0fEV
e7mro/TLYCGq3eVz8suWUJpJG0H2YONBL5vcGxGLEPt35zr4B4b8DHFVgUqKlHEp
Teg+nxTVPJYoOTv4n8EaoFljnqz1TD2RISonGlUv/JRo6ytJVpXvQ8IBikFSOtHO
dOlZwtGZzBF7rpWKmjbXsOn8BPJEHRIxbQsrCJWb1Qf04GSCOo4EpnvHkrzgKKZ7
fkokJ6yQ3XrX5x6rQKSWetKh5bSQEJUWcAHfLBMutthcqy0XZDizpo2NC5JzyGUr
gr2ixCl2cJNV4j59HCAzvwkp8g1sBdc0+hSFnGTeBE15qSWU/rrygNgYyagaROC6
h6tnHGgL11OTCrL4/hdj1kads40rubz1xFCLUTGd/mRXC2q2yqngbksMVSRk86O3
KR/6Ws0HpU6xbjdxgrhXv2MKBX/mH+6XQ65FnNYl3dMQf1jq9U/P+SpXm9DDzYUx
v95TyWH9jcZFVdqb6K/srlJAjFghSH8XcIbBChDVNiu1l/JVF4JX7a6ZNxOW9fwb
UVnjC5PexcvLojE5AVV5tcYCBIkleoIDGNvM/Cjqjd4pFHKDn9LY18mqMNShtNFV
k9fb0k8XqHy/kxNPncW4rmfjDZkJyH3f4H7YqgH4pXWSDb7I8PNb0s4Jk2kSOPzN
DxlVTYV790fpJ1iaq9XY/C36b8M2EhdP/Gy6e3i/gPP1l1K+Cp+EwVG8RpQrod5U
fIBjf5pPB96zQnZ/Y6YB4ShZa4p3yxVMRhdmyTdPHuF3qLLaQR8JyvvuTmSqRNt3
MPVqFerb61+afs7i07a0+JxIhgr7eyKtjMNzQrkgV+WDM23xRnDYsF9z/HRmUYmB
XiTE9b+doUQ++tYHnIg2ZaBjRbWXOpBDZqtIxXkdQKTI+GP26YSPqOqCZVHqNcUw
UYjzfgtqF05eExxKuvY0IjMRylmNzIDJrw3Bcrrf+dUBYJ7UC2oMhXNayOH5T+fP
ICvgy0M/WXxqY1V2lwIqHYvLqkGEC15rldZTqve/E7qnDy5SXxFl/lTlIQTxjSza
vXWeoWxNJVdaeyh8Rd/+F9XhNMSBjtp7Slp2J4jlbLwGSGXE0Oh5c+wJlksB5s0s
7nDJsybMFkF0hpbMnvTRbmKHBGri7V5PPg9PCE3tlLHb8aBV7tcTdMsLrFouOWPr
+KXFbnWMkeSSFBphmPnxZAww8idA8quYnXoLjWK0EytZfA8+V0l3wL/Ull6qbmq6
dIHsaMdfxTzhl3P545+7H7UQSUTDJNAf55gIVQUavvZnV4X8l14G4gNi4XMZtIcF
rmP57r73yPayypTnZcoJYdtwxILEJBfqxXL8p4J4nBMH4hRDdNYzgvavJdMB9C8R
eUcuxw3cqBmlLR9eX+aHNKvDA28xSQRNf88T0jh6IBYOBY5wh065XkIpAiuySbJd
3EV3htvO3rC7Q1ziUzo/b69klwHVYFAoTwTxdDIRzilbiCoh8Lx/1P+AAiAGetKg
3gCaSSkz7LUNG99z5V54RC4gnV3P4Yprb/syEiFKalQqitRjdDkKqPynxCnZiCFA
MIIBM7SKcg1PNNNjF6qRZEYPPe/ivnmcvJqK8q8ng37IVKeZz65bAbF2h67hqi0Y
yNUedFMCEPV7cZrcK5z0IZlA8w1VxyPV5eJ29b3P5UvYErbw0hnPV+2pB5kYRRUb
FY6NNZ5c9RZL5mQKU9vEDK7dWTnXfrmHNmOplNz9jbpWvo6v9zImRxVPqOpxAhXT
hoY8tulR7jXdeukzqZsxczTTXzNMQ+KfQ+D6U+9hutQ2C+gW2Uoevc8yqg5RNi9n
664ieB6DdtzKoITDkGj9bi62vMEJN6m+vUvPXJ+wGWZqNzmc9XJnLjvEc8KwqOE1
VOvlqscMZaELp8RHZX9SRp7utoqm5hHj+8+QPar2jKjS8i4POv/zm8hXV24zoXzj
W17lkIlxQ3DaIO+XyoCc+m8iXTzpTE+PA4KkAw4pg4HHU2dsKQOhef8EuvhuiA/q
QXH5MXM/u3dLoyqSwNvkW1zdDTTiOt9N+MBggu9+AnU=
`pragma protect end_protected
