-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TOynWnpCGHwSLrOkIU8g/tBDB0aQWekrpmCntPBtTY9UubUz3S2wcV9XrUcoa/eFuxAAPJp5DAQM
WYwl2qFXw9G5AtrtTdNuCf6q8XT9kNY/fl2SW1POq31PCHIkyL/TYFke6oGwgbxbn3e0Ei6eXASy
3cijXucLm4Ae4IHoTVUjXi7uTRB8IxiKfm3o3I5MBv9LnZXZ4pfQF+n2bkBFoT1ztObPxS1lGpSX
wE+DN41ByOCMUQjEU+LCJkSviOtFgWUgfOtAlRsJzAAPeni9cZS1MD1vrLUvf3IlDwA/iG5SIzda
9Wwc/JU526ZUIkMETBRP2dpnnCkjKx2xIqvnjA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8048)
`protect data_block
BhgvlPnSQ3JA3jCDOpVj8qIR7DNwYztQlFEwKA4+OrvE1PDpJqFQNn1BfNd4rN9Lm+jISvACpncw
JY2qf8fu4Ox4h3dE1pWhtT5NxPyZ90AbMtxItnJRIqBARdvkWCs1f5e4xY9Uhhq145asLOPAdv2O
SUzKUj+ULXwyeXQynvpMp6iIbeqfsyutAxGNZmHwYmte+V8sP59WFjZ2gXKkjgmdVuu3V/u5E/74
z0ledX2gG7C0l98Ywbj3bTr6Wvg2yKk6XDDEj8F9qd14x+bct6n73F8iKoOkHYwNX3ee4Fr78CbW
S4AXRvAH4rQ7KoUN4JG63Ri54CBD/KRxoTzvIrJODaZAZkpEIzPBFtZigqLwJlfOE7j2a+MOOowm
zVZB70emIy/hjQC0d9hMFC4NO3qtqbOdbBtY+LvZVFw/a1hdW7nmY7YdMj/QbXJlcTgXfjBhb3Yc
3EkOEgTKAl+pNGJd2RPn6P35bv5yUrcn9tnlRPPxc4nnrSJxAbjHsl/QmburMCGg2Vv4wYkYVX+i
ap3UnHt/x3ILNn00ZoBpe1Y5NnjnpmltaEmH/VYex7cAEsFXDrm9aazPwlu35lVLxVzDIwDfrQFC
TuR8ZLTJMIonEiSibF34tak1y6+F5Slaj4eNggRlv0pXUO6cN/y17Q+60sAFRM3jFzX3/7jS4lF7
UjgwSZTFuhaRY7UDf6tJom6h3vDSlhpqj3VVd/eIQCvSBMIN+86KezKa2Jq3FErJDlzSaDAdcMLS
tOEtMD+itfrBla2wZ2uiGMnuZsa5wuQmW4R61WeWrVrkivcrJkdtiOuQVTUEbyx4u+eTyegGOP8P
YSQQmkNvaamiIOnWEc8GKKSsUIRYukWgZUQD1C3syeHfNRDBDzAQOx3OcmIw7kqxZ6DN+A+O3cX7
YLH3fV3Q7OCr2RQ8S2Pb8qXlCXHWHvQQz3EV+UBP4ePrlqA3Xdyq31Bon53Rw7RmPxg+ZPb8ZiyH
dcS+rqIKC4XKZY0kc7Y5Phq3JNlb6VZKKT6cCfjyaGtBEu99TAwnoEzThyrFeQ1CROZhcKmRbKyb
Q6PlWcQKGA2L8WmyD9SiaSGio30FyvVFnbpPG/wRGlrLdGHOaoOwRu1l+2pqfa+DvZxY51haV04s
8w9nGAoBbGcmWyFRDIqzSt1vPMOkv1RscjSe0mVO8+DJvD+b9kMweBWDZ1B7dJAJvekRtQRNxVhN
RLVZAHfhAXGMsPL12f3q9Xef0+dGpRikm2qctko1POB/R4H8ckI5/vlOGQat/d0Hww2XTgi0r4iQ
vB7HxQ4xtqs8pjiYxVUvcgyCUJD7rwFJwJprydDF+EENb4BdWaFZS+0ojHvvqhpVcWAtk8ZilQto
orXFEWIqLrzGLolTG+S4ULq0pAqGg8owm0/y9ql2sv0wLaXePpKBh+/5NseHk/1pJQszCjbKlFxX
CM2yQFSd1gDDHxQnznsTwSn7PzmaKJ0NEd59Gv4gXK6pSC/M3V8vyoQqwlZhdru77Zef6dofQTFF
pxtCpdiY3SfF7NHMkG9Y3mUtsGFIQzm9+1jaM1nqt2sxh1O4/+BmYjcPqY1v24IqefpJbrkCaEZe
XjTWzUuLSWNhwEp8KR+pzH0YoQsvzzYajkSYrG+11fXDHwBrlCIyrE/gQNvBtnh1xHvgBbZftLaf
uSs11cAI5aAhchlR0MpBr0Ud2sqAtPS/XGrml2Z/s5v9XmduKTg65M4YIVhoePYqOvQsBlMj5bW/
Qf+xwdeHwD/+H7D3vKxkqdxJF2eSgafa0Kt9ZDD0ROeWOExTn+2z8FOb1llwUAdJLsSUQFQ8DK41
eeN+jaqHce9ssEvuxVbp1cdcppImH0flE03ZAGI9VCY9Gpd5A3i/NzdpEgXBgDRF+De2ZhSmQK6n
CsNFTdkH+wejmrwyXnVlF6V1le6Y3ySajJiYOsr5+8dYy10LH1+8tV/Ns8Zlqhp/KNilQScfyW56
UDTBEYEGTRKUiCD/4DSZbvoP8FoSC63No+BZgDp+vM5XRc1InSf7LoJFy+i/QynexMmbyMJrhP1E
2ro2+MM0rU81YZrCns6ROsNj3f9NWtyHkNgaSO5EaXBA4nMZnN/aGiGcwGGQ2dKGnDR4Q/dxV5ij
5HI/PSdz/Ja24V6zOE42rK8jaHT4VNC0OCC3sQ0KWX3pIgcVN3SyR8bOOo/X4LWAWTRmiYQzm4Xg
Vo4/xo4KqTHI9bpl1lqo0WeVvTiaOizy4voI1JzKreGChvpixkB9zPi6s3XHSl3oQNKMJqWUubGU
YpbwwSEGsPt2vJQ6WZJJ6tGDlr58Yzl9PCF4vTWTyM9NMCjUs79ZR9OUxl/b9cR6GS4hF9wiF1s4
vSMNOINBA/fYqRk/Te3eZCvSv7qjWnqoPKhx7Tx2oxhhZXJG77Y9p4UKoiZiCfnPKtqI2KG3cboP
nZKthBGW+Krj7pk/NDP9qKDrZZZpQtz+Dm51wqErocUp6VpvtEhcdzNooJalDC7Rl1SMz33XP3oY
Oz9KtWdkGgXcNWETHtn076NJ3QGAm+Ul4e1CyHkBae/Mp7an9rCzjuiPByUIFG0pdQN/rfCaCbXy
/lj9TwNO+islXI2HbQoL47sszu7DT9r8JLdsrj3ULWByfSqSubvrGB02gbmlyyx8M2/czzJYljUl
eB94d9Ve3JUAhDPgJDuB6vkR/dk7yCzxgkoR5pcnySURSx3cfYHbpjCG0msNPfIyNPiCv3UNhea+
8+TP9agCjSNFdxoPT+hW1muqLtCM2jY3T9TAHnOdiLqPXc/LMNE+6l8DbrYn/VdImW6dWLAPLCAJ
hAsfeNf6cnMNIR0yg3rUAQi+oZHQMTlxhjb61CNfj0tl/mwRq6eafW7YmBcDA5H0WLcK5CfIk3Mw
6YfO3fUV14nbFeLux/bpO650aPZlF1a4wOoUgF8jMkurJixl/nP71GvVxsElU/6Tmq37QtsUFnq/
HQGeDDfTw6A1ClAPaWgaysopH1+MkdwdnzjO2gbDdAdw19kttiH6fVl/Z1lWRWW8KXSnbq+i9FrM
HKMaWSQj0Ju6Q+rlyYGdexYqXOA0ebiZ+VCgfIG6BSCNTmpw7D9Fzcvj9Wfxvix3f9AQ6wjd6IMp
FEtDsjyTszUj6J6rblZG70L4ULKJIQiF7lBklXgZuVOKW0i2WDR3/AdhtzJmS7GKxCfCsZ6Xs8Dh
ecwob9ludYXoMpIPzl6KkRy+ze2SwpHix8eOtuvcW2cMI350WoSPj61bt23V5/wtwYqYo/HCIV8Y
Xq/3X1duyJAbiYrsR7q8sgnuIsSidOLj7lORXipIguSw1CH98W4FX4cYSwL3n3ZxFPMoSM5bVaSI
FyX2UcwUiIDxVwodHNA4FHzUvMqGP3Tg5CmIuAlkZGvV1kyjGsC1PTtpgX+2TsT45qZBmvF5DTF/
Iy1yCge5oVckvFQ2sC3oNqgx9rmw3F/EhgK1PFzkVs2+/c2wHjvCRN/Opox25bz/zD+Mqi9CifOR
24YwFsRfjBtLBTaXBWHZWVDpWlyoorvFkxCaLrJFiL/hgsXgZbL6BCYnHnQW8hUPSguUMd9KWe1s
qCnailDrA8FlzT++Yt6m12SvBgqgoNclfhjHD7M5N/1j/3fbGaeqvdjx2g8e9ubLqqYwQ9vEHcFa
Bs/CSb0xJA7NsJVVsmcWqu7z9GgsUXkzhq28nB8ma8136iNvySwWZsnEuVmy+eLZ1Satniulc2eZ
G3i92nodrR3CyoJoVxrDZ5ebMBZEgXoLsLw13OxY624p1qXlE+/iX++PvvgKjrofP3gI4mtkEGF/
OknCg51mvVrk/nMo+ShCNCbWZWT+KaatfGR594p4UIGZJB/slTOA765lgKXy6gvlZhoK4R37l+MZ
jDpwFrOb/1lvF/2EgigunbjGqhsim27DIZEDip/jq79846SDIqre997GZKc0IyV64PjbC3WQ4C8R
FRCbZoDG1IL9K8dhljJsHxBkWTMKsLIODAIB58ReTohygpimPc4lDYSIhfLnCdzoAm9OJlBtl3lz
VszsObKKI7yBS2au7c9iDu+RNeqSqgPTD7lbWxO21utZiUjlDYG/YSmG4wMU1xkUqVffZvU2xMB5
HApagmcxqSX3J1Pqm6Km8HMzRyruUyvN0vC4d0Opo5x3V5kIuddYybKg46gtO8aUu1LhH4OoNlyZ
8H3bDr1uYc7TlM6h1e2/cJWQqwXpjeTRLBOzHk5uDKJnpGtJa2R6WVyBD93mNkt3emJcE2qsgaog
xHj3duOSyvpgjvBPJv6MzVtq8QFxnRiADkP1mAnxckMmmTF5ZYaVpDu+Tvk3IdcjXSrU6RDEmVmE
9hQ/7qWtuGsK4RtWwlA080Wpu1taU+Smj10NLZjHLUT8+tfTuA6cmtm7bKZRXR5sQW1QxotPQYiP
d3FQ52lQviXizbrs59R55xXnoizUNd7JUXWGqMkkyCtbHafmkZHPRKi0S63Kmw4ikoqFwYhc96Kz
kAG+qNqfpJasWdPbNx5xSHoYJGWZvmCQWmPeGON8RwlpS8nkA/ap0Y4Ouhco25jlSAr/xOGLJNjY
bEgrWcwWmTAkkWYJ2fJfV5lItJPgj/Vt6mcY5rN1yzlD4VTvhG9iCez/d6fj3EmEYD1VQT+7Oswd
cjnMt4nUut/iJsG7A+vLbaZTWrwYMCCXe8SuJwpO4jxbPoH3KfrHvz8mbF41Inpuz8pCJd6z8yXf
w0TxrA3cZBBElPzGlXelUTV14CPNTU8vQNqzP2plT7uFVoyyxdP/ePTENJgwAXqgNYI2+/IKRtv2
bhhWlFCjwEiImwVbvV3wuIXTRgSCblmXk8uZtw8nMc9D5BiOBSVGeGRAk0+qrxfvzSqQXazlShmr
tXjLMoA4P/f6J2VpK+tPvLl3pSqh6TFBwDn04BipGxtUIfkV/X8fIuAFXdhV6pkT45TfcbvxeIpB
95jjPYsU7/IV67t+PYYcjHfRfB1W45IHrMo2jHAbLMD10wThymeWDA8cZFDajr2s3uw4TUTomQVK
hkUsLFYehenLSJk/5gi7C8YBcTYILTtcdG49VU2N+r0Rtz7XhOHiJEv/joTZ09DQE8bPySHxOoH7
n6MuGfE6+2ReXH8x61jIYJM93v6eOrnyPHrAhO1YY9/TB0PZONkQBjTAd2F9fMY+8t8mZy6KFj5E
AySBg1nYENS4bUKkFR2Wak0fNLdXcTlnjgHfx6o/TSaFD14Iube1o1t9m4ydtTBRrjvt2/IJ23/h
PEEp9eivEMc+Muggs4OyhbsrS7Xs5+DWDTxXwfmfBEWrjsLBSGu4bmjzoRH/TKLbkydZjntyDyCK
C4Q1V7S0AshZq+0SQBpLEK3jIrY3oQUGT2P2H5SodJPuyBlTEETSmG4gVsTOECsk7d4Cmd8vlLJj
1xqxNdEqTUBJP/2ityzgCPbpq5lbLLxQDRJIOXy1qYSmooFgzyt0WCnyMjuJROuUVeta73Iwifh9
5Ac6DNBgscJ63HcKLTsmY7ZzsINF1zmqBLt0SvH8Dk/ajU9uWqrJpVrQrZxwFuqRuONDH6QSmNNa
cQZ8TQbbX/scYSRwf+TZSrof/pOVG9ITtXDKxY7KZjjClp7fUNhvyq8yD9XIDnMra6TNa+vaKE4I
Pswb8SejgNQ7BjW1jRORNHQSls0cpDRZ/o/6WaS47lni1fzWOpRrekhTNhNdNqJde6BEWEmrnEtE
zorMoEMqjOykVru1CCIDnpVa5H/fsLfgYYasblT1ex3yn0bdHkP0a7qVHhEQFhL+mU9KeaFKqFBp
aTR1jGDcMD0qE/7/kimr16EkLEsy/wmL/jU5Z1gusR/2yef4C/CyN6U3TWn536evXLlDY+ONm3bx
Dya+F2rowg8z892s0Cp1m1gF3f3zTwAoy4bVXAATyc/Y96TM1OYWwMGzAYAzftRUJK+pd0KOMpSK
pJWTvtXaWHtIGj8pJt5UWMZzvxuVUWHaV4EODnV8cpq9PIwh4GtiUSzY1nmwv5zGa//5u5Q52L0B
5N0nLEMqg/dleS/dS5whKmn783NCc3++1hcmnfRjz0/du9QWz2fAnwcp1xQbFHsIcT0VRhAtMSjC
AxnYotbcs+GJChXP8TPUFBmJGx+b6BzAihWbQyfeTLMJQpXTJyP+oNK6aeENDPPi3avptRorhRpB
Pqwo7CEMOi4+r15CPYp8yywch8+jQLNncRfYV6Q2DUQwhc/QsgLg9rkWSgEASZWsgRlTA+GP4FzU
rKcW/KYnYH+/Z1+wC/2OzRp7Jdzgu7GjngjBpzT31rZMXnCV3dpVISyNHzIw5epd5hFPuDXmzMkO
vNKsuzByU1Qchqw8dQKhMPf9wOHdgx14libshB7qnCNFeImDZRPq+IZyffWfptNL9FeMpnlFMnrE
rjyT1bTzVPRqthJubuBt8Q54DhB1RjEqUzJ+kvt3xEXyKBCcaaw0RIX+duabcb2PDVyzecOK6DyC
Ose/Hf87klN5cVUq0VhkFZnUd39BIa5O7b+oBpfvs9FtLM1lNdtWSjT526EAggPSjk7v1DhqYhjh
fkS24qtY24KoTClqftAM99Ni8EWlGnNHg/kXcZupqzZG6NS/ctbDHcILEedVzatci/Ro3yPP81+j
ILEk4DT537hmoE3SeDb1FUqsOEA12DtATSpXMfKunZqwrFasHaQ8puwHQgVEFEepkRkyf0XyhBPo
xEoaQy12YlVXWk1ehPJvqdZWTnoSnfbLYARpsE1rsmYLWBUs1k42AZ8gBM4lN6GJ6nT98Dzpmn60
RqGY2xLZRW2IEpS0MwHmyDK1bX+nYLYrQlKIRsCNEyUSEBWDQ68pry8x2a5FutYz9/o/NGjjGxXG
MNlvhuZB48WyInNH/4vr5NLdWtj7v5OT01U740XyVgc/OHWcSPR5LWQAsvbCQ2JdTboAzuWkBQ+E
9M/NLRJvSkeM8GpE9fhN95pU9gdkmJTMFziwnqj1ODhTWsvK0TZEiImzaiRspdklM1xFqDo0Ksnw
/8q/mwDu0eU2ZHRy/40sOA+sZpoZ9rDb6fEIo7bsgR1tgwI++2MQdrxlDbPRINouFH6HHhpuaR7L
tvYhW++A4octgQAcSjAsADGvZ1RwTqfUYr/f6DXCvuvdMCJ5ST3O4cHpteLoe9jp5CbGYeCWbL0W
fwRfHnT9G+AcKmipRwq3d86SaoCWPYi0ONogFnr3Eiq/jbqYXW76XWT48KVelkkz73anHIZAsJdK
HJnnifWGsasglg3g44Fah67aa8x9kz5ob6dhNy/b5dHZI05a+8T84EB2W/IEBuQ0pWzZIP5Els6p
8hkEapKB8TeBGbCNBlPwxyjSzY7WemZ4DfB7OuK0qCi8PhesFkVuDu6xnoMq96Ts/uGMg2OvqEEB
058SrVZX7WOvv64opgM/ePgLseGXiSK4eMMdmFPK5D1Gm54LCMlEZzARGfl5SRP2ScayhKIxYk+t
eWTi4qEKFybAhyFH6T212mcg73H5VzbXb9RX1TLTW0uUdGaYF21PpudAgeLefwVyhcuh4lIx2Ovr
pva/ODY1Pey+oNbjwRojndrds6Cz4bYjRVdfVWAnnyMZms4p+adGWE/O9zrb/biqzfJKUbKgdu7z
F9ORITyteGdMGNOfqW0MC/BX1WagmqFC9PDwIzfHls35EqzxGNw2X0aOzUWiPE1d8ijUjygxmmpn
gZ6Ire+z26Ru4uru6mOV8n1GGiQtwtNIScyir9lYfIDD8vz2Qti6iM5oA4hcZq95cFp3K5uUFRD1
TECyRtn0s8kUUGb4EPDLiK7ktWU+bPpEunR9shtTHfFiqikVkG/J9SmQro+6OY/oXNj1BnJNZmsY
Tjr1CAMA478vECn1keIIYgKKcKODKJTk3f79cfdzlmY9+gDCejsq4LuFLXwCYsSbMMKKQtWiNPC9
i53HdErxGqho1QqAt0CHlqcrswH/l+FcUDMfNdPPegqvdFs0Fy0XZW12kRUHGkDio5GnAZmUA8Q9
iaSBen1/5pZ21biZ6g7/Az69muT1uXdnYMVyvr2z0Gd4yAqaod/fyof7VboLqkEXRtHZAsk1GUYU
kY7eAUDAd6/BX3tj2HCI7F8Akq/eUKtxHTk0r4pISC9GqaHJK/ZmPEN9Y/p0KKuK4StCCdGrxNA4
JYk2psERSQl5l8XnueXxAbkWzjVmQ9mXFm0JqqF2P/dq5wN5REEp1d4aA4Qz+Fi5PvnewtizZpVE
NkrLIGP+m5df8J4aUmdyzObAZ7pMseMwxDawMYnz9tM/ah03EfBR8yOuT5xVG/TJPe2KUGU89+sX
5phCIAGfPYwhG1RQnyUS344uxptlrK1OVlDFSkSggdnSo92ORgyiW8XF4Pd/yjNZ+/P/A3k745HR
whEUmy0tBcoBV+58jD7iaoR3KPVAqxvmWDk44ckNYpT/sod5OgggMqKPACZcO39pBtgQi41KiPja
6IfAGAIjX1+pnL89rWQBNG55l/fnfoVrI1rutmQ+kvgxxHjtZrztmLYZcd+c/ilFzAlP3eXY2WxT
aZ9XyduEIi++LgTmpmFM6JldAPqGdBOCzAzveDDjkCqA18HZcywsCwQFEzRAg611xpMqM1eK8Ztb
66Z70nuHegR4zFhoRrf/1m/2pZFwHIoqIyyKc6+YqS73strkLKBdwIuUwE2T5dFIYDJW/OZe/oEg
3tisoEpnbThD79oK3kNm2IuFOs4qY1lET56i1lpfNvJmH5H367u00coNjG4B8RA/pMMgEiBGzGeX
v9rtt8PzSP7dkMJbEGVpPr8sEKP8oj3LYEil0VCB7E51oGsxC/If/iuwiyEeyCMaNrcoSCgQGP/E
86zygY2lYmlWoJp3cgL2+uEj1R/2yqtyRRO0iOfmie4GhcBN9oibWSoMwLqgt1IH0twMEfNm6BGe
Wd4lCzO9K70RV3gJPCpsO0ve7Wi57PmYK1zBmEtik6d1RRZsQGIC0sLhpwhoKz7DlNmCF6O5AWhy
R58SNeSlYRXV6VHdYrebgsxOjx8dQD5azSfK4fR1dxreHH2ROfrrIue9o32vBoYqoV2jMVCWJbGq
XfDacS1ideH6kbe/qlgtq7ZUrOzsiJU+E3IKSAxaFFokQ6YKuAGBIM28IPAE5k6YWlqjA3dsmbzg
PyulkwcSHGrN3Hb2fW9a3b0IvkRPPrp4DFMUq3oxPYme5PLmv+zVS79rws90bZ7L1fYCwjTWRHhG
IW0R+n8MhgEL9XPyCWVsXCoz2DNj4n0fnbY4fsIEf7CTaFIFm2IsqatHJQRB2ldGvenW6UVmdl4Y
SbJziyR3STERQBukI7B9Dac/QaoauXy9NT8bTIbJ22K8DY4i/u3CHkyWMRpNjnOOPW4DxAeUJIem
0FptRc7NieTiG++uYer7mMG9yujq/5mwzzwBGqoMYMmhewdz5GOeUoRh3O57WQAkXF4t7U3almVq
QF3VXal8Ee9G3nFrj8ca8+3sI3BOFs1w1UVJCRp7gBBSQr0SKbrrxSpKs6Av+N9nWz3P46MDFO73
k3UalIkxx4JK/X4HiFjNPrOBjjqZqqCWZutHrc0oy55hVNilLS2jGR0nbHyoDPDqKowFwqnm9vme
VEL+VI7wDp0SLczWoBufvtgVquTPrlPnULmaIOxV7C8+2ImHSWvYZFRGnoRMjgEH2/eKbI7JPM6v
sOHp/ETVN8gBxyCrDES0PjuNQkRsQThTFK5oRyzLggyOiye4vmWh9ohWOtEfQUB8GLzulLLsN/T8
z8+IiKEoXxE7exuJI9UwQo2aqgMO+ciiyhiO71BBkYbcKw2w+KPSSUIgOKb3ELQX7c9hUJNHAkGy
7/9GFEi5Ja156SZQ8mpCC9NOuH97ww/JLXQ/EmuaE6+PSFybvwanUr2PBz/qkVfuMiakQ0qiSguO
DuWPpPMFMsp1Am0LxLOiMlHUmNxuQ86Ou+faFsePMUbY1EBwhTswbpmOqF3uJTkbEd8R7ZgZKaL6
B6NKO2O5wijpCheky+0QEz5UbSfF9bGbieuPEerhqUW/Tj1FX1h3Mn6gTCXkE45qfg5L23VSF5J/
/kf8LpAhaEPjkxgnoQe5IU4RfFh+p/fFPtITM5/sMFg6o+pwKtvHWxcUhKV3MpupzBUZZsjWE0UU
eGg3XrKcDNLVSJd8cxbvtgS5t/Lefxqg1ZQcArofs2N8dV5Ec7SHLRE87CKv0Fc2fYAOyIwZjx/U
3nUA9pQP0oy6D2p3UP5krVXO0fHo+pkSDrDcmXMCLGyOeKZYdtQ4s3DWHKB9lBiMQcprcgmih0gw
eJfasSkZDmAYaEkwHY4UluGz+xKz8Kx9F+0cIrW9r3lDCOqQkadBP2NriQKczM5VbHgvRsRMe4ix
56jATPAzQmjgMcc9Ug+FUiBc4ccxA6BdbV+DDKddzYWWrRF18ckeNGK9CpmTt5e649iTa/8SqJsx
mIu/F1wUsHnByCKnRLl2PN5qqbKZOrnunNmzzcE25DbJCOUqc4y2DpoIGfblmcWIRpp5/zhG9UZO
pFc/5GDhvhjPKCLwUxe25k7+4s2Unl4b1bUAD9ofEbo4DDNfZM50xl3k4bjZSSqnwePiF0uEzXh6
0ocBKi+KdlwOq2Gt3uw2JFJDKPAKtt5k6UmK1cAfRdlcrPLyrQN4nHO8szCItTB43ChC8mrShXWZ
EWMKN85s6EQscxYw14oXTOz9fs7taSexZCi864FE4CZTMoZkOpstJeSgsUHaPzbzGg2ygjXyNqZ/
Y7wLzHmuIbzC3Lo=
`protect end_protected
