��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l��ӡ;h�>�C�0��-#R�&�`8��2�_E��6�kI�n[�{e傭q�wҴ� u�j;hKb�>�$'���a�찁�l�f�^��xGL�Q�ɸnp��݂L���nڜD��Ve(z���j��ǭ%��H�$e��~~�)��/ޛnI����ܯo��{�k�yl�	`���#•�<#�`��L�C]�Z���B�Sq&�$o6�f�_exa�0���B�\j�kPؙ���wB��z����	��O����?_F$��%h�f�59��8� �d���Zo�<�~;X�d�z�F�4N�S�!�_l"r?���S�L�y֮|�J���*d�H����{8k���*_i��
XN�E{1��и�n(�(�v�k�,������A"P�=��/8b\��A��,�0����<���A,�r�f�Dh�t���!_���X�|�3C��Ja3O���i\#�3`O�,Q,,B�|�q
��nڈ���Nv�@���Q�r�7��U/NI8���VJ�J�}+�ܨ���ԔH:�C*f����<i�CR͔�\э9V.�#�#�6����?y���Q�N��c�oÍ�k�}��i�q���db�-ؙ��&��c���+Y�L�韂g�(
�O_���Cz�q���.�RĲ1zVb�V��	s*���a�j����J� �p��v&�]���H�_z^E��	B.5�(\��D��zQݬ:a2B��]�[���7VTޛXlF�^w���D�Үw���>Y�']>���{��׷�lD��mG���`�B��0P���'t	g,N�?ۉ��>��W�%��g�P󵊘ꉥ|�*Ռ�H��N���� ǫ�H�d��c[� ���4
�w/,z��
�a�/��L��h�Z�;��N���mu��H_�pM�$��F����?�٪��4��-ʫs��w�!;%K5�X�+.��bO D�}�����j}���#�el�;(�ɏ�>Hv�OM5�>�}捿Jia^=E_�R���S2!�������BD5+ō��w�L�l	q�n�E�`.�sI�����}rQ¸mbunN���p����D).*:�� �}�JK$�j���|�!o��XGO2�j���%;JG\�)�j�����Ɉ����j*'|�?[!��R����J
+GY��>�̀gj-�s_0P�g�����Ix����|�YC�ѬC�4�Չ2�X)�����h��3�9�OÎuΡe7������O�A��d���nL�`�6U�t�~��	:6�=Ę��=fC�@7p�"��pN���.�������5�W��F�w�xɿ�γ��W�x���&��U�W��e�;m���@�sz<Y�N��S�t �%���-8�=��1���Ιr�r��+�$������F���8�"�}B�B��2+�t�B1���	t:�ߖ{g�&�ٟ)us��Z�s'X��`���z����#�#eS��Y��(¢���n�Q"&Hs���`F��/���-��Z
~��; �N]|CG^���9qT�+&jr�������R������V�Cڛ<UT���o�*��3�%y@&�픪(�&!�p5�� ���- =�j5����Ìk�\�*S���)p�݈�[�	��%N���������'0 Hh�*����Ci(���`�=�I���ʹ�aHe�#������ �C�/�c�6j:Fr�jwmo)�Eb+�<+�_�������5�TJCLJ��m�v$�O��J�n����Y��R�� ��}��LL�0nb�^^)�'6\L'A�(�����EC�hz�;/���%�?8�x�n:Sp,ԍ�a׹�nk \�C:��IZw�����p}`�7�ä�2�����qQ���g 	U�s��c�k��6IG4�h�e����h,K ���頳%�Y,^^��=�2�^P�	���$yl����!�ӍJ�� ~Ն�?T^��L+Fj$�1�~��H��t�Z�"���+�斯�k�68g[�sB(����̞5g���AY�=ͫo����+$���k���d�&�z�Q~�M�F1'h��\ �i��kiټ����S��q�|&1?I	i�ev��_�xu(��q��zIߙ����Yekq��?���qR���	���ӥA$�6_�e '��L%�WO��ǆ�%����x�k�CqG�H �, �؛�$���DO�Zz����,p��B#$�݅o/݂���'3h8�Xn:F�[�f+��p{��;���n5�&Ʈϭ#���b�s_yD���{U_(�\$}��{�k��V|��>
�TR����/�^l`ynLp0�Ywp�XI��LH_vGy>=�|��7z�A������x�v�|�I�V��!OIԉ��=1,�F��tp�  "<z�̒�O������Fʚg3��������9;B�p+�_�KC��>#�=��a8��W���Y������4�-��>�`-O=*�B\�aϐ� ko'�C���pV�T	��j3]@���$�sS��/��?���.{���}}cE 4)xK7��-��ۍV��o�J{�.�A��[�%&aF�Z!LT��Wj�9�>63�5B��7Z,�H��(ZYx{D�&�;��3�y=�9ۄU��MPפi�I��_�k�M���l/ {/s2s�5�>��`}�NVTn:��;ދw��у?=¿��D٥����Tf��(���y>���Fop��'cO��p
��X�o1	��|E�v�Y�mk�)���hY\�û���%�&���?Om%�%�X}�YѼ@�ԍ��0Yӟ���Ä�R��<n­�?͙�Kb�6l��C���-�����D��w6&�fAy����3�.��c�!Z�q��{CP� ��	�L�*�
��ڒ��Z ����1]�)�y�|����Ɇ��?���w�wyC�Tm;x��f��`��� Ɂ�������e�	"/�fTqLU{��bwI��B$�`媇:�5'Z��/���_.A�Ч�m����ǘo��n���C�o���,����2��JR�?��63[��R܇�NJ�޵b0�R*�V�c��К�(ma�
� �B
�^ٻ�s��XŤ詋av �Py'��hi����!K�cC��Wϴ�:SF�͙�-�	�4������(��e!��)�a� p��&��G����A��r�B�`0Dw@u��'E���C_�r����j-a��!K�cn�᰻�8%}�
����;���5Y�!`��I!엁k���ܯLY�]aTL���B���nE�����̀Ll/_�������Ȫ������nݎ�R������F������7L=��ɦ,��TF;�a�4�����M��|��z��xI����rcE:���#.Xx�gxF;Qyr!�!�!��H2DY�n<7zƹ�-얗{��5zs
�|;b���3�[��_�$��4�>��C�%��^K��a�c.�1�������P��J����։��d�;��
 ��z�f��(�����m� ?�ysԿwI���.kX�Ѽ�q�x���*4l���^� B��N&���Y�r#�NQm�`Gh<J�����r�Ooj��ϵ�7y��w�
�(%%��Q �x[���Y��������0�<�֍n�Ó��V�ʴp[eA������r����kx{��`��Fr4T����U��v�_�G�\��c�q|kF�n�!�,�m��iռ������N�I��Ph�5�$� 2�������F�$��D���氌� fe�n��f��q�]��՝rP~2[��Xd͗�̏6S�HiX[�+J�l���0��	�A�+��
Ɩd�7ey�p^i�U	W*�9�pX`)�a��DlB\Y.���2�������?rT?k�ߠ�"+�s�s�,`HqQS0N�'��z��x�¿v>׿�2Z��2�2����G+�6�����t-s#�9�.�F����;��?��s�ah�Sl�$Ëu^��3�禇�)�o���q�<E)�> uRԎ휋9��C��y4k�7j�w��}�ߙ�iغ�5Ǿ!���m�o(��k��,sޝ7�Y/<v�����a�$�?���f8��f�|K.�����~��-�x�QMzE/C�+ߤ'��P���#���VY���~[�3i���Jf�c�#�t7B�&�tܼ`L�E�_��(�x��!W'�ηw[k�	"�p�A̗S�D��i��b�����f��3	���!�X���.���>�J}�C����aW�c;�\ԅC^髺��]T,s��qf�
�u�y�፟K8�ew�4��<
a5|��)�h;�,+�<z1�_���vO�סּXĢ�$��KN��8�F'�KnS�B��5��g�`�rtS�N�����n�d͇ H's���3PA��f9��g�>h[��8Ԓ
����Ҷ�և����L�C`��I��E���N[�r� ۰���t���_�fii�Ȇ׫r�+BEY~��iu�����y�,�C���o��m�XR\��Q���I�����b���mD\�J����ɨ��	����~P0	jQ���!W*L6�	�`��LU�Ivw��+�|���{�ciVW����Z=��^ku4_�V�EI֟��^0k�}9�{���͑���}>���hs
� d:FḠڭ=Y�?(Q�jx��s%Z�F�l����2۵rT���n��u���C`�ZxG�����i�S
����,�����D�~.�P���5?o|�,��\(E�C�2
�a���?KAH��>5��GV��~�}�/8*�ؠ�����vߟ�7�0��P";���i*�%�ܶ��T.��uF�A`�. h�ؚ(	1��V8M�EV��[HjJP� ����&�b!��X
��~�q�}^��H�Y��O\�t�I�3mIl�P�m���#�}d!2�q 8����*ɿ��a���v�tpQ�������C];�x��uE�5+V��V3���z�N���w���0���Ul�����^�O=+0�p�4<`�+������9����t���r��iF���-P�۝�!4r��Q����y���B�8����M����@d�T�F��hN���Y����^�U��c�So���r���3M��5ҧ�g���­7Jm���fJ�l�0��\�ʑM�n9I�V]i���pAd�Y��@���{)��L\��N���z��\!t ;�]��n?��Z�>J��?��8>"��O1��쨈��D�ҥ�\h�������ϊ[8Y���*�5-W�^δዿ85&��"3�Uѿ�8>�9a�6/a<v��b�ZFN4����mތ�Џ����n#��4&qw�̭�ps�6�8�R2d��n�C�nʣ�9�A$��FN�jv�2[!B&���WYxIr�@��AK8'`0�t�Z���� ��%�Ü$�@�qޱq��!}(�v�q���RZ�#��s�|�<L��=D%�K���	a]��0ɱ&D�y����{�E�j郷����u[��39]0���!��TV+n�n�X��h�.���Ứ���Ѱ� ��Q���?�7^uת�T�" �Ue�g#�v����%P;*w�Y)f6�@�]�*M/��NY�v���dNfF[6���dgȘ��rcE��]"K�O�m���2%��nv��<��٨�O{[~9Dٸ �q�6��~e�4Fc��{��qk4;��1���WN�]bL� z��９�Ρ��$Ԡ)X�_�K��+n����Ew-CAڇ �Ά�;D�"�V8?�����'/{U(���6�K��@���2�gL�s�m��P���Q�����gf܂���{!��c���J���Z��?'��8��k�w):�����;�TP�]�ӟ�������`y5���Pa�ׯ?B�
H$u��;�,�n��TS��Z�t���1�T���衿3�=k�������&`s�:(�X������mpmPg^�mM�9���f�|�>K�9��/-��}�~vx��F\0��3�q툑F�TK���cv���\'&v<���8�N_���ˤ��qB1�q���~C���/���!�6�R���c��ϵ��ox�C!h�XX�aM*+�ft1g\oy~�68��-�,�Jc��������f<��P�JPc�\�� ]̳�� �n�rկ�)��
k�o&m�K��%G�O1�JsY�ۻ gU�=*�N�