// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 15:05:45 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ch1PQTFVzXH5PyIskkukCcBEPby14tDxdaqzlXIuRkMxi2jW9ISsx5wuDjV5irpr
Mkfm1I3oiI6AdKGmgyOv9+8i9vT8Gdalh4Dweup1OK044iKvAsngz+TdjSkdprt5
H1xZD1b2C3cS8JxjEYoD74UrrE+dDZpbPNerEc8x9o8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22912)
Ao70INphvj65QFaN/yedI3bkYdUunRyBNqxEMUJ3n4FIRuYzesRyddc1eL3+FDyl
0MzOVxVe/fQiDsivuzPOf2SllzqqTPzqCXtJcOZEcM3l0AawJxKRIO+1Q6EE2onu
Ywjg8U6BhNHOK3oW6Redx6+x24j9bXZCELA79vWtJN5/GG/LcixTJyjlOdE8Inlw
pq/j2M4QXcIw0wkd23MbhWzhx3WAnELw5XfusC/85ViKTTVfQIgpriXWi4Yop0Yi
OCWVkX+Xe5h7X9izy+dK3vQhwwXTQVPrWUiRgxOB0DYEr0f4/Y4IzxDCp5M6+Rg/
ht4CeoT31MEbicdCyF67U2JtNL/zznT9dt4joVjMwPybY/jMmQIXwAfakuHOzoLL
Kfmxce59/PZzni+JnpnHlMhVEBQGt1IoQgH3O8QMbeQiEzzyRndUPH/En72Bvq5s
AGh3xyXMcjQfDMQKFyZEpnH6mPQrNcCBuswB+C2QF7Cek0MIvr1aWqGqHGBB1t8B
uaMVRTuS4WQiijN71eU3FHzOcsiPZlyhzGvLnCtdrHx5hBifSWU5hje/Tl96m8qE
0zBjlDJBc6OcARkTO2d9u7PiGdn5WwYIX4dBMcp8V0pntE/Calg9zo1MR5bBNJxH
mn4l7o5yib7PBc5y3kV681qYi1Wx5/w6fgKk/RxRbvM3ZMBAHlGTCFRKTl0x4mtc
T6KiHrwqRdrhWsfCo7qdt0dsbB6vbRArXzeztiVoILA05t7rTsuJarXyyhhq/P/l
sVv+K7xRFPRlvxlGx7bhTzzswBLkW+FdicvY3a9bCCq7eTaEWQfCJN5ETOwyj0yT
C3NGp2Qaz5gh7wCGwADTPwBsF0keKyJ0wfq6WhjtIlkdn9cfHtqjAVtNBAn6ugJb
VyIiHmZWCAaOI9aJlmIyAIkTFUAdfI+G2WrLuNbz2SnZtMhwYeBsoAvg8dq773+J
tKIoWbYn9CP51QVLyPxKHA/jRnF4885KSNkCTz35iOuAigryaH1ntJ+Zqvv8brg0
4RVY7nP4xs2Hfw7qXyQpiztmPXLPXL6V5eN1Fr4+y1GsFGTl3o7Bzl0bberURzy6
SB9p+Wws3u3mg2+4dpBAcbyLZb79tL0H7sbxWJO9Om+EVMqcErsktzkrjf+zvFQ/
jXYOZt5Ozs0cRgEqUNWviVVGv+awjTqSfX+OyYrcTdWigDFF/NBQ80s6dg038PIc
FZ6YmhPEJ91kVDJWiViOkyLL7sQLF+c0Z+Ickvpq/wqd5MOk8l9m+9lvbRU7XzxK
pfxgKv6/3UI/1nI6tSncrqki8nXc+coindWNHlyPfd4Itnj5IR/9tY+uGce6TNUx
PQxFaBI0FGKTCtzVNiHD7ylWvA3RUUGtzCRMOvS0cjjYXa9OT3Zmm8PnNuyDauYz
qZKgUt6XVupRC8efmL4+ZN4QHxzPcYCfubX80YWTeHj8FG5FF3BUaceKJNzd9yht
1ENMI6kZPLIhfeomThZseZpmKvnx5FaEErIIc+KtaJVhpnzIzK4hRzE2sk8Xx6Y+
oRiQc6WMKFqDUMb/G0+tpzMGREUooCZIjT5xHU72k7zPMTCLAhm18ycGSY0kzWS9
HpTutjySHzzcopH4Xy/twvrdOhx86KBTDqEXT3P0jBpdBbTuHy0xoX6gkL5RBqkV
6wbS1XmnOohQIUb677Nn4eVbXE36Tv1LQ3UVJRYAUixJpibMHg1X2xoZg+G8d6iC
/L3KgUz/FNrax6/28RaOnZ8Oq/PcYJ8LnaqmET15dSTvID3yKfLPzLSeiD/1chl7
l3P4Ag5vbBQYs88pse2fjzeL8ysmFAPHvwZq3H+3wloabnQw1noTKNn//n7D2WT4
6W5nCkZHr0OvwcWXx4/KXf5GCTA75AjyXu0FWz4cfoPbYbW+Kr1YL5Fajg8JLsED
Q8hHFN3h0YGaclOlnltPiyqxqm5GSijx3xOeCZYmO9FR8TqsawVKHs2EWAKSjWuP
MVOcSgpuTAIrpriI+qUpMq+gvL9t20JOs1gDbORkWTopMu0Bhlzkp6AXAh8HFFBv
Y7tnTFX5hkad1ZkLXBTTfkrltg8Ba2QUPKWMwJiP9yyJwucMaVqVzXy8CogxZwoj
QBiVNEd7uvJtS53YhGF8AFor3hAiwFGM5AI12ctu+vVRf0TK5RQzKu9HiAqo182y
ZWTiBuxOFr4UgWO0+EO9JqfSG9JORh2OzV1CWxn5EKlKspWIhd9Vn+AMCxvJ2Jnt
M5pzfrKzKvVAq1vQBmvjs4hLhKgTMASvTsxXc0GqYwoQ4cin++FFfQV7pyrEUyf3
yeB8jMRJgUtOj9FW9qJG0CQf1jE8bqA48dsjHOvlKUbRqCaCkkeSrFXuYWKH7JCu
7F2JUf78qUwkbSKGmZtT0t4eDAmq16OA7/An6lT2KR5tDl7D+IJuJjP0umHx5XCo
izOI+HSC6TNgJz4Fki83AYp4zzttM8XCPESAYs8s41SXH/L6mKffM5k38edjKwK9
FSTrTjm0JwNwHBlmavklZ76DusR+wIfu85Thtyhu+jltY8Dz52xNxJJKf4/zgBqj
eZX4/eYkAVp6a09ttRwroAxHdko2CRzzRWwmTUd8v4+XOTN48Z3GyvPbOUmCJT45
r9cKYLLAvNveepEWZg52OZK4uir5/50/25ytDh8KqcQ19Lkhk6QE3bhDN9Oi4OAs
xYNsuqMBykEd9bY+W0jmp7LSdznYErizYsRHden6mJU85XgY0gkrRwpulXFiK0xv
KM88h1tLkwdt1A9/g5O/DvPViEmO+mc0qxkomMKSzk5MKjrrfaRefWIu/bCjTZ6E
vbabsQ0jCK6YCPXy+W1ZuYOAaBHSNWoeTyVIafEQaSYhYvUQFPzKbt4dcvMjG3Jz
kXiTy6U5gPVP55IxnPu4UPWMJNoCgkVipvuPDHzxJJTF+2g1eqw37EaYNtsa/Yl/
1i/kBOgb2nXSPOCDzcfHT6DXyZyp80Mhh4hXSee3Wx3xTmhy1S7chcmPz6b6tkCa
DOjuFOVXfXZHsFlwIVGHvRdD+Oo7Ku8ZzbBhO6SZxR8+ObrdHy01qAMeQmXamCX5
MgRMOqx5d5gSbsIipqmMi0hsZU65yUaNl8B6lfIgZMSltcvwmhQIKMwlSUPakEkx
dqlqRgzHIXJq/FIbJKLcqBWa5jiED1fDLECaIBgtKbA5tYHtOm+gr6n2EqFbglyw
67UMd6/1n9CM5C3ico45QhfDBpB0Klu3+lY1PybH7THQi7Jbv31qCC+M46GCKn7x
0/ddWPlO9g1yh/KdNOKMVf3jrF4EbbkfcIf7bDvR/9/khhIaSmDyTELNvfx5gFdn
vfZWejj+Sv4K2pD59Lf8rLUbFjpr0S5B+PY9J/Ef5VFj08EtrrMdo4XHTzSi654H
7/2MMa4HfxTADPmBHLuJOajchyP0p3UoqMuqQEtip/LFTgkBDYRIKi5ZwcbQzf35
3ztYkmlj5mF+WwKdXgb1LzH1xdFJC92yb4AAoU1VhTyvIx5DlQg2tm9+KX5fWXK0
dJ2G480Vqt5ootR7FUes7BD00HVE/RMod2Ok3F/nDi3fsO10mUhgLRJ84uwR2OYQ
33X8mW70WVFMLkBkqxIgdMcG4U0FeWpCAXo6y/BqP5YKIbIEp+J/8BcCBhGSey3e
J0hxJXgdPt6aJ0Ly0E5wTIXVMSWjNlUe8erPWxm+59p9KO4DJDHXYt21HVUR/Y5L
neIBYYVEKV+Mxeb/A0Kb7S9A9nM/nRdQ5GZLmdrXBsQF0H37Vynfo3j4Gr0lB049
EZ15z+6kD3/AxVX9bIZrcuheapCnaHdP3qCbb3W7RSfUTwX/24SZttHMs3c/TLBZ
1vYcYzlYwXBI9w89rHUmOFyDPvhJ22cQpSN/h1foENUsI66BGnJykZGhQ6w6WfDo
YbiTpqLXz6nlnjkco2xo5DWSnkvMRT0KMMXYvlP0hIxn94xGIUoDT3HXC51YdWH2
KRqFBqJH5r4BeFUP+T3ptcTcgY0a1DhhSq6RggmVC450DGp7t5mIsvxDUIb5atd6
g8AsTIztXlR5P1cqqn9kb3zqbo/oYHTjU8xFkbswaKBDiukV+wRJLy41Od/Wnprn
f07XUKUFdDQOg2aK+g/FiUTqlK6hofYnFbsGhUtDGA2c8hZVFsvlPdtWza9qGA6u
Gtz0okZxZ9RYuu3pGt5Z9dcA6UhyZrwR3a//47m2sUoSleBW9EluQMdQqx7HnQi2
qMfM9psauntMN+2bfNVCnpXXz+f4gtHCalFbsi30w524SAcVtVVcerDwKmVllFU7
oWFd9GEEFwSpfFfWrceH79VqtclX66fZ9wmw+vjhipwvVM9PZDYo+SoHErZ9XWWN
q0dkJEel7vpp9NZflKGKGSW8ozK//UERwbQJuQh4pkNnKF9SJOE+QPaiyipMdLdN
p1cixAY2gYxyTb2Modelg5UfU1vEc+jMX0Z2XtiaXMi6/tACfz+xEhYxOIZ2BRTq
w7+GP75cQDFkV9g7QYMlb5J6K9fZfCU7LZx6NJtaPK4Y0wuF9qSJSME/E8YY7Um4
eINuNZ0XCSUFEbp1a/8rhBil27PeIJEdYBOJduCY8U7jjK4vAss5nXPu62t1Rpze
hpik/hpFhGl98HMw4i37x0DbMeWAc46KYYf8tQH3uPjtkM7MW2SieTZoeZpA43KH
o2bRDEq6KmN4OzLFLDM0zy8ilMNh9PGX1N1fVo/Lwl/vnBRk1B3fPeGK2eaTlpBc
CupYcG6gmLHH66pwIMn5i5GLlh2JwW9AaxbCJXhMfVUeCmKlCA+atis0jR6HFfow
Oy5+pTO8NTAMePPZ4uifv9EgULRJppqKJtadTm5qErJBWYPA43+7fa12W+A5s1U1
3JguxtgL4iPlda1bX7XyhMyd5YMgohMhydN5z1XHa4qW2FPf0wtec+JdQQp9JixW
YdDXliiha8zXzIP78diyyTLLdo+x9DAJ8vzxZc/zTA/ifh5yHOj97h4aPlIsvenx
GpUE6BpiI4RnBiSyuxcAp2pSmE7kivKqyDrOZELHAp7jcWQspLZPsBjEDvq6dxQ1
F77ssF6pJcj+jEthoFIMoHfipUBm6NgGVWv3lNVpOVaADDd2cdDtIM9abj9U3hyz
ucFZMk4wL0S9bbRdfBZCIElGDUTtBM8BFGqf4yVq6ibIsTADrH57/bu1sT9s213A
1iAC41/fcWswna/u8bkfB9n8ZF/NyZNctYWMUiLF42ObiS8b4aTbupT6yRUMwRAD
9kpbKDXumpDReMu+O1NP4NitTkqbSuaC+HCpz9OKih9Jk/FP7hJ36pMN7Z9Y2fco
gssFDtaLWclmDPNI6QagPfS2vgkWxBXg1F5u4FvpSCh6GqVj/5BPXJxPNSg4JRr5
35xixFVeyOwBU3MK+baku5mIIBip9XYsDiqBrwyZZ6eCozVPM1jUlHjegtbgnZvU
LTllRqgs2DvW3UCQx7bmrNt/tYtkPJFMKb+VJiryRKI3Ww1ondq9Oh2UWMqisUqo
MptzPZ9z/TdmsHsrq3EJ/h1DyDjmF4lF5m+Ig8ISZnkgoL3hLSWiTWAVXDSstMXU
lcrbOroGdB/Vscj9EkFUF7vGBzZ+B/jzjoxlOhk3pPv4pJijz5Li/Fb8oSpv1ckp
oqCQ8EJYNzIiJc1SvSNM0ZwKNHuZnlskJFkuoi9vrpzcb4HlqNaGas4DtwZ2ca92
trn7dM/+tKk2EQlSNCpRnIbT7wj+T+SO5tO9yr8hb4XuKKf7TTl8+dnotI0Pvz2j
vqdigPpF90HjUDagEgxNP7T7274eUU//fvtG4e2L5eNA139lX5hZ96gaISr6Aro8
7yjPwYOL8goOiMEQ2SV5McKmN9jPIPKR7Qnt6C6FMzwVC9skk9NjZ8e+yLhZezsC
2CmF7hXUWg4moIqiR1RuaIhl213n7FDhcP9pgcjY2/e7E6C2e8BYXcz29tU4MM5l
0JBZsjOhSKA+pOLBQ3p+YhKxgCzOENFAlrO7/nEW7NVdMUG42zZStc0FJFgk9eZw
S1YcwtEogw8eSPQ0xKQ+I1d30TpYdoCkLvzyzLQRrnDz1RDwu/UOiAC/LBejzrev
VSGsam1jKG2+26MZuGGtu7QB0/pOB4+FozDw42u1/5X+nsyEZ+yBej6vH9jmZpEy
eTN5a7QJ2KhLQBWfNJ8HPVe4V4qDUVOYLkU06nY9JP76Ip+FKfdAAoJt1kE01tVI
HTYRfJXD1Zf3RZ+GMlRAG6c6JeIRdiOaje3doPH49YPK+Ne/fFMlxl9XLfflrzoF
dF2GH/NPpWBIYJLl59NdnIA3x35XWnID+GMHb3PyzWEouejqqdhK+sWhJSdC9eaL
+8To0AoSmd/2HDy4plim3ZkyaO7YAZNUzM/0r3dqKknW1N0l5tG6SX6fpq4CrYjE
xBLOZ5QPkkMFqvdJPiPoAOa0/4MNkSvqYkrMAqgl0Nl8xKPIOb7KD3j6WQr2N+5P
wkeCfD8GUIuxH4Ti1kKShz9lXgughFzD/MYvt84M4aFKg+Aoqn2tCsBBmXz6k7ZU
60d8NUtCLbLKUXo+Q34i9j4pMjNwVf4j+xIKzYWDxnKxVjrMvwLlMWU59MhpIIkj
51x1Vv7OmQcCP8OgXxUT2+K7FhqAg+vj2NMhYCkskTYgmur+ktyA3S3oSH5+gyE0
XlSfVURvA3j92St8teuXeVTitmoXfQQRWVJYWlm7OWBlzr62Lu2ddPcAilR80SL6
UxmznfGUJVYNUxALsd3cgVMRCvSGLtICcGyiDcEHooVWqB+DmFP4zUHljmMPOTLX
dHn8iiskJTOBy3LJHvnvzL1TRPJJNvP4JtYsXxdcJosPq26GGqRB0UpPR70hc6Ki
a8fapGWzsCUUvNBni+0cW78doSm1yoxpubTSNC7K46Gmzbz/b0vDZz4rxH+Yjy2E
yMiwCYM2HVH5EfmUOY0K/+UnrZph7mMT6scQC+qV3h6zpGc7p6E8T8u+WhBbAnsy
TXDVJaUOvZKV6LL7hwIF0ZSkxhm5atDLB4zxo0iKBD7RzEGPI+3SH0iiNxrgC4Zw
wIDsXybn7Q22zmtt/UCN/ORs+qwzJHLH1jW1viwMgTC6PsWnITP7DAkx4iaOcX26
9npFFU1iGmUw8Yw0ffVsLo7sAt0SxQvqsx99luwrC7R50gAaHLGL2vuDaBFkvNCd
gS33Kse2V0VR07gHMXsahUBImzw2Fv9S1QbaXyNi3CtaxiM/fIfpg2UeSq+RRlV3
pw5ZtfHRjc5/TyXhLtfmplOiIzJxQhz2L9vOhDfoNozZEoi5xcf70gh1UV1YdOtB
CIVnxUkY2USYsat6Mg7Dl5NfZ9etbOsp6dwNHhpvnQ3C5jLHyzD7cH5jNsTisJkO
5qSlMyeMQBtt4aZ3v8Cm2I1140WyvVe50aTIt+q0+2qG0C1JAElHr6mNNx+FPgO6
vlgUbm0G9n/zmk78yd198KVy3FWkWa0+WLon3fi7x+UqkWJ4xQ/SyRwc76BzuVlX
wNxknE8ZHMu7d6eZCNOVTL2eVKwGjwa3YYNXFEfzrsOT86xRqWejNLDJBL2xF2/y
nbZiEjgtsHWDzw0Qn1UMldJzSt/WFrtPDqxY9bZv8U+VnRivFgCth+r74HtHZ+Xt
8YAH+0lXOBDFg1a83uOIVvOdSdKniItTyBHhzeowgbdnly+mXwLWORO6Y8Qcgd+Q
JaAgcbWx5/Mbz6tVauZsktNyz0tLPhk9XUwk87bOnELXXYAWCC05GeOwBzU3gc1e
zBpxyxk07ib6dN7LQopAodQcjDg/WYW2LOR0J2alQpYD0O6hPxguHzrZ6QT3kj3L
qQkXMfVyEeZ80fRZ99ra6VMGXsPIGw/5SitylSxS2cub2xbiDCxMQdO+sFNVORfI
utazjkWCae37xkTCCmem2Z7w9thT29RfRYoAJjvtbsdKFaPintoJytZBUL4kxzmi
iZjFarmpyzbMtO3UwjVp3Kx8dSg1ow9oCiGGOyztcta5Zx9XK9Ed/c5t8q1ZGvYT
ScNk52aovAcCYT2okW1hvypk58jZxmq7KB2Bh5KfWnzs5JujEY7qAo0t85l1NHYp
AHWnch30CETIwiEoRCdjCrUljgK8U4DuBu/1ROpHM2KdYLg0w7H7+zUo6bITjwye
Hf8ne6WPbYkBxniC3i42ZXEdH8ScPl0MFP8ThEQ+LEhtpD91OnjgicGOLuvQ5vWn
6+a12jtrwIyTv8gsLhWu9k2kW+1avVIVd+R/btNp6R7FkiEHoK4Hu/aDzoOWCP4x
WfaNWsRhXrqjUV65p6UXkRcwFYIQJ3dYG6vgqgU2IOMOrKox5ulCwAkjVCex+1Rn
D4YM5Z40Yz5w6QoL5Zw73I1AHxZmVEHR+5adiK2GsNjtlmgVUW1UCwg3kEFOhRtQ
U2/l+eF1ml9GlJ0bKTz78m9A2sA6sTnzRTUbx1pvlE3oHtzbOXSQdEPaCG2qu5ew
NyZX0EhJQl9tQfuBf+EuZBmhr1XwLk0aGrN/85p0xAMAia5rh9p+XkjY/WgNctTB
UDKIad2CFYoH3YYU8hhxqkhqtm2i/aR3fgFXMjjwVnlR40mUbF0SJOe7YcUkFWN9
ZQS1Qpj4v4RfvlLu98QNwr0pLT3KUlG9ufh8FObuSfAHMX9+RmkEiArfyksGr8Yb
uABkTc/hjZ/3SZVbGEhphjZPd/jh07rHYDi2pXxxuchdPwND2D9bEdV10X54EzjE
zVwtZzBH7J89VuNlXtmd8XfwhLBQcigoU+1mjsqCjNqsw6brKdxZSyDtK+dnWlFl
HP3/vIYjA9YfZRQLYJx5CN1CdVCHNBgqLZGv+IKjDRWHjt28SnlHxXGSRpcvjhVM
Na9Iw/xqWT4Sm8XrYXM8nAWnRrxpiEExTx3mlMobEZis4fbHArkEHKX1Ho/WLS0+
0uvJYUOiY6BVs0X11P09Ncuag6LBqF6kS6rUpmIiORj2RuGSrSm8L+vA5//Ll+Ql
gWtG5jyHqNLEdVSCbm1MPNnANPd/WByQugJziG1UdpTYvOZ5L2RehQUZEnpbxl4t
gP/Qn5nB1ZJp7sgalf4n4E0eBjSTHNlqTREkZRveqMtkcmrQFNiVi6xNJCwZBssL
VAw9p17SvvL/sEQRcy7Nr6ZWTMD/Z9DlzgBZb21iJdgb1IV5hjCc3PDm049pfYv8
0XuHzVaMR7rZ6vjgd9bgh+1F9HMr/P+MDrSmT8GIUGfQO1oj+Oik34tQqA0TKOft
PJq2h2S38DDdkuzds/Nc/wE62kDZCkWhAoWb6dsrt6LXPEXwH0v3m/Tq/hwsdKh6
IL6cmOjBsUQ9Gwvfln+0lm+UN24iC08OEeqeI3AaUNI77Q18lkOB8Mnk1y5iAeFW
7980mI+tkIYul3+/o+DO/gLGshtxIzQiS3D9MWECQZUsuAXpWvMlwNns2r8hHRbX
z6ybLJjsvxFK2YdoQg5fm6NtqS2ElUKUcc6uQsOJUA7j+rO7Fiz3tEa8HcDpJB9+
nFunvDg3rWpxwDXZAmrmSvkXfVzFl5AJYqZyEVEtbmh6OpLghesjfMeH0gTpch2w
oFnn3rDF/5KcLtQstgzpM0xsoaAAr4xjO5TCCux+lXvtDmy3Yfk1LJyJQsKZFh3Z
9LWbVlldn/UmYkigVG06cEdrs2X8MLpq7qdxO2f51bSF4UupYxyBYXDidMqPuILH
pXz4RKGTcedgy4lXyGCC0TbVt2iV++cj1CzmHPmZ0TI+W3gLbemuDqn5Y/5r8nQl
XSif17WgK8KXZub2YDNP1DPiKxqXRDHNcur2vh1I3KyaK/SSTbqcyZ93H5MAwPan
nhFHONH1QcUFW5lsQMjYORTmDcOW+Pbtu62JajUGI7WgpoSdUn9Qq5lVTDkqTrtX
PuuiEiQQX4ycW9FDmabPamZArbUlFH3ycNjeZuOv1KSX8D0VmSriktG0mtu/sizi
oVYk62skZ+EycuwbdjQD9SU/eJNyBe/z+1JWgYTDZtT7+FocECznDAuPL+dmE5es
PXy4Z4I60vKElVtrz2Lia0TKmEFr5JLZ3WHdBVaFDPq1dth3RggyW83w6MRRPwzv
1qljCNmtOh1gwul86NQigD0XuHp0g9LEdyU+BaTOZ0s/dseAw5lI5tYpNUpnXIQx
Z4hzc1YmWgIxpOGoyv/sLESFxhNkWYVpJzwyHPcRZyqsBfIUxhEMl70lRkxSfNn2
lvIHemJIFdThaAV/yrrFDUfBTiUxuGMztMhse2yxKNwxYMH2N4xa09gI/rStom/+
eUaDH/1KISGEBdQpA9tYDCV8y7zdhsFRH5Wt5gEWDfI5RayPBDfAd9ppSyY9lXmh
+IfSjJreSlMkzlq4G+nA1pcq5hYh+fru3xSrTNpGEw5lBpSrda6fHGzUuR4zCDOY
2OxnLSszDgbRk2j1yR6KsX9ZA8MOZDFid95RXJOUx8bemScUORlA6eixmPegbbrF
tHRhVJMAFAVVunqINn8teOz4lODaGwGhRC8tA98CjjtzoSff4MJouhYucWZliGg0
jiPRh1AZ5dPW/LG7IG1gyTAipX9ovd7Yte+qlfoPbKd+8BIA7cB8mv7i7R7SvYol
FJ/dwaDPos4DTf0V27CMh2u1B+GOiGZQI446p7A7BDEO4SGmsWPO7BiBbbmjZeO0
7g9uZna7GvQwT74nxNberklgaVJTd7uARADntRtvgkVwkQE6h8Z1yz+G2wXqNOgE
NwHP1Od4KbWoPAXuvTRQ3TZAQr1eJ29M8+RB4QWXHcEUB7phVmrAXplp3mqpyVL+
on3B4A54ZShvMX2mKy3R4RQxgv6sh1+T1qzOaIZl3ZG/flsQ3nzCFXanB+iiLtWB
XyFyMADvdSbhPZnVWzB3kv7AcSMdbitIz0EY4FoQ7Bdou0i5LzUKhhsQ4gEwAMK6
8wjqk3cm919hn8nmrL1aoP1ZIYjM4W4aGC+6XnNUcDuwxvPYNJTAlGGgQwhwhJkk
dbU7zXHslRhbXpC1INGsTQBdFPPMWKNAKkAo2Phb018AO97ELvlD15i+IJJ0026j
7amiiQwsPen5zUXn58vwFPK9EtKmWsUlxAr44RR8+fBDuU+dNu6pXNoPwkEoxim9
D3ksj8hOaoqkVG1wMYzpOBl9eQIztlk2U8Et//923eCsF2FGXq34uCCC5lAyig+3
/RyxeM4cbhI7Y29DoD1iPdWqpAw26tAMtQ1WetymeyUWOKzJ6WniIedzCet8iwEC
bGvg7uN0qWi/TpASbUQZTpPkE690DxJHOvjmUflr/DbyTFviBwPqU3A4W/aPo97y
7cNxhN0pbOMTqf1fwUk/xV28qUE/fEzcoZcveHUiERZYPsAPpKatUBlxJOWoZBcC
09YI5AH1nYGWhrPAfggKl4t8skoaUISEZtpxe22kyJarfIWZJigVmrHuF7dhQwtW
jYL9STPQi6UUfG/EIds8LLYdsKq34TmDtnPnIBT8lzXrPWngEHe24IDtiJtM3JdO
GeVd9Z8JEva1HDf/dvoICfkjMCzqWgSyupb942EOJMt8p63Id9od6Jb3jR3RxLmO
c1diUs3HxpiQyjzSdlWCuF2iRLJ13w61m2nbVkupdxHNmiquJff9EpkDKk6CWaBi
mqnPeomhqX1Qgq+lnH7HXAo3Fhhs0vMpYXTAJjdCud6TfDjErykujoVI9xIPcDJm
pCiXOJ43Vt/jJNlHHfCu3NEJgd8mXukqRXtitDP/GbQ63Ga9ZyA7875vnydumvHe
t54bTKR3NfmxJFVGVqovfymOWldzjT54NlRbMNvipoNH/kkVOnHniyxrGreurUgK
nHzGlDkyvxJaxRXJGghk+hg2uttixjm9mojFFGJdFghe2k30bXPHvFTyFBDBU46J
6IbTtmpYd9ruMkqtE4QIJgNzVYeUMn1UagPMus2fj/1gkqAVSRd0o8Q6WzChvGKY
SMCPssd38BMcCnf8qulGNTA+Dhouu964+dn7XC++aDrF3GQfv6SgF8LXlyt0eC47
wifyTxTYcPaUEwA/hUi5AngP7JcECu8yc8vDoQK1dfHxQsGc6BruzaF1MeXssaEr
H0fG7vWbEuD3FtZXskYGh45M5clMq7BTrLGhrcctPAVj/kqAFthu27y1hkx6TBiu
ttKRUOnuc26Vys1JD0k6A1CpLz4jv79o+DTC1W+BpCLE7m/NTTw49WeF0kqkFTRu
1x4+m+zd6TbTsCp+duMHCUVUfWst02qX0R/scFtx2siHk4zcfsrTDJlAwL4GW4gd
zCjSvQ/xfR9PzDaeCH4LWY3p7Mv5cJteIL2CKSc8c/EWo68AaU+Q09umaXN/gYVw
yuqW6ClBb3ywqTXPwwl8/dLrDmq+wMVI2RnHj0lUqmija2q4e0TnaZYhzjQ0QZcK
IjZq22YHpcgHKD+34z07Hlu/VsbBH1ObIuH7WxhfAJ8NAKPq1vW2BmQusGam2NYV
MPb0AkYDSUmN3INpBOhaYPo8PSC75DxtzKsFvMwFN0cmioDbjQvuwJL0oB27OnSh
l80XKZOUwsGnoA6vhA5z7/a8GcAy/vJKdi07qhXYel+AP40vbzenSnvl8ovumnd4
IehfpMuy/dmEtAIHE6ZhO4PmmS/rI3qC9ZPmXWUnsyr8OpW3Nz2CwYJ1khXbIogb
990eTT79Ai2OWg2bM1TThcyavItPbprezYvCB5z+qnmbmN+k26zyT7xlxAMaixUz
y1ARyrQ4MRinDu+HbH6jcthXmj72Q3j/AdrEi/VmY8f8ehlf+evX1kmeX+WP5/PS
T0i7Lzh9nd7oZ6YKgIuZfIuRbX808RZReIF7qGMizTbCxH62OpvbekMG0m52gNN5
/H6C0CtMc2G+AmJ8mYVMJM9MSIlL4KX74LCZSbp5lr3vOuP8v19SO5+j6qlFkvHF
HtU3HNBWziUPZ+U6Jks4D1rlBVWuttKpJiCu0h0A+dV1u+IBzFnyAijF7b7jrPYi
+IVmRjxqAM0EiClAMX3ZIwd3AQ/oFzUBVDTiEOuPjxVcYCMsXBselNWy3XjkEunO
up42EGZmVe5kwBCdxmMgdHE2sl6vS2lnxwdHvokGO3uSz/mo9RQibgmOjq6vyrDA
ci5jhwNrpCJOM+QyF6ohamLoohw2UoeRKDpSuGwffAMl5dSAyoCOaZAlcXxKkGuf
K/NfkzT0DG6Me8brDJ6QGbi2aaPFYIq5upRnq6ZH1WJbF2z7xZz1PAcOB1ZqKWGv
HugpTgyIaUgaYMTKCKxUyuLnL3jy1OERAXC11OOIlmx92MZS/zT9ZR/l1rkxvlKP
YCdgBi6wiiaQWPjCv3I4H2HcjmNS7eNHpMhvoas2nUFylUQIIHe1EysmHFUz2thY
BsiZaYyvb7JlZ/VnEUIlguYe2LiY/02mHQ+jS/3RhosuI+Q2ICXxyr3Eb5Go1MDw
OxN7j6PkuVc28pwYI1GhpTrayErFE3K0suVIbEw0/BKLsXcAT7tSrU/Nmz6bacp5
mUrRuqKfOVlGpI7bSp0XlFGmn6+qdm1mhGhD9kOoN3qdrhfH1NQWVtghlzQ4lIPT
sdj5IlQuFt9eaHg7MUAhyHd9iH4ctRkRQnJOvLKb8b4DaxyPZm+CIVnOt39eTBBG
1MLSYgogyg9lx4B/KaiSfqyQhpi4EL1lvfSABdD9UMyJkyo3a1YfVSER+TcTfAng
/Mt8P92nNpTlu9TsfNTOzd1nijjHcv2cWfnaZc4eJlH/6qtEr1GoecXZ13xZRqXh
uI+W7UOGq+zrpnWqBy75v9QWV/XCzVt2Ir36w7qPw2L2/CV0TY2abEi2fPEIxz0p
oOV7uDEXrgzWw0kKFNcgyvTZ1eNNUqYr0Suz1i9wQX1H5254qu81qd8WWuemHVBH
gNGzMgwllBiitMVXcFXH1uwiI2XP26XvGBFC5Te1tBWGJ6pOaen1QTDWFL0vmH7G
nTIa5llt1rjg80du52W4Y0eNWGZECTXA1it+bfBElZrJfPyYIJiYz3aJpA8mhaIQ
uTDMLkEmZgW4N3eCX/lEVsEvpl9LzAvTq2KMgmf5OnmKZGDyQoS3PTWuNl0t/zyL
+Bm1zQLi7hwHuuTSR8JluuAC0dytgzQrZQ7FbLfoLXrHuOT9dIGz+NY09+LwErrO
KR6FnG9+c+xzwl2lKqVwcANmxA2R313VK8xr7YTRtcXYDabPh+EguHMPoNnhuoJT
5aHOa/BVEHBzKqSU6X+WA9aPsvcScT0iZCsyy3RBE+slgyWfI14nAvD7fpiMjCxU
tJJT1hK1mRGMUDuCNvqsmsZVnOutmlicthZgrpXSZq33ov3ENQob1GavmypxzkBB
eOHIdoh1liIwhBSh1BBmUKDqwhm7CqYd0jRfViqcDjtOPX3YB+hDUVy/tIp2EzOS
JTgk0JniU5/4ahY1UhrvVe6OyzEcdiiPFPT/cw1ySUAsYrU52NX5G4rVqm4s/N5v
ECNTHiwA6coSccRgXMU0MIBpRHfbKg91ScDjfy5p8M+WrYiEuffmcl6mevHbsH9P
D5+ja8eFuL8oiTJ0s4Ei04QjyEqA1Hf/GnI2hZbS6Jk44DWpFnE+omrPbwFxVc+t
4F4ojIbzhN7oP85GlAIm3Q1+nxMlATAs1Yy4r26emO4NGUzkJcnEWVVeIlyq5CNS
9VQpuYP/dxaVRdXr+Qc3HkwMrjyvIcVHcOu3++mKZLJxWUJ8a/Q74Wk0EEJLyCa5
4j2cCT/Qe5nSrUxeKPvgJPDR6UNWqzkME8X8ogpjKy9ZGSRGtTBLnZ/jV9WpxwVD
xMltoXFc+0JtmdvV0/YwL/+4v8v7ZdLHER97I0pVpZ88jf1dQoNnlj8g26N5E9Rb
3r/Nx1rNsSrDK6jHkHanF161FHpwORHu5f5dj42Eajsne+VJ0mGkcHcCOmlFeD9v
ijLMp2qcHPIPGmPCrFrGZZO6UkYO4lTc8HrtHGSafeVcPR5K4iJITxrvCDp4DiV4
H6T5DBsg3m7I3wPTrQw8dqenFI5sr+20SuX7Gvl0s1CYsHethg7k8Pfq422Ccr/d
FPcq0a7lMnL0bdzDn7WqH3pG1SbGYryumVsDel+cRMVL9Kt/2PUQ1vU8O+YGw0ol
eBolw8dNgi9ElyT7DU8UeBSeu70BeExSFJFm58Lnel2yoojHNFI523mV+me/aojD
R9fOmEYk8Xfw5yNttYbBpwR06tDPfQk9mkWdbxCDirGDmpr+I2mI0FKH6c/4KKI+
DV7fv21H2WZy+bGiJWdkf+YwDiJ7N2H6efIUcdlknTBm13U4q7ay9xQo60yWXHyt
ZDRfX5d/JjpQUcsVjdO05WjVIa43UrBVVoaA2/rZ7Y3oD4z0Jfd+n8InPNWtAncc
r5w5EsIipJPjILCc0b8h8cBvIxVywmhtCoYGmpxeGyi9d/izj7XeLwRXcI/73Qmd
RikLyCDsMPuyhQ3zKi79J0tleChAsBqkaQk8v0xWfZx+r95CeGpVh2fzylgRWrF1
uijTrJiq4LQTO9ZrpDNFbHl+KgU2vDSxv+HXvQNoaWfWE/ujjBk7/P5GmBQtrL0V
KhBuo/hcRLxp6CYOjYORy5JFA+QgVOzmjJod3ZXYTlWyuUt1uwsp0S5nEaTjYm84
0Xxsc/uLLiC7uzIzPpjld/Qkn0J/awdwzCOXZ5IalKjRPLkK2MK05XKMcCJwnsb0
DJ/LNLMbD0DdVOrNx8CyO+dHBP8eqqN8gtBT2X7wVOR9hildiC+O5fACrAWl7PJE
pNWUPCWmQyrmAHCSc2dBNHgt0XdZxS/Jsw3lgcKqlN0nkC4p+MbrvV/lstZOZK1F
DfO0pAR+9UKtDYe69m9YJ47OGJqh4WflNxHzjbGtq4AHNcKNya5vV7VoOyJhyQ/A
xoSG9g3OH+2+IH1jU0H30h4ClMX9OIuEVvHRXwxaDFz6URo9hvP5zoOFDS9fvlun
8hXXDAVvoaH4q7FwBzYTuj9nae/Y5jQNVhZWAKhj5oRvMrfsVuWZbswOVuesSEUg
TFDw+tQid3qwVWZRj9etgW9ySTAOi5NNDPU8sAB51C4dSS65YyDuGys7ZDHiSsr7
QzEvQVAhSZ7X4/reG2Dkhthi3X9xvGms/tC6zsXf+h2YVJEv3IHaiEk9oGFCdisY
pW8h6yV7ZooNc8c9DceMmgVEMu84EnesAKTLSnhMAENe0S0/WQMhr/o65no82TDv
myvN4U6ZJlVhBAmUr7dlux1F3CviYsJefmyFqbg/dX3zTfn+KAOb8EF/Br5Aer/b
9dD1T2TOpcz2DztkEizF46SyNsKnnNhi/qoBwlelZzyE8MGFM51B1Jy+UhtqnRJk
iuUZbAag+0L4DW2m894ujjlERCC7+cCKe4VpOL/+oIa5wIbokMYVmJKJlKXPgSfF
OZvtsPwRnA2CddcI/EtBxjIuE1j8O46wX8uHsr3u6TtlZD8ikc7i2Cpg7haQV2+3
fPapWaIu02oWH1hhSR3MDB1cP/FjojvfhsxC/sFb/iarXNL8xjupsC7vCqX2+Ri+
I3gGPO1z9WJuTImS8fSz7xzYYsc6KHamwB1bVn+7G+/ARsATvCJgTZCm5lh82P4U
Nb3hnpwlIoTzvZFQpxx/14BRujPjdbBAGXQvrNxucuiAMA0whphqyp43TlNZq68d
zteBh2UrDsN3EEeqr+DQ3eTH9P50EomKfzwvlnyJSqchA8XYKaTZmjDhjPJRYv0e
5Boy+JFaPgZnCCyToy3sAwJ69SVv4p3m/yV9M+HuXd7Mf3RPP4k7O75GKxNpCLgl
rMBBG9qjqoHWODgKaYrPPJZxjJqHY1KRUy0JBF5lkoJXt4CPNI2u7VjDp2ZPvHlZ
d+9IUKfp/ROp0vj/XIaJAfuLo85YHYczVWnWxf8JtZlAW4oFjfXXmgJTwGRHpQVZ
kctlFMCyP7SkhBjb2h691XnxivGbQBgebPBbk26vZZpPdrMbuWj9KAkKQYsl49a3
KqHGbVHYtFevcpR7CNuGwqBjDSYjT0DyW4zIpR6ZOuGNjG9fDZgJP+I++8SE+S6S
j6xHCRgxMO9wR4MUDhGy1aijQakKD34ivNB7zwtj0uuDb9XQRTa++F9fg2hq/tHI
r4foBa/g+JVLD8PhU9Ua2E/z/kELMnPTOswSCaX90zeanQSJ/NT/07MQobnsVoV6
nxyx4HsTLp4/kaA6zqv92eHCy/jpGkf0xrSUtfSTk3DYiJ7qkxilT+BZew6bo0rz
mLLpfk+Cv9n8Tvvdz3unJZShgWrxRaz4JQOi3p5eSOGE6Gxv7sIuPOTq3QijV5Lr
MQqXOablXO3yAb9vV4VWSuo4p/rjdcWl+samfDZ9lZOtuyMit77GgYZnUUsgtPcM
X/k38RMNd9bouvbH2nN1YnlJr6o1I41+Ka34no9RC2YBX0Xn52RB4Jv3qylCHkzo
CxWeTPLqyQ2k5RTv6P5qPtVZMAoYfQDhBDBxY0jur1IlgJnY3Xc7PyCXbu2dBS/d
cHQgqh3u3hGyNY6BsKJcqSGt4IW3WDaEcIAA3gayxAzHQTPmglpdKrzD8PvB4gJp
u0+WnrvH3yIEeHLTGdFO8hcLvEbg+bF9yJOPOIXz1VKM2DOf9cXljWh1Dv16nOEf
RVXEQj0weDsvYesWvI3xn86TtW2qmAR4mvfnvvD1NWJ1mgW8F+5zbWRFTlhst6H9
eZuwUuVh9dJPUAI+BeMLLJZrTXTNEbwgIG/rQvBgp49G8YEV3lh7/vwTC3IPs9gn
8VQ4DXAemhXRV6FuQ5vP0rgwWN92AiaD+9yaJskQW/u3VqJ0AXdXv5TdM3AAmZ8t
1QpHAO/qDLfYma776/3S6httkpRQg8Gg6kZcMkNvNq/epfC77C6WxEC3/HW2lpam
Z85cnt/uGhsjuLZoIEHvKM3nbLKF8Gl7J6PUKxlpQOn+qgOlj+YiNYzrX5+/gzTF
lUt+qKpvg79Wqwjg9qKrFkvFptH1fzryOUjJ4OE093BnTEeZOuzXS5xsv0h/IxjK
5UarOs2p1ibqHLLFNPWWsgCsQbICq7QRzED2h5LpdXU4rkt9OGYz1Kk+GOEkM4AN
Qkia+Kn+A8TjYfx3Et/xrxBiSOaqOmMhanD37icLC5KqYEVxVSYZuga5JWr6PRU9
qM2LijyZyUXNJm7WkEqP+3c0zdGUxSkllnG/OiePrUbJ5Qmqx11oE0i/lZPhVDtE
oOsKlq+uhBJMJFDU/MqxC3f5mw8SIz6y0QiZI7XRrwqbZeUtxy7FTZfdKC1vsJTd
RkH5QgsLVAenYseX6Jtq1s/n2a4FOKejGpcAV1AoFG6NA+Vc4cv8tUq4yYlTLKCk
ieCHhfdgwDhWbFoftpXtF+Q3rR26xGHyOTLRNX3OnMGNaC6L/3MWf9iN3gwv5Axc
wLeoZQ2LlrNgHkLeUgR4fYY+q4s0OLyOiSLQkV5vIVKeaMtQeUWq1aROcE3yFR57
yZ6faISXZaR5KG1YiDqWhEblmWmL/Ofnsdx1ri/p6WhpyiQkvC4KqjaLyI7hutNR
/QnmFu/wOrcJW8KaYklaYA6F7YnuLuYw5e+MDuyq83/vvJx2qSCbqPWkviEfeeYC
BN2BvwfdfsetCXMb3CDe/YNdyu547Y4R63xV/S4MhPD03d4z6ncFdUPR0upkqXrh
PbnIS9+jdoHgQFMe2yXMJirGyZmrEp20JwOoEsBIZX2mjTUX1jP2ybGRhIxMEnKa
zzY3guxvb0XLcVJBX7Z353fcHYnojJuc7hCCFubakq7KIl43gkMaeJ71OSYIvaWG
L9+ZDfUUib/RC7sZmZzlF0+NX6VfDKL2h3iaAliQnNCz4izuQ8dMCQyaFn8LqAXp
roH4mT2X/PAJoDLKGnltv4BpzL2W5ObwOglt2AyQ5O7r8ExxrK6p71FewmfGQ3mp
9JFCOq3ok5l1IjTIYvvfAOIMhM8HyJmc2zNeO3MND2DgU+4NBm5yW2t3bE4nLGBB
Bs0/irj21YoY5Lz1T9Dily3S5UPCvjG2JfuuPjPVkuKNJl56gmLS588AYxLFbP5E
gZO1OxjkwlayRz9O62rDNEODrLTX/XGV3YjWAJs20B/Z/oRP+q/smJ7IfScslDtI
CC0U7Cjc1ugYpqHtewxk0luirDyRISuiu0Sup1Q/MNNXhmEnf/IrR0nXfuyxxNnP
eBdTuaDiW6K2g38NJY4pYXOUyioH5qPuYGSX4hGlpLsuIFli6mWklMJUl4JkFd4K
9+OBY8jgFn/Bjf5Omni4YR9tJe84TpPsTviSIKXYqT2DLNLV1LGg9AkxAvgKFojl
HbIg29t/0DBdl9AgacE/3Z+8cQs1Q97m0/fZ8/mqtdZJnT6WyfHKNbalMrm++BWA
XIwG70G5+ZGi8+eQtc2T0EREjZ2Bt5Kx2pJVmRUX6ZLTkPfyYQLbSY7blsvx2BMD
L8+YjetYIZNwQ+GIy2pN1WgCcZP2VkaLuSywAu4zZ7EgsU9EjAumlKgNaH0rZ4wM
6IionsoZVSb78fYYIy9s1nMNUyC0P4oUebIGoHtXTqAEdTDLuxGrPzUynoIYxTXJ
jgOn9EUpGNTR9JgCgg+w7GgxOsiR38CN9vW0NcveCWY8e31GlPyVbJy9QpOTuO7X
F9oPfhBf89fUQw1y93iNUCR0RgUxmfRei4JDfxkfMYYXTlRYfvQSIBbShOrQI/JZ
wJrzFM2a2ZEZgLTTlbmNuCJxI5ixLT98YNlwJxxDF9FtiLCc6J9wyyWDh3EEjPAU
pzgb4mIxdlcYCCDWK3kLppE1QbivMvsEICkHbx7QsLRpbABlzFgqSR3P8nGmSL5k
wL3yeuDMMFXbzv6LN+2+7F+0nfn9IBQhXNSU18CeRmWZelf2f3+V0ywinEO1sJWK
n0LPjU4IL3EtuDXB0TExj+kbYHLCJ71oN9CT9ZAaIBCjP/baNAnFDqVpD+796knq
+p7+360hz54gVhnC4P92gnzU+g4/oy6R65o69E4XvwjC5KWm3vkrAQgsZgLMY9gd
0x1IOtkrAamm4rMi7I+znWuMIKomtnWAhhhc/bcwj+q508k1cUcCVSncsb3xqMGO
KnUyH7tOZwlFYucogCtEuaFtju8PhBvlWVbc9K0RzqX5oeyPCS8XTmAxK83dTcaR
Pp6zQbCZlnxXA+tFtLebnI8JgUAW8RMEhsObIQ5GpmYKBJehDky8xZ3sdTdzGYZx
IDcEGycv2uvG3952SxM49e4MY0tUTjZ7UHcpCQB+m8X02spOE8UtZMZYC9sjpHTV
XQv+FIF1Z2g75z0jdMx6H//4309RkKDSsNYG/Ud/owJHoSgmAM6B6aYSjB761akc
srWn/Is3/3FBvMKOjXU7MBql0qBmshsTOeug0eRE8lmO7HBbTlgcmTQcN2o9m1wq
0C8ebqcMI37D51XjjLEwUhPO0boLGaXsgqJcQIayj6zl31/jxUB649S5mM2jiIFe
+8rpUvrS6SzPdQo/aCVVlnLHmLTs8ayRMeDFgVnLe9XKTYUnKwb61MY8uPCBHXqN
2FADz8qabrtSTivUZyf84ttWdxd7l8eSCIDLbdkBQ0JWQXCcCr+nq0ts4hXtR37O
eGW3ICJgk9PUk9Eia/y08nYQgbWBv2ut0brgrHvf5IpM3EgTpzNPcAHXi7MPct6X
tRGFlXludR9H8tp3dLCgSKfceiRDTUDty5/V/gAH/JsXou+Zi7Y72rOP4Qoec9B6
4XLrxY/io+hqmjrqAzimXqqq9ozgzo/+x8xe638GZmyCWHjP3SJn+deo6kOe3/Oz
phUprkhJjXaVz5hdeUSt3oEqqPs5kqHHyvMJc0x/vk2poeXi0Zuxt25tGRzyv5O4
6GXtMjS5wwu9sNuDNshuf5fHCnFRwBVBA4VmgI1vGU6ur3Dm7Sl0qybsZQQH3Rl5
9zDmChM+WajJkgRBnDSmIqhD1c7kni2FJq+3nN7Y1XvyLWve72tKci8/oi7v731i
pMuGp+iBIoOHhGNSRRnMQo3nypkGYtilfU43G3/7XBIVGQjOvYJ0rVZb7GQI6j+n
wypvwtFq+8aAA275tiTopPoZIFj+pPxzC+ijx+qqxs2qydhhcDcTyJRoKb2xtiyC
83OsR/DMDEUonz77rgedRnsDOuehDFmt7zY/5em6SeLXg8xTMrJPqP1xSs3trURV
0Care3GqCugzbmP6MJCtHKz8B4w4JApbB+czNaiUnVJQbWt0ATsKJZJpM6gGFgJA
NXtRxnK9m7j4sSuSuE/ntc4yfe3/bwL4mr6E59Pu01p8rcB9FsCjI6NI1NKWtV6B
mDE/V8EWJd9MwZWXcrHL2ptbkC8JnlxNu0gZkqt3jhUaFvxSdaQ53hW7d5JwfTUp
dxxQOJkWvERqn2PFAAF/lNBMvwg781WzbalmYvOQ4xrkco1mOZsYs/GD53uHt13W
gHv7ikNndK7zfCFKqHK0qCqYwYwRzmEanNzDiFteR01uUXjXflEihW5TiWcKrdH4
pOYfqJkqBVqCL07bdK1DKsQIY4RvRBEPwzFFwpeDA2meSiRRzAwmAtgyF8chuIlm
UvQ9d+tksUzsX7Z+UW5+jjtJ9l4QoYbKX1zaO5r7sYigiZ0adDfK5IAoXjPLYbLs
X6ig3s9u7nMoR1AVp4U2274gs4mYgy6tAsmHZnXqMPs9GHM0YHy12WCRbRtLEiMW
pf15QBYKl/Cq2zfkzQ268oiChvIJ5OZXiENSa0rHWZfYUCz8TaauKzbjaM5CC6d5
3SfgyZ90xMrk8kR3hKy4jVhFjDVT6MZrBVy5CE/+84rsP/ZRryDfzl0PoBVhIHaj
jU/m6XpUIyHl6L39YMJMehbGUZ++lzSTCXW449Cb3SnWdOoVrTBz3kBMn8wpVKpm
HgQo5MHexIIohzXbLXU1AqIgkzgAmDveojrpboYLzmJbaD7Q5hTN5ipfgtyEDxlN
KxZW2D3BRizgfprIxowE2ETlOlm9BTeSxwCc0AWe1iLylHqA5h2U4DrJnPVJ7xyb
j6RVzyP5MqYdmGJ2pLXIG9fa7aHa9KkOI5S3d0kKfU7327cUcI/5/XYhflmzCZKl
OpDp5vhK2y+zhMp+mOnRz62EOWj4iYsvAAV+oQjQOchVFxpweFe6Qkcl/j9Rnsl4
jVo1ywh7sj3f22WeMsX8aZSzCrYhYxsvFXaWVglbFlQP8bTHSUG5sbWW8mSDYKZl
i2SshFuA4OcwNsohGPZNpV9NlX7ZHEb4uGhkpyGYJMTg9aPjdrtfePkwG/YQIYgD
ULgI/bI6JBrfkjgMDv6+6Vy37fDPMwOcNIO26aSjGqGZiB4UcaPA2TfOQxniML4n
GW3Vrz3/hnxJCYDHOgPlGOPJMi+SmRKxAszydm5ZYyzSlmnXng6jA3zLnkjiMIQI
glyN14Vi8ReSnKDYFqc2saseXO+IkpXtrDKQCmshUGcOspRipSEn4+WJN8V57kzh
8nmkCp0NS/TlZPIepz5JbqRbKhd+RC6HLOwFLCdscjyuUYtRiLk/F4auURq+pedr
VUmaF+LReCA7Xsw2aXMjjaEZ4pTTuj1jn38Y/hJDmlkyQm5JPlhNKU1WJBED0uvr
vD7+mifFEQy7bxGXgCUoGDTFG++YoQBjbTlHh2n0fYnV06ErZVtUFc7DmvS8nGR+
M9DInNgThvCPVPpCQjAPMldoxYByPII3bSPuatleU1eEvxEV1KS1BKImXnCDG+IO
g1lZfLpOvnu7Mq+FYFGhygOoh8KhhhXT5RRirHl5yIBH9eN8AEteTSNEl0kiHzxt
V1PgrWcNTbDRb6Nf4tho5Jsa1yW+SIREyHdwR4QiSy2N3aA5/IkmOXoZ6b4QInT9
abZBG55TzdqnqpPFMWfqr6aBO810B3FeOG17V0MjBLGyUBZRtMu831quO0YwTC2J
a0eEtoBSLT5KQZnFx9k6KD3GSNE0kIujahXEfKo5d8f3HDoAztqATDOk0Y6MeXdk
GQYzi/M0+lKyDIDc5mKM59LAq1J3jGYNkHdcGKulBwZ7EPycdCsWOzUsRVzc3GtH
WkDvZ7bTwi+tk2f3Q9NyaF68gZwC8x2BzAE/R5rqRXV4y2nE2Ndm90C+xkDTRLep
DWUmpJWsUC8Hqr5zp/8ZoM6XrcivF4BFmXHM9w6bAlilR4ZiP7+WyyPK+C8cfOp1
hr/SdRAenlUlHYdt3Zu/S2a8fwfvnOB2rut9zOZOTDAm4QGA415m9HuoPlIJB/qU
TSwcZNhubL7UYORYRbd+eIsV95hX6OI40FpTP+CORFgDPTuq0S0JJeBBeZEobMq+
8bfJBzP6CMuJanQXgBbssqg1oeWhX+5RflyPzuOAFsDyLXpAGzhi61Mt0noYtM1q
Ik5SI0XCcU1YgE76+hwxCNdm0erdjLrc4egH1zXXvv4bC49Ix7ls0mghx2Wyab/I
ll0rowSn9pADAmj6OH56zxNh0zSZgFWjSEvFXY84F63hUviXOX+lRrOMg949bJYE
0ZTP4n0jNuCOlt6fjCCHQ0ETPjudelfkNTaIaLk79Osf7fHuh1MNucAMWe0B9b10
3HRKBvEy3yfGuqA8a+Y2N5/rcV473O0dc4vLjqBnFHdp8ittKPHbQHp4rzcyjTkf
p3KpqqIWJzI3y18nZLotUrP3pQoYViDVC5qRsPdiX4LWAeIxCrVrnpk2++h3550N
2aTOvA8haYnoA0TyJa9oLcsQkDOTP+RbeFKhLqDmlHFrjbrLe2OvkaCFqOxpoZ7K
zHQBnO3jDue1hqTrY49pBM5F1T3DywP4q+bCst84BAfuS7+CU0+MHCXcKaJCIITZ
k1Aya3PzU2/vOAJxiNbPhZ98UOrGDIajpTzuEvjCJ14YaR3erRwX0UCb4l3MyrqK
TaJy7dvWHuN+HheJ4fN1ingLCKrvSCQGZoUmJw2wZxEGxJ59p+a8pluCyNum9kTm
H00DZSoaVwWee6g7cJrgaIs3xAC1Tns3XYqPCGcXYgsyo2MPFTLp5dtbOSF0/MOZ
TQ+4QXD5uUA43KAveouaWGTYqfV52cu+V9VlPsmB0Tfy23BJOjlEZIfI0jV/k0MW
D6OSROcGSFwqaLiCKS9OGkBNUJ5NxOGieUWy1TEBGjJmOqkLfCxNUXaqlVlCYwJ2
XCqdOl1hY9TmBJa9eTZn1c8KHG4OHFSgsppe29Z4iDl8xFj6A/+Ve/de8f5/4b6K
G/qjWXzEudmSOGFc0H798OQD0MdKioPQFSNPSin+zdOjZhS8r2+I9cUMm1dL8IOK
u26RZ4pGqz5QCflgHTHyVPzG9Jw3c+K7CBlEopcdWLEmN05emWLHMdSNgTjnSMFr
EQUdw0mF53kJqWuElWHQ1xzIpdcGHw0JSPxq67ulax9ppSCKcb5Z0mqUjnW+Otvc
Hg6WM38Bblyc89CZA7ELegU2MygupohWUzeTQfCGGEHweQ3zCHGjTFhOEwmaGPoX
C7jub5itmgAf+udUSDpoukC1CjOHXqIVdsUWOAXV23j0XtBzEu+hF/L10xzkpKDo
9QPBSIoO6KijmUWoUqV8PZxd/1LPtwgpHn+G4nHh1YQhKIm77yVPR2KGSTss0OpY
GZwJq32fNrGBchHt8VWotVOLDB5YkOq2Rb+dc8NBpun07sRsSqpSZw/bi7ZzcYQ2
eQS+fB7ELJRpWXkuQY/V3f5mgsHoGCorep2hoLAUqtFGbYitXCBg3IqokBfAEfCi
CKMzpCUbgvfdx2SbZtBCcLHov3oC4qpuB4SkHFMA3pvVErVf8f7lOBBVPNWJHIwJ
SwqAmcnYXusex4sy3YmyO57S8etieNbOIvC/JEtfPGIO2WnxAqGJ4HXHZ29XksGV
fpsHRPUxLcj7frpHVs63ofH5lq2+F7FyyUICnB4EljB3WVWxbTpPFaHEdpTb2Qwk
3cWxVjuBVFggPxkCKb9b2GtC9dgV2HmZ0cUspORx9QCBe5M+ma57mcir7K0xSWNz
kxItrrtV/7DDHGqT3190TdwC8KzWiEgbUabeKbAO16f0jtwLzCvRZkL0WFOlnRpQ
Esph3NmZalwKhj8DZUCcTTWgxaLULs9CPHcqlr5WT3aeCUrp6NJZqh1h9etM8IoH
Zn38YzKUWXzJ/Nh4KhnUkqn09o8knEk6uGs7gECgR0j4ETW1Lt5KDvcr/yuF+Esg
HmvPkLo+Q1B0NCPfUbTBr7RC2N7n7Sqnps5Jq0syR4y6HDvx3JCe5D47btbDxB+7
HbYYaNAnXHlTuh0J+KlnUtwAYgOZBvqkccb2cXbe19FpZA0YrL2oIXOP199Q7zbI
xWnO4Gs0o2Tb1JgTtDCej5Nnkw6Fv3nqPkGvLNI6YwTyLjY1Hh7nzr6B+yS9WXMM
V0YkQz51dei9WtfwnhmcTuYmBkhFut8zoKTu+DQYh+WU1HEcM2ARWRDzVQDBbHRv
0yBdjB/InxamXkEgBLPFvA04sKODD9WtBJwBCty5wHfWB4Ycjs8l9O+KSltDRVig
/zsk1t8uFFCOPxnjqug81cfBqGYPK/9QtQxV/yIkQbv8/r8k+JIc1GReBU85wF1i
HV38E1BgbqL/PrvyJIDXK9+Jklaok57uCeXBPtwPxFtEMHZieRfVN4nJV42IITqp
9UhocrFXc0kBGi9j1sEX4JMTC4T2GzC6m+nBMhO0lCXM1qnZlaVdu8QL/mHvvwXF
Dhs7P+fWi9Iob2tJRuDPzWuzW2PpVaSFk4ipO0WupWVwfX4vt6KWXq1St4vGm1Hr
CXU3aAaW30GaP4uow/bwjvGUnBxwJgsvh0dy3Z7q4vNHE42m69mhMqfz3FZ+53NR
v8ztxy+tAGmhumY1UX3oW/vvFXS+1EZt6CRKqLMpeS8ZKEfW7SLlVBJEAoDDNeo5
HEGq0iAWpIFj4r/4Vu/TROIxqp3PPYeTxG/X2cUflqdmqdS96R59ybOzBNGGX+nj
SQ1HHFhDegt2UgcDuDACfH9yGmxFojDD2bF4ezd/F3NTA0EG4vQkfl6JUcOOtMhD
a1yxN/QEaxW5CtauhOg+Xo69MgJOFVS/8eXnG4pqqBaxgds4UnX4hsUTF06AY7Zf
wuWTENelRqBQYm08F8BRrTMovTe0lch1dGo0R+tPTdGbK/x27Wm2U35IgGl0P5Tj
lOuHwt10tTHssXR70OTysJlFqI8peB02UYhTwkC7w0uAH36C+0dOVtR5WAftGI5J
w5Ul2xNfe5QIm99k8wmVGt5LOvp/RZ/DaOvZy/qZ47xx8hPcSOvnyAKBpr8mZw0F
eWm2zDtcjl7jZxWG/IaQWW/VYPW0ov3rImu/sN1Is1B6Yq2aQa1dqwHcZmTCF5Dq
qYXYUoUasLCG+fmqbZykqNdg0EDXIRVs8YOqqxZ3PP1w8A9PyID5wtqNFUj6hwyv
5tVnSHHMPRN+dL8p+OheGHpdgsdW89vVq1bjhNufV1qnPEvYE4nC369b54CKHen7
QFSFAbwZKd9+mtByI9q2C9asMjgNeiwizm+I7eTIc4ihgNdkXWkFTFF3H++tFEbX
t/Torq/vqIp6a6FotkSHmK6uqdPk7nvmQADCRbfYxXDYZ3izHS/YFu8bYlgaqWbh
p1Pi5uQneHQQTF7XjD6ubrMVA2jn9hHWAgUh3Gd1M7+dy1FHVfZoPe+qtTs5jqE4
C/6OA/2ep/UCKkVuZOm2+bIRRDNS645PXEcyNLOKfL3xkXar1B//fakD+03Co64H
RdmVr7h/LdVtBK5MG73uWPTjiO4hhB0aoCRrG7D0wN0HGTV6lzAyMpAN4nkUUwKd
52rh4Ej/5X5sGg7PkRhTYw31gHcYn9VkbIrT3kQvrkhkXNWdOaUoahWXuoqYN6Eu
q2yJxuL+ObV9QWcS/qbc2+kWkeg25sPMpjfSu/eDXN8z7jGpBoOfeEG5ySqaaX57
KQ2w7azecdWqO4uzRRBdYM6SWwMtv+NDdEUUVMyEcOK90NKuQB6z1NVRUx2WRnx/
sWTppFZ/huvb9uG/Paw0SRLT9TU1nVVJdgV++0t23aQT4BT6aCBCTkwoGAdm1Prz
2MFRRDqCZHQSyX3J1Ps13+azLzevxauBuZ8rEVWaizBsw0N7Cd+IbodWLOeW9VfH
gMoQoWhIjfcGBTC1utd638yKyuhDnh225QHFfRse7SNCZLxBYzdk3NQ65BVhVEji
MV2bYsdWg1ZGfkNA6t7BgLNuZgHulnyOY2QhTU59okfMaE92dED84urVd4aOXM/v
OzH5FvZAjcUSSDHnQsakajB5/GfyYY8BAR7MOLvyjHjuvbqSfcoK2ZDt/EBHwP8j
lUhSXZR6GQADiTTQ986tlxh4Z01/X+GpxijfGVQszGRHAmQIrhSfb8Y7zDEERJwg
svc9tgdGo72idQqQKN32Cpz/UMoz0305w8r6EY6bJqbZPgfy0nxl2U1Co82Os8tU
SZ1+haMR9t/QOIhpqdjbVO+9Ck2T+0Gu4aK4umGDSBAFj1MP22d0gpApRL8UJ8v7
kei3aksF0aybbP9Xl+JSj9JIlCXcJVktYr0D5ougm38ZeveNEImYrYsjrY69jXEa
UhvCiAwv743onCMIAONyzidxSIpMP0CklBUp0oJK6/z6N2/b4yRhObUuuw/nIBKG
zohLj0S9K9hoakpnCiS77DkRN9GekgpiJiPKTJz/Z4UDHWE4qiKGXIyKD4rq0JiS
/bZQEmHOAEGlmB5QF9UdBkCHqBhWB6g5Bx69cXIUi3sab5CZwSOCGKUsXP83GAkp
Pn8e+ExX2YvYHF6aVrDB+H3yNWBS0fQUpItQ6LwKU/1ocv+85uZvi7tBgbN0TLSF
kdmFlgBnSr9AnvnxBleE5By7jCx8a0z9XyFMGPzDBsHMuAwz+q/7lETVhrdF3ivN
8tnP//3iXxwUfIDJOwPLMxDHaMQkVUr5jpsU67B9IBpUarzq9IZepwwtTXBNsRKm
PF0zGzN4F5msI4mUw8w053GABuEy8SJgihI4xN/GCT83MS4E6lZEb1If/oN75wV9
tlXrsqzAKNC2ZCW/tS+EjUEVxQ2NVbgt0cpG12tUMQcbr2Rif9ExcynNJgSDzhLH
9xtxgxPUg+OuGEe+ZJXrf/4fr9roDmOnfrOlrUMINoM8QkyLlzFG+F9asVFYAOZ/
MQDaeBByFvyS7gAPW0UV50iPKEPax9mfBMay2/UgZ4pOQN4F0sjhcxRtFyOolQ9L
CxcZxA7wZ6TBxRIbazpUPEQfcnC5wsS/kXI3sx5T0SLoL9BRM0TqraCUaoxZx/eQ
gbNCJ7L2ZNq9RLW3k9lqEFZ/x35X6ktEyIBj4Qbc9maBhTCElr1QJ1JICPeKpfCn
XZfWSmoaFArlZZsqVThjOGZuDvdqe29mzXNU212EiV5tyKEw6sOE+Ver3mzSD0wm
JKMpyOWhgnC+x+Xnt1ye426MbClj9jgVNQbLBTEfGEq2GgTpUkOGRqUGc8TVMbMb
FECewO+tbB1S4dwS8y2q/8rdMZlOd4XKnsmRsouZtPvGkhM/UNPBf9gc5S7TN3qI
PDeTrg+5ev+Fsubo6x1mrSAI5/O6sN8Ben7THuv+byIaOa8PPHpaAIgKMXXaKy7n
sXAiw/zW9UgLHenp7ANfujrQgiOTc5KDotxTlwudfGQOuIeNngO3nlTbMPWQw9zK
yGBY9nXCL1wFZBYkpD5OZ0wjhbv5vkR+LJZ2jvNLlfXTTL+a/FFBKy/5ySiKKi8X
nB/2oZQDwSddTgv4Jy9bPFghvs9I2D/x82Fo9eki2t1/7rptDbG1juaIl0rhdi7M
RDkkIRp4q3qsG+Eqj/z1Z9+30SOVgLlIPcIKgp7os76mahGafAjPKqMP5Mxgv4bj
Vdjjj68etYLGWHd+50k9N1KOvnPuKAGlQU69FwpzmVOW1ngBkF9WkBaM6Wmg5k0x
YV15BGZCJk5vd96AyP4JsR/wMMvtDagMYudGll+if4OKZDQ7BnYBlXz2T6RnWitW
GZ5r6eX+HYX4zNH8Fw0UO8HiIYbTpz1747Ej9Cwpsaml2zfj8ZE+4l46/mCXYP9k
wsUDPBwlh5US0FpRwpYcL0rz65P2UR+8OaOILdq9wWwe9Q2TEYHMGjgEy7cjreR3
uBaa0uNqt69lnI+XABwJdZsPfV1SM6hAQiJPuvpiJbMZ0J3m9+ZgNZBxvJD9Wq2Y
OmlOqMUAbkP97jcKO22807pe0ppNJQtMuIaRnndN0cfpNg68AzdQulfcdmfKA8g1
MWo7uLAGAKNm7O6I81X9gFuzHevy6JFwDSbqStdcsgWjdX7gTtTJ5FjC/u0tZJ/Y
Goo05XdxVBfS2U1rJq1IeviwPz26hrrOfeix8M3wCFJNVYUpTRsv0jkKeufFS9Sy
xUk1CrvvXjbCk9opqwhHHn5wx5v9PiN1I6/Ote27ewU441EGOz29TVVpt/etYtaO
nA1FadvE03WfibvUfeneJWP2iy3xxBgVbqIwrOEWmmLjreyDYQrQaLOuBeBOuq2Y
WJtznCBxw6L98Yks7IQoU90S0qbI/ML6zVu847VyyDnTL1r0Aw4khvgUbdUqHr2Z
0VMTyNc2ovhFiO6KbNTFM6WnxbupjmxeHOy4zjS28u/hlvLrjSqihn+6AwmYSkin
zgHVPEekXETfWuIlDQnE+6SoYYf2sjv9QdvLu+9uzjKveNtu+KiXsF5WKmR6Rwr3
uLh6k5JhkCOjpthkVC4gPahWpvRfZqdXH5bhr8a21gvAxaMdrQb553uVMwWQBuxO
IKfZ8DjC9hG8NlXiY8nj9MicauZzpxnya5gWfsyDzk5jXQYTR/dOQYO0XtP3Hg+m
IelfA56W2wXsr2VOtJRmY/NcY33GcswIDjWRa717tKM2xVvyhupNUI0WmrCVYiox
ztHAZKsJDPccEC1O8n3QVW0J3M0buW5LxgogXb8ibQK9c3GJMiedjS7zL7qgS/QN
pHxVUNjDYfb9petxfg7UwlqeDGOo9/0WZDCAAdQvx8Y20qOFNi2lDe5CvLIovlEL
x0sC/PA1LTc/RHGLnvDSpJHxuDTxF7yWQOzvQ3EloLVlS5u/c1M/P8kqE8XyaA7u
ktEBmKdGOL73rL1fimiRwnHIuCaXUda+K9HKMb5EUDuTTUYUwmS4SgZqFd2l5SQ8
evFR0Idmk22f9hHymyI0XGGSMCMe5JmsfxyS8MEHr0Kx/guBUEvzuOWPHw+Hi1lQ
ea0Sqxlk3NMUG53j2v076xeuNJxdk6jFHIpvRw4McAwWe5Qpoi/tSiYwK+sxpP29
1XlbMigLs7FSuAPkg/SVWPTcN/MqlQuBw08DWzHBd2AQVIOsF7Z+/FrVCBz7xDxs
kQKkjezH+OYXUc6cD9tkzznjzajqAQm/78AIyL6anc50XU7BQTGcSvW23wsP3tQ8
UWAeSc8RulXZAIStP6HCIyyA4ppuo6MuMu8QnEmlP7EmaRmUyQdTjLl7bbsPPO2L
Jm5IAK08fNclmQCvdvB06K8P6IRmEqvlA9dMTijAAsLhe5AcVUwytxNKT3A4WqCQ
XK3flwILj5nuyfdKM7DwzGnVJKNy4Sl8R2WTqkPu9LD1hNfxfj1u0/vAMccGlDyL
vw4UaDpwhJZFYLPIHzbNpWW1zESrpSUFp0Pf3h8ZCGPyAs2ZRQ7Bm6OUKsR8+OO4
sf6a38htLNkATlT6nyLKw+F0M6hCF6mz/0FGSxVizeDYcnyI6ZzZ0nB8e3mqy1JJ
mmqqbkm4q0DYsfrQ4/7aPQ==
`pragma protect end_protected
