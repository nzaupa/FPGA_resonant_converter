-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
j7kqdqJcBLn11Zyn9ETKFQOmSnMmLZd5McaK/jyttSwSAw1OOmIsMBT1Mx1MpX6rIoLVD/roVXXs
ii4ZXSpSwTADm9sIDFA7GcTyB+uY8/TPcaeCzqGQWyU/jrgTeUbycTBZl11GoPkCQWOz8Yu8PwFb
ZFTjq4/64nH+qEzU1Orw5QiwHDQtPurxmZcsFTSGyM/mvrVYCObCxsO1tUoU7u/+D1zhmPs9ojaI
uyMEhWA5mvFqr/Br6g/Dul7EwIUbfdc9+o8Gfrf4zHmpQzmbl+M54yL5VQ02ODvwTt99XtTEn8Xp
CR4/uzIDSoyvIfTtIBXH0WLz2pREp5CvcsRpwg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6672)
`protect data_block
Tz8wzg8EoSaRI/b3+C3r8pjtnTc+k5RrZD+KyFLBy5V8ig6JG1T0qnRlLsyAdkAxokv4MMEwl/FE
6c57YSO9gUSGDl7loFRj6qgC8XhN+1mFvp5mEcn7BtvaONfepns23v/AQ/URhjCvHUjNpz8RsDrF
q0x6YXsFi9bj8a+M1/kd69ZEY7EPjGVntrOJvhQ3zfwVd3IsKq6y4wutNedVLuRxeegLGy9ujaTR
15DCwGVy/DNg2GAtaYX9LM0jlnk3B1QnRYJoM/btfUb1OqhiuqxvcjlFWprT5wR+ibhDHYZWIPPa
4Mi2WBRbYwN4BUCPz5Noua5Xc8MbOwSQBxydsw8ACmPWUYn6v/KqlsETSLD9zcTglvQHZlCkKW1A
NWfYE3Sfkmp3T4Uy+b0f47TsNHPBEdwnZyM0iEEkxW2aYn4CAEs33X4St93svJODZxB+U0dUQ/tG
biAuffFvwV/RTigfM2PIbTWcNMGANZTcx175EFPx6P7y18VYc9QjB1L2M4z2vIxE0IjV/a+hgQTq
BiNSr7M6Y6SBEzE3N9b+4DYmc2HQwfM3FZJRdHLhsxFNUpiPYhEoh77uSOkKsfm1DFgRAKETgh5R
KkckP5kNH9dWOHZWayMyyvLaftyqBGXN+bpBDTH1z4hYee0CQVrv6BNta7FHB8NCFTijqpX2iahS
1pBmPuP4pTVbkBOs8AU0eGvwPlq9bJTsjoEg7VesGJqS8E63GYHJRqDx3/tkIaAHjGiLXnNh9l/p
+O5P4RDnVKL7NT1MnH/D1sySqQRL8h7L6iWWwSPG64d57VGX9ydQgvrRZLW5OGKNkplmIW6+OZ01
qdSiocc9hDSPml2pOIr026LFowKqo3PnSH9EIKTqfGuHEvqBl2Wm8wFG2+XuoVu1MTFtlBdKNowH
jlhtsqVTHnVpQo0jZO5eQVpex9jKweM6vDU5fBTbDkfKrC6cWy9YuiOY59i0OFpHekShFmQ1/22Y
5VewHp5caTLkwx+6bBIpqewmS2injQc5HpC23iXCNcw4D4EGFx4OsdcVmGdczRI5FHErJX0yaWGn
SKKhFMW+iaADWIGs4JafThu9UGx5/sENTsEQoK2UumFoEu4ya2VtdgYqpqKEl2LcG3gqEjF9eqUm
26jDDrYiji8BxLjktGxLNa0meoYbiFlWtLAL9bQwlt/vH8prXUYuAoALjk+OIiS9YF/tFx/RWDbD
50OXMFLg/UF220dPBYBOQu8E/K69A+RUjzvp0/IGWSsWkzxerMOxtEXZivc7mK+0asheUH7lANDu
ZCDxVyLm7kAdYuUPNEH7dCINiim/mDlx8W9No+KzyMeVYj1OWgwAT6EDuXjCjv6rrZnOQeCUugJ0
oDXzK17OKwI7pnZbtNZhcm2HcjSJ0fKeg5a3LWjki3ApwxftJ7pkcCvDIr84TZZxL+1m7qaVjH4F
g6S9f0GjrkLAY1LKvPiuhn7TSMRv1YstVhflvWyWGLpcCGZku/GbtLWQkOQxE4VZLmfN+YiQGq8n
o/m4s551w6RcxqV2s+4G4+A+MPWlbYVBfX1GYKYCyUrW9Om0p7Px8hbIGNG/DA+YxwCv0t1RH9+U
p/DHLTQ0X5XNPnx0TqaB8EBAJnDOwjW2J7SHgJyOBZL7peyheF+f+Z/Hh4yX9aj5psZYX/SuGASw
1rryPzzMj9VfZJZL9/UaVJB7VuwAE24tnqHoBkmwt0T2/XAIFMKyzcfjrNrzimRCI8izMfcEpYD/
MszToMo9fa1CyGn86cauNQ1+r0J5IwX4IPS3R/6jzGcgxgMKzcYq2wc3ZeIPlfJg1BaCi2Qwo4k8
oUaNbOfRvN8bfe5GSzK8sz3mW+xuHWvl0yZWYFLnkdD2UmTh4x34vvamJykhsaolF8sPa3u1yvoJ
PRmjyAYupfzcBoXZeo+kAoZn0JULhUrmnymS9uRy7ilCnTatCGbNBoYteRuGyXSOr05Jzj9Mgf+K
AsozBJUvu98f1fjVoxpBpq7O4MMTR8B18zlZkr/mO/ht9oyLvOqbL+94yuZ6YLkiosSF8sPecZpD
JQOvlFnJShUhjtaLmqKxDuGvZFDyLebFV8wO7BgnC5bZhKgEM6FXYBQnvUmxoNa1kyISe8IsXCg0
TQ1rgMq9Pn6B46Ir2H8NDC6hwO0PyhIjvfg3nUgm9qJcL7TVm8dWunbH7o059IcJZ2slqPYE3+bw
mF/EADbri80KLEvqXaPA6p0X2R7LAPVdtfvhizdc39gCeNcu2JZdV5busP5Ln2fpvreT0lvy5HH5
bTi0C5VyWqIuBYY8UWOeMDnmalz9LdiHKuP5aNwLp2VXvhjWbk9o2wuGiix4bxA/rdkqjzUyPyHq
VPsE5rhmS/9DJx8jIot2rlqDBZer3U12KM+JKHwad7fqQAj2PbyUFiFEkBJHBLpf8J9TJBTTbG7Q
pF9qNLVdQFowo+KfNhBbgbF1G697f8q1uICBLcNWaa2dH6RnyCVS+OrRAGrLZDA1/Loo91cxoUii
6gp7KxEjNSb9UJRNBoc/Vnu5mMshjxL7kSlEcxxRemSLi4iM/W8Blq14nWLvkKKt4Ul10zS5wB26
+vEapEHFG6yZyKKIjthY72LARtLPTMHsEaYfrwgWJSzNIsp+Xb9IbL0PLa7MGFHeCV5EZjqOd7iO
lQigRszRSqyeIMaru8a97KXCKtU6dFJnDGXZ+ySykQvm6Ozlte7PXET5zKUvbkOTvvWOFNR1qcvD
Wt9mvXILzZwEi1cpQplSEmkItgUUsYgVwFd2X5ie4Gq1xCAPMuUx6bRh7DN3E+MDFxZ8dZggGwKR
EYb4J+jljVAlWUBvravcCewmg571sLthT+6/mvrDhesACPOpUKOd6WtIebcgFX8HXTvWrmJGi8N/
CiEKz1tpSV9HJVjXA2gDU+Yow66g/xysr+hTJgbCXs8d0jMbrJD/6IXZIA87zhaH9+YMIENvjxK1
Lt0lH2vWUlzcZ02goDQgykdWmp6YuavdQh6T+JC92Z84gyLLUqzbfDxu1anD0SLgdVRFlsjXrpfd
gJ+ibavG7v2ViGEvqTCj252ZxIFXSratxzDKyIC6mOu+tJnG17do5e9DzWFcgNPjIcrUIxBqGvIP
iRKeeQwX7LcITx9usg+vZ7RCQz51SteNhVmktU5YlqhShy28PnlqWRGhiAimnmP6GcCoCo9GbEKS
wFMww7V88e3vZ7GexKIk8U1t/mIgFszLUE+DR+0iTLgD5Z3x8JENyPsQ+j9CYmd/zqSPSHT1N8CT
gE3iwb8BurXlRMOGZyinhGePUSPtDJm4965sQrSSL1FoaHAzqvLz3eP66x/kOTgiD3ftbxwiz3nP
LSakm80QdPQ4DIIErML8brRPvdA2vY0IS7H6r+7FHItRQVa+7J0rALmGKDAiInqw6hIi8CmMRKbS
UexEkg0Ihy20GCOCao4WNdXtVojAyUcLe2z0I6E+bPtEkhUelfFAg4wg8c4F6dMFK5CnJtl9+59R
J8+BtZ4zLwyfqqUdMz+xSE+FiXbRFoNEvZMgjmJmirTD0iyTEaBsxX9k/gEzcAuMiyIBs8FoebS8
qjXLtR5F5c2wbJMbqqe37ab/6OknhL7pCvVXld9pkYwC1Ce0qeHGTVXj29l9tNsr+YjLOjGo3H4R
lgc+Grq3AxhBTfs/BLtl0W0h/3hnwKAdzwkDG7rimhPg08qUxFndTLT7ywJ8resYUa6Fun7r3Mkp
I2bTtxIXETROLGt9GYosib6Tw3ygD3WWZ/BjE23NeDtT2SxEfh73mDf9JcAJewNAG2lTsFfuR9BV
YsMRU97Ke8CDuHR9nLCk3piDgdoVUHJndcu3d5u/oonjS31RfYdq3ZNc5qt2yPUw23tIP/8dQDx7
GWO2OiqD7hH+tcn6TdQUVEPNjv/Ltr1bUPgnBeyL87e/cYXJp4i8oPBiJvIiqnesIHTCebYfybGQ
D4CTAAsF4d0Sh/hJDl9nJPD6x9sV3o7+Dkf6usrzk7p5TEedYv8PYvLsVNxn0Vvq/BWwWqBDJOWd
7YvW+TDmpsmpnWx/mL8zpd/OKIIUn44H5wVZcMcEo0Q6MbxGSEYn2UNVvbuRz4jkllM4I9RPL4wa
0DZxVdhcJI48o+9X9CHJ5uSNmFNwwlrm0/DEtOHjCCBQCtkmDIp17o6XZ07uDSBlCVXGANm2tItK
ebY4lU0dRga7UKKziZLF2XcywEOxeseS5I9iB7SX8Ktf2dEPnJV4zcsT3R82KWOjaBAD9s+Xs2HE
IK+ErN1pqrviV6F/v8ESKuL7tsOT74zFdjgIe3x9JLJHrfYH5iDlqePb6QUFt+e1p+1nxXICyg2v
vJlLCNpn+KXcsXO48VJQ6ctQkMJ1Z05Rn8GMd/GC2wq95s+fW6Ca/c4eHFm9mVp3foG8ZUgflsf8
PTbROpwKMhv62HaWRTm9bnsTPmYcrEVU9Ggl3vNsHHExzhlVWUHX2oymy2xL4BKd0if5JrPpCiOQ
cB6y17MPfvs0eNKjZnaI1wrLuGuLfVdJuyPBU28XIVh49uvIeux5vtR6kDlslZC/mYsmG1pwfGvk
5b20aGWnTSwFjTvkPBHyUUesi5G9Eibt19NqtLGfp8TerZETyIe0eKTa6edjxgu+rhQEXqUgOdqB
po2qdzvj2d07y+N2eZ/JTdcewezFkCbA6A2LWsEvsl5tYPULL+FHODpgINTQSZ/O91vHIKYL0f4K
z437mh30871HcfgrZgwJOFebCBCi/USr886u01IELaau2jVJ374Pdn7L49ohKM0u5fzUjy1nZJ4b
wz38EaVFFJGGXB13KMmdTMShs0FKeCc4bOzGKOkhoED5bandVVOC3vueLXqZWx6rPmGW+rn0sKuF
HyZQSSQQzbdmP7HJ5K9CI7D/6GTXWxKpHZj9z8UBBp9WBBLh5yZCPTVzF38PSkvzZ3H9gP57QicO
Ly2TEz8QdYePneiHLoiXaWN0QTfOH0VUhEyUvbZzOwuOpWhjhS1iHlc0Lxd1ZLN1ShvhpPSaWgCV
dw30nOWPPXj16CCrzkf1SnA8pGxUFSvIS7wFS2cY8pzG0rDqsri+yurCtUz9hb8DxUIevDqJBE6L
3FeevmWgSqx2q/vRrdWawJIB0i7FfhbQ2JQeajk1UtmxurCvN76rO5AXx31FJvU+CZvAckOmrlvB
2lGrG4vnGkAdUGknEhFhEpLCjugk31g0Yhi02guWhpJyugW4BuvC1EN6cEU8qIXvQUPlhvbTaNPA
aL5TQXFzZ7xn4e6bt2uyrKu1n20/iInzqVOpzXZKuS3aDT1omfQxd8os7kIcsOHWP9Ugd0zPixqy
IDYJUzDhiv46kfuKSHKGOVzYmvynDsBpZxzvT1XCBpTMbS553KJvxeX0NLtvcIkm9c8yA9hJBPHa
34cAnNj+d/oU5KJyFkwpzcpSNAkUsKcQbb/KRhcclyQb8+7JyjdOYWhev/zuTzZpJnfYaNwTBm1s
BFRtYeSFk/pwQbP8F+DcfARg1OTttp7TopkLA/4YPbHnR28ofjEpr3HiKaWoL84K0oMOQ/VeWQBt
H4vWjZa7DKVULdevBbU0yGC/HMnKyqKR6F0q5bZEDOPpN/anBdilfwmaZB9YKx3vhHOrYgx89+hv
Q/LiIM5VKEb3z8kiSMriobF2Re/i36KPIcQB3ZhoxHV4TMgr8RvWd3DTIDFkgY9CuIIosfLKVJ4x
xk25tM7Zq7tzkPY+bo4CPX1aKe/ixnXUFZ4Nx0a98+4IC3FG/iiKbKMd/QcsW6gbOuxQxG4EpRVf
LSAmLpumRXPB+w2uTOnqIL7THlFa0hwmLGVTxtKV4+/oqUkcMAXlrEyckTnWcI7A8qi+veROflva
qDm9XHhe5DYehVfIlfPCa2JeDjd+p4Zi578NRFMbMPyZPCkfjsHyRlhSEJRd9YGCf6nMiJPzZOkg
BbpFXDk+ApgTeFONnZger7avOgjnd0sBwrl1irx9pHX+LkEEsYeGZY5M2up57ds1xMNoj5dMMWSJ
Gtw5ANV29ZWguy9kr4ZfaD/b8DnVrIOYitmRefxKRy+Q1zoGPj6aK8C9sAL46336mlHVS8a0D93g
cSUXV4KzVcpfUS3dElOmQk/Bj7iyQ0vyXWBKVo7XapeOUmtNMt28r9/OW69dNhSMgz2BpV85qZSi
wk0KnU+82tmIrwicHdoUROiuc0QLjFjJNI/6JbF1qUba7B5IfaruK03AN101l287Jtm+2yvFUGSx
byTDgSsFCeDeutblLUcrFRy4YfQesmkf5B9hCDYQit/KuX96IbaG/bwf6iRjt3T0dG01yFn/Jrke
E8OsrZb8DWlZXilEJi+GedsjSz9D1VuT8sOTtcHoe9vT5xkZVNN/hBysUDhlaXbSvMxzvZRR8inE
j6ZvhlW+s6mFAEdy+XKJvrqJUQUpt0LVKjccR8MWdmoO7BPBGMM3SEAlXddti4ZFsVYNZGcqzGL+
53LpaW7Q+0iXglFGJeteOAxfkj0FICTqYTPlPKA4qxYZ9j/nUs/Szzzch3mBLbc/0TVNr6cKT+c/
sSMf4olcSU21ouylE5vkzQb/GBcx29f7Jw7Qqi8GO8dUyGkW32h4iqL2wtJFGaEZGRV0qAZ7H3bp
3Pr3oe7oSSlz7eu45wZiiDeA30owHETJH7deDfmdj1BIfHE2r8QUekhyCPFBsDFufTvcpI+rssvW
og8/q8MYTpeqRvfH27vzShx93vn9ipmEjkg8OZsqnMi8uFwXoZdKLmAQ1r5I6+xU3F9h+YDZJnTz
tA2hp50pXKZF/C4UBu7lEoEr2WP6Kd8WdeCWk/06f96/ap+TkLcLnscXl6rL4KriKNr11am5CeVK
6Caa+X6ii1R7Bw8tVjNqa20YzUi4i+Dhu0MmCzfKRvuNy1D3YNmDg/uO5oAw0i8GjpK3VxFaa2FH
CCMr80S/IL3BfWIOYv6RIGBgRLCMocKG8WDDPVanvF2+3UXEyCiuMOOAuLVTNiF7v6KLoU8YyIEh
R//oLzxb9RfP5m0G3FZYbAKGRVsPE7diXO1C7FkZ+dSKE4n5NfDKp0Nryy5kI5eJNqsXFn+B0KKR
ibQ4t/XiIW40e30tuOWiJHamkg3vBgdyZ9zeLiA2FSvCCXLsliHSXRJiAiKqBD32odI2QK/wg7Qm
PboyA33X3B4WfhFcncAZtKHQDg1y30TxFM4YiTz8GMy+RcEYVGtzq4ccKtmVYhpTr1vgIzNAfmuE
qsocjQK2goHzsrPrw4u1hSDTqAgQ7ETyKLD9P91IRPqBXHD9hTmsviKwUCMscxOfY24+daZUX6nj
LR5dMwpWJrrrnW8Job+fokto0uxjI7Elir/dyji5VjuGcu7AlBbUATa46LbWKblJCyzea+DkL4G+
f9MNJEPfUSgBxVSJb34fgeU4pU9bM/ytEQXx7YFtloBzd1Qui/mpt6tXtIwQz0cQq4bBw7NsXvEM
pbEIppKQEhn0sYWpoYU6jhNeP7V0I8Go1MPHue8VHoLoOouv4WbJCvQnihCLP90Nt7LfKddP3iaB
HX/sItqcj3ODwpqvhHftPYXlyCXCXQL5kGL0sjCiXk1I048E78AovOFtWhssyDDC2cYHS8HFkyDF
NOti6xAdptimV25uNy722skH61M05Uk4gr5PqtaPo5L4fT9rpAz4mqjE2I85i/HBMtZ59+PkQTy4
GWVr6QER4IcftAhFU5gpJGDX4U0BsyGPm5n9sf0WfRV1weztsBg4rno8yD+klw2TsLc2CwmRC3Ii
Avlm0TSrtTaSjHY+ncZVYY+5yKn3wWF9Qx9xAnfDxeXagQI+9zgVeMzw4/P6NlE9bywhaiGtCWOA
iw/pLXBLuwLQZ2HfeqAW36Bt90KXjxjBKPLwqb7kYxbTNvI0s9KeXy+jSkAkHIMT1obvx2Y8lcAa
eeubYOQmboWTmdLukhEZqvCryar/dnKSTPx+Q404V980RSnzobDe7xgAbcaMVgg/GO3N06guv0zj
MiOl8/mVUgWJMcD4q7bZPPn0U+vq4RTyR4K5rFKfJ5O7dWarj4T447n4ySIDPZtjz79Tmh14SsjR
0J7kw3m/286AxY0aMmHTx/0YQyGgbMEg9TqybzFreGlbIy3eYlL2gZfZ7k3kKCaQOYgtbkaYkJUq
7T6zuC2AkgHcsHxnw4IEHLvR1e0qBdCGhi7oDgRrteDMRL+pnchEa+VOm94DN7G963aisHJi4Aar
Zd3RtRQoZFgBTDjwTguQh5tU7mN6V3+v6AHbZ35ujVphxlTlYr1xueu+vNttHW4owbfUKfoT1NkD
ot6z/jjoFPr0h10pbK7hkd1kGr3wthkmURVN5S52EblmORwdeELMMDqBT5G3y7JEF6BOdvq3B5QD
H1I+VrIGxOqBZd0KKK2zrcK4ghmRBR36zSsFDnAd2D2wOpQtcZgnv6bq5n6mlQQKPHwkC/4TbEyJ
Q1qWD0mDP6/K+dqtsx5Zy6rXl7ILY7eZ+GWN7fDQme7O5rwSBKXoOPtpkGJjlD+61uPES/tk6KJe
Lz5Jw+jPU20dLeLtlnMWXnh8x1Vnw/urgkMahFvM6Tgxj6GheRjF9HTCaMtceAjSYyfAX1gT2VS9
ozu+zRQNKl153n1j8tqwohUcoc43H1Jkp8AtkGF+L9ZumYwyglYx6o/5To4QpDfK/N7W5JHOv8Bs
QjHyC/YzQMvpNY5TYjXPj63aBuekrh35NK+dk5+IWdCWYJ+AODnCMgOkNpeAc5hkdYtuizgBL64t
bWgha8Ao6At4HHWeNmxuW9lkmlHmnRAI+W9srnBxyq2NAvXs7FxwqQVz6eivD2OZTylMOsMOhbGC
a+A2T1jnkYMyMTvtjZwBSKu23huSZ93VUPm48h+lGUyES/cuyELZ2a27Cv0WAwJ/o0NrYU2oTKuq
t3T0
`protect end_protected
