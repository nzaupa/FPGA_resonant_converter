��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_ܤ�y��C��RǑ9Lf�%�%X�/��W�&r�YG�u{j�x�O]*t�QH�:JNa9��ˍ*|�5
-Vj*��h��Q�8�n��׍��h�Y���R58�/�$i���Xs+'�Tw�����^Mt�^� �n1dk�>��A8��[���_���$j�ʎ���0��g+��Ԕ����G8m4�B~� -I�/��)�
�D�	�[��V�#Ա[�.�^]�:�.�v˼���"j�,�w�́�#å�t��~�5�g������7���� I��b���SBw��t�D�& ��V,�\q;�Q��C.��������".���r��`�=����,�ڃ����sx�~�'��\�5#���>5�Ѐ��#���u��~PP�#X9�Y�l��K I���3;a�����?���mo��Y�R}Ʀ�j"3�}�=蓖�D�-�`���_J6��B��1�ʯ���8�K`�{��}D��)��/&�^�����,�C�s#:]��D��M��hg6�֧��a�$�p'�M��L�`�4���f���1z�*���ZO���;�t%��s��5�Ǝ����kF��&{����/�z���b��^P �K�I���ˡ�؟LC��N��E�3���w�A�_ӽ��Y�jm�)nD̘��x���_�r�a�{,������#�ş��YE(�f
���X�������S��%�AlY�mY�+7�_x��uީ֜�ۑ�2���]��SzH�ٵ/��m9 I�\�:\�nX�B�	��$�˷)���3ԯT�3��'��9�e�!A]JO�p���\��~QOl�{}�m �_s��3���c����,�2����(�N�8�F��n�m<z3�"�h��_J�#�KW(��C,K	+ž�����@Tndad�>f JL����&�e�=�2`��=��4�����`0�&�M�)z���x�+o��a��_�IL�!*�F �NH�|��lEi}�)�x�K˽)VI�+�ʄ3��}{��I��/ k��"�o�'����\MV
"MY�Hx!���[%�g,O��|��V4��k�W���8 H���{? �3�A������_�G_���n�[١}hp9x ���N#Y��ޱ;��Ǉ�uj@l�<��@}����^[�P3]��[3�F���Z�;?)�΁gI�_���ġy�4N�E]W�>�����ך߶3I֍=Q�����k��W�ͲRX�hD�5�7$�m	B�'=T+c�Lf��bBW_率֩�����u��}��*Y-���&J���J�Z���?�љ�ߋ ����y'�ϯ��2�{�3�	8cp���Q%�h �;St*�3ӤN=��z�U�����mx>�E��	��=t5r놹Q�[f�&ҥ>0���D�=�~aVU�V���ŔE 'ܿ����,}��{��(�~@�"�G�hŃNU�<U�l��Ʌt�hiey�I�ֹL�{����D���Eڢt�Ň���G��%y�3��U?�m�A���n����Cu1�}B�/�h�2|��XlA3�L�"�����͞�D��#��Kr�h��
�Y��Qs*{��^x�<�9 �R��60�p7�����}O�OP���4�$���6��?�@���k��z�jRI�e*�5S9���>o�;0sF��`�IA"����|�/M	�+��?!G�'�V�:=;!��sOxկ0&���Њ����Ik��S�8��@��HR��7�Y� �\��L��
��d����$��-?�l���N���3�M#`���M6��N��Is����Z�0^~
q�%��&���ҪF��,�:�Y��/W���ţƴ�Q1砨���h�= ��\@o��|�J��.��]�܃t�� �A�l�齫�q�\�PW��f�rA,��|���x"GFj^vN���v�{h��|�*���R�E�W��s�JYs?2�MУ�~ў��?T:-:r,q\,s�L-��@4�9���(SS:������ea	 ������0�äC0Fcۛas��<����a����6�5b
��� �<:/��ݥ�q �^��	��Jy ��#�d��릻H4�h:��
�����.��(td��#d.�W�0�W<�y�(��]��4H��DV�EJ;�!�·��$&�X��M��z�vFM��8��=Z����6?:��?]ߑ?�2�?��piT�
.Q8��fk�S�B,O�%��J�k�J���P�o�*p_B�Ȇg~K ��I���wD��Etִ�_�MX��۩۪G*��|\W�Zir"�5�n=r7c��0��E�Xܽq��$�ْ�a�D�x��J��� �B�m�`~ߧ�+'��'�?��ߚ�{05@	�1��uxtF��+�iݘ�S��/���RB��� ���S� ���.}?��\ϰ3א���!m�:Y�`��`����pf�Y���Ƕv2ǰ=~�4�K��x׎L���A���uy�gS.�&O!���5�V�%�Y7��[q�QO��a�c����'3y���Z���]e���[���V.��~2JL�<tVIePȝe�}�Y��ޓB6���-�C,�5b�4���83k�}��#�@�[pp��5�bj�	n��N��[i�*��f�Я��s�G�u�Y���fiր�d�U=�.$vIp^��|��yQ���3L��*N>�n�����K�n˷����]s�˂X�̲؃f΄id�+��;�~�K�ط��)P_���*��{�s�SnF.�OFK�-�Ȋ���:6N�������ٴ��[;ʀG���pŠ���#~{5�����-�1#JǐF��]ө�ʩ��A�H�q�-2/wgQV�"�2@<�:����,�8����\�DM.p�x=� ��1���hc�N���
ف#�ʆM����ri$B^��0���
!���I�M�3�ϓ-U�%-?��I@��P����G��p*s<�p�*��hu���Y��׌7���b�%�c�{շ��H�����㠫��x�kچA������}�a���`U�)mt讋O���V��O�J	��>�?|���}������wƨ��i-����KwI.i���ۚGh;�yv	�Pâ����)Ѫl�p}���/�>�|��ת�{��f���T��X����ܚK�� O>'W�'.�Yx�/P>�q�n{��P��wA��������t��t���[��BQ�Q�&���_D�Q�֤�`D�6��ej4Ō�l�5�ox�$Z�z4ذ?X\�֐���Z�Sǝ�8�C0��
�6\����h���x�k�˅��C2c`#���_��P��Fj��҈�5�_�
�a܀���N���d��cJ�0���Wn�WBg�8U̧u�5-Ղ��C@vk�{��̂h��F
��Sf�؟�$�S�����r�:Z�0|p6�� Un���;'��d}�˝F���jE�C���F�J�Q7	*�(����c �`� n#�7����O�ٽ�8�A�_m��3n�(L���V�{I:ô���9f�*s���o�kI��Qe�����JT��qdC����vj�OV���,�11c�]�DL��r��6�ru�DH�OM�Vi󊀦�s�q�j�ɟ�g��՝�xm=1���I�w�187I����w0�KKKɤ _{?���Jm���h��+&uك]�T����Ga5�z�p�`}����	g"2�d*��q�S���̅�t!�*�*�-�w�]��[�@��^�`�<�ru�@��(�o�eU%2>j�� �����>9�rp?�\D0�y�wvL�"�{��%Va25�Fˁ��S�� �� J׊�I�$
��6W�#َ(䡱����xA�i��y����9����R�NSykz���<��u�{�v��CE6Ѫ�4�*�&TO�GY��|a�}Ve��
$`�}��m�V��	�A-��}��:�J"�?5�;�ě|�����)��s�ת^~�ңo�
J���7w�3�B���t���ZC�a�l=.��k.C�2`��z���d����Ɉ��QaQ$�UAҟ�j	kx�x�UҤ��xO_(s�u}J.��o8�-%½��Z�R�q,0h���&������9@�@��ܓ����8r���I:I���.��	��K6:R�\[��{H2�����P�B�x�H���oX��p��@�o��w����(�$�<��>1�%�a�Px$��K�$yP�.��XbO�1�d7���߁��Uw���'@GF.�s�0�Z�=p#��}�Cí��i[,�J���#����Ig�`
-o�9��韼����-Y�zj ���خ��h�Q��4>��)mԵ@���B~�&�\����n*�Qh��#�@�,I��`���/�[%�3��/=p6��g������eM��Ax�))Nx7?�X�\��z6��D"Eu��9V��Қu�?��7�t'l�d���{�i�4�Gt����sC��.����,bNt#�	�şE>@Z����J�N-�1�=^&�LCB�P%oɘT��21���/G�^|'���qMז�g�gT�ΐS�3��;_�a	DH	Ķx��ͅ�N;:<�^���m~5+{���3�nw���.wqд �]���N����cl,�܉� q�Ε>�ɶ������}��b?�zv���˓923^J���+	����^�?���N�'`�Wk%ޥ�����Ϡߐ���0�0+�GA���C�LD����av�ݞyH,�I$U���a�Gv$�������v�V��C����h�ò3@��˺�vR�pȽ�������i����y �=�|�Ge�2p�I�d�\
����h�K�òrݣ��T�L�I�"�;j�{�4�9���6E9dm�|�֐��M  `D��X?U����>��h~ �3|���D�q{���E�����N��@�٦�_���B��rY��A�/w�8[ u�KW������L�>�w���g�6X)�{�#��Vi�x�ru�z��_�q����4L
(f�Е��k��Ժ���*�G�/;�*�.��O��'>�{��_U6�u�ibkD_.o�}FH�p(.  ��\.V����fM�n�A�Ɩ��j4��W6�9� �=���(����k5���p˥� �,�,nGR��,�xx"�[Wk���U�"�T]kZ�ݽ�9%���aQ3�x���^�
{�WZM1 �k�zb��LT��	]T�� �֬�$�����i� PnMC�G-y��㾼�*�߲�՚R���l
��ax�
�[2��S`��A.[�֕����Iz*�D��; �2ʕx7���
f;���2�㔡��$/;���0���R4x��n�20����SVx�ύ\��Q�����hq;k�������x`ϝ����O"ĕ�8v�^P�M�]+�7�&�-t�5��-��Mk�İ�5��P?�H1���?�������_IG<�)ωOeX��Pª���*�����i�����3<,�/�q��Rޕ����4O�
�)2M�u��jF��j��=I�t������~>�ܚ�>�<�>Į����Y�û����&/e�:4�b �4��ނ+!%��K?�k��%w�3�'E��j�S=y@�bu�n�;��p;�Z|��h��!������:�$��>RW��0�F���D���Ll���x>�
%�]Z����7J�&ݱ5}��#���JAx ހ�-ф=N7��D�s���]�Fu6s�U��.������DR�TY�DixD���c2����ؾ8����8�C���UM�@B ��I�����K�)gA����0@x&���yI��ߩA~�VS��5* ��EX�	�'���}hmܣ@���M��%�=�T�f��úݘ[Du�G1�K��1�@	�����3?Ա����(*��Yy4�]#���Yl��5��<i��a�2��<0 ;i��[)�E_)8Q�b���Z���an���H�Fc(�eb�*��E1�QN֡�9���]Q�Q\p;�] tr�|�B�&�\�����	�a�4a��FSϫ��}�]�1���@�s�u�iƭ�`�����X���Y���[�u�gn�Z�G��x1�����@�5%��ct,��a��6���)XaO3T.�T�WoI}R�w^J|A1�������+m|�W�r̡x#�煱��
����u ���+�"��
��K����]��.��kѬ)A�"{[���Tt948���.���*�{$Ru-C#'9�,�J,�Kc���
�R�o��ȱ��,��Y���`�l����بګ����+;���.�ӌ�kb�#/U�ۏ��a�$V&,4�W�'"�$Ȅih��X��W��2��~��i2^��v$8뾰^�b�Б�(Jϼ�S�l�6~�	���k�̓���,ĿAs5�-���|�������*o�l��!�t��O$��y�.�X�!dW���.$w���~�@8�{�����ё3��.H�q�h_�����bV�[�y>�="�"����C�����f^Cƃ�T۸�TRG  ^�w��h��@q�ױ���/0��������_ܡ��Y�����x���8�:��JF�v	K��X�走�]K�y��f���"]��=-"�m븊sf�\�k�Us�¡�fh�R�sj\�a�GB	�����v�c[a�k�t�H��3=�P�x4��f5ga!���:�j�wyݎ;��p4Wk=�	� ӂ"�\_�_�f^C ���h����E�A�.�Ȃ�p٥��ٯ6�3}{g11�!J���\��@�лe������ye�*�e^ :�ϼ[Sh���'W�H�2�����y벱�@j��2���s}9Xu^r���L(����#���0�:s��)��,qz�՚�80C��'(���HB�x.��S �Հ��5�|���4��c �D񫄁��B_����q��se���K��O>�fuZ�]i:|-T.��Y���E�y_���:w��`7Ko`�씓���Gv��[�6��z����eۇ�!<��by��v8^Fd���K���(��0U��5@g�:0��Q�ќ/z�V,:(���F
��=���*$������+_-�P�	�޻ܗ��RP|����$N�{9Q�_�ZH�2F*��	����oMfn)E~x֞x���Xp-���)���7z�׎�.h��T����������c�J�����������s���?��"7M�/��N�[y�
�ʴ��om+�A��f��\�q����Ӱv�($�0AW�XAk��t�<�����_"�/A@*-yn��(��_���Y�wQcRۖ��l�^#g����j�Bz4�ϵ�!�65a�*.?��m��|gay@z�z~+)��6�d������ou����V�1U����v��=�VNiV���\����ؐ/͜���'��}�(s���
$[�T-m/�����ou�g����Vܣ^�'�N����>�2���~܂�@%���ne�pm���m�ˊ���YeoM��~(tؙ����e������Lꘄe��x�\"%x�0��d��������AG)�J�3ϋlLwE�g�*~S����WO�3�����3�P[F�k���ް?~�`�5�襧sE�Z,����"��F�a_b�¬9Pg6�v�^�u(�D.h`/޵�� ֽóB#W�e��E�5I���]���6{��@�;�&LjԞ�1���O>�o��/���f�T8Z�R�����09�F'�	Ĥ�ûW�i�."L�&@/����R#��4��Kŋ
���ס��+���9DL6�z�Mӊq\W�z���`i�L}�����)��=���<?E���)u�����3�6��"
�(��~T��;M����v.��Ց8c�7$Ԅ��:}<C+�m���̩l]Id������+y�n�����byM�(yȁ�@w��]ƥ���W��h���D\y�]��%��4�w1u��{\.SL��Z�xy��<"�$eH2�1��A��]�8��H�Jů:3ɧ�g��1��z� ��w�غy.��)���-�*	��O�N`w �[O�$(�Ue����قf�J�鈋���<Cr^�4�G!x0Ml<uFkW��R�����^>��/���{h� ���ʇ'sB�Ȇ;POĕi�T�;#���2�����-����p=aD<OO��$��~�ϘqP3"k3A��|��@��HxYE�!�Hq���_�ι,;��B�o_з:�\i� �p���x�_0
'�S�l�����O�iY:��Z�A��x�{ƻ�,�I?�N0o�G�+�Y~�Y�X����f�wz8�=�H,i��ө�=��P� Ŵ���	�h�H[�~�t�Q wM�\����E4rӆ�L�
=��<��?X7�m�݂�u�b��"����BV:�@���b�ԕb�Ȕ��g��z��;f��T���ݚ+�w߇?�J-�����P�J�=,��=y�
��W>\�NB�]b���;���4�Қ��̶��-�R(x�'���ϱp�tm%ëo��B���
��\Q�ȓ���1�&i�!�i}�w��&��}��2�s�Q�`���b�9v�=h���3��g7g�ȩ��Ӛ2��M|4�����h.�/&�X�h����Ȇ�a�@��V��E�&�O���W�YE�?<�E	����߽{
��u��!�-u]��Xt�G2XUѱ3����2�a�^��ӝ<������:́5�)~
@���GY�-=� $kv���q�y��cN/+�T�>���)��S$�Q�V�@�PS�G�v�D�ȼ��A �� m��A +T8=5n�m�sܵ%q��՛�Qgb�9�I/g�5�.�I��<ܲ˛�yZ���ݔRډ#�e��&&=���?�6�iZI:i�0_i�j,����!����;mGBz�F�2(�&�UB���Q��A ��������$���f'8t"%�&�d��P&�?C�wW�AX�7u��U\�1D:�)���^2oXKR|S[���R����{o�9)S����.�%ɣ��������N���(읽��$D��@g'|���}ך�~2���"�Ұ�Dq{Kq恫����u�8]c��x��`���� �J����*��D�#�A�jA.S�I�a6{����)��H�N��Ǽnz�um��(��2�� GO�8Y+~�8��YkZQsq�}oD�r�㢠�� �T�dkZ-00��� ���Ӳ]5�jU�@�hLյO+ʥ|D�4�ޠ�Zs���= Ѐ\����55ŉ��u >P>�`˞1D»ĪRB)L��N,� \���ɐ�,��mwe�R��5�����ڂI�B��$�s�r�x��s)5⑼B6����
a��Z��"�p�RM�b橲�q�.r���!��lp���fK������j�0�z=�܇o3�:���m/!� 4���]3�� �!<ľ��!��� �pJ�(lS6�haʽ�6���7�^�m�pX�x3>0S8n�93���`�W ���t��ѯ�R�ƣ�DK�b&&Ϻ�}Pd�&)_,j�$Ģp ��{�'��>�ҁ_�1� �;+��jwJ���c�j~�H��o�;(��'�{ce
J>k3�aIoI121e�<� �JV���nDm�lR�8�O>>R�B�7�o��{�n2�M��c#ϥ��m͡V�3�2�N���VM ��.�ǅ�%���;�Hu��r4q��b�Ǯm��R@_�OC�g4g����ojQ*��LԕB�C��<^R�OK\�x��۷�y|�AR4�F���n1Pl�ΰ���vqj\�O�rT��6�01I���x89d�Αp�T��Q��B��a��<��\�:��of��*uw��������>HE�8�&���,ĸ�>j����*��T���I��_uģѣ�$zS+c���K�,�JKq��s�x�<���2�R�)����˺�z��K���#me�����������ň�k�Y��[\W��LG����7�<��@o�\����W�u*��pr�,g=��/�Yָȣ:�<��g�;;��T���r���g	�υiK��p>��Rvܬ���è��;<��qxc��m��V
�Ցa�%���i2��	\���B<�Ab��!YsxF���4��z,�5@��s��]�G����ꅶ�l��z�}�]��*�"��x� �����}�yFuPV�fI�^�)��H>R]�6x��GaM�ȾH���o�����{6@
 ��sm&.�u]����ɞ�c��%�.���gm-�3�.u���n����
���U[]ٛ��2���,�Bձ�5>1*K�J\�վ���]��Ĝ��P����!�7��,�G�.��A���J$�{��bn�Y(1��u_�c�ں,Q+8���B�$��a3���nU�ڧ!�-�#>�J	R�ϥ�o8%��[p���~v>������w�;�ai���®eSe0�]�iӌ�� ��<4 GWord�guF�*�^L�"]˨��ͧ�Ut�V��΋Y�����6�+ �a՞y�5�ߞym�vj���_p��
���D,2��	q�ߊw��I�ς9ಥ>
���� �0a1Ã����r(���0�AB-�K}T�I���}�F��쟬�{�X1� ��K1���kHͨפ��/N{�����^�'��:I�A'�q	�J*TL�6�ڀ����r���Q2��RZ�CBM�]�骤	>4@��h�ı�2�#3�ն�����u�+5A�����{#��V�lx٣.�����`���D5#х6U�S/l�١{{)�ڋ�z��jь��4e��Z!c�*�v�˖��H�g�d4�B��g�ʹ���%6$�Ba�~i_��]�)��p֠y�a��"bwC������pM�у_`f�j�H��1�}Q2s�B"���H"��BU:h�ЁX
�� ��
�o�r�%�����H��y�L��*���"��aQֲVƈ����?���؃�+�!�eώ�@&R�����4ʴ��4��&�.��;[V��ȧ��8LjC�* e����V�0��#�jN��1=�	�\�~g������y��z���^�_�ai��᪇t5p����{�1X��*� �ȷWS1��4�z�ޕ�k���V�8��<�S�E�Mؿv���7*�[����8m�l��/4>�ZJ��H��8^����!��8�Έkފ�K{+�������C�T�{�P��{��2H6��'<��鋓4�O8XR*ܭod U��3�, ��_����{�M�ÅA�$�}u6V`����"}?�w'��{��ZD��g+m�U����Y�̪%�K S\�;ܻ�4X�� {�g��%�6���1�_ql)S�=����J��q,������"�3��+���F��n������&w_����+�şi���.Z�E�T�?�b!���bV$K^5C�j{�\HT�s!��Փ��K�������Y���k�ywN�H�R*�DM�y$kx�� �{P���WH���*�Ǯ"����� G��5��=ң���!� gD��w������A��>X�8 ��Ҷn`�t�oE����D��: ,΁!�f4�[�N˴���֑}�6��b��?lS	ݣ�R~���X�֩�.c=�`W7~��j\\Z���/�x��9���ޡ�����q�p&�G^0to���O�}6��o��m�vL0�c��%��p�^1#�)�^���
�Y@��^�R�e<���~U�	p�>���P8
X0+/((�x�4] KR�3(��<��l�Q�'s�� l�b��U_�tM��re!T���CM
�fg����r Is=�_R2�y�C����Yv�g����ܞΑ���&������{��c�����@�R^x�N<��I�E������~��O��E��f���|-��>�bE!E��DIǀ#��\U(��J�![���`�֪'H�L9��L%�0��)�Dz,x<,�o���ƭ�*�+�$N`�]�ͽś-?����N�8.j�]xR��h�o5�b����D/��G�SN�8ɿ36�d�/W���҅R����k'`x޴��6�����FҴP�HV-ܚ���l���3�2��7�!�,���2�D||x� _P}kD8|����)�!����p�Y�)ƍ!;!ZD3gb��ǐ�ℚ�l���=g<oQ�C�˷��,Rߜ�x(6R����y-�[&�k�A����F��_N���@[U8OȸC|�~]��0[�Pi�`d���.� ��0T1�w8��8��ش�<;��l}��o��H��G��g����9��G� �`k�~��q����;ھ��C��;�Y�K���-���"d�V����pX)�W���%�4%⇳�����*�e���׵�p(���!�x@�P-�u"X�"\%��nt^����\D��{�MZ�E��ϐ�����"E �>��)��J��]�_{t(e�����|q��L���ܿ}Q���77*@�p����um�}w�dМ쀢�؅f�'{0�t+���_�5Eu�)��)a� �dD#Jk�͌c�O`�-�se���]�� �_"��x:zi�	���O������m4��Sa�T����$�c��q�A;DC힋���Z���[5�Z�h�i���Q0?Z��ko��t5�*�^�'��Ռ�@l��>
���20�ÿ�A����y���5.��uN!�9����Ox݆TJ����Ðz:I`Â�����Ue�A��s'Q��Zt�i3h��D�`6�b���SvaR���I�h4i�b�k�Z�Ō�9�o�TQ{�7�!��J���H�u��Hʚ�'~t}3��fԖ�C��zU��\&۲j�FN�z����E�]�x�� ���;����JO��Y��4jltD��Ht��uW�E��
B4S_���C�Y�օ��i���5r�tyUm�IS�+��J&�,��\i�_�w8�p1D���y|���lX͇���9V�ψH��9Q�9	�	H�'���/�����)��r+������2��Vֆ td�:�q��82�26v�4xJ�C��LΪU��6	o9~���(�A�ҥ�7�2�NTN�w � ��l7���y,@M�TQ��	��ܺ�����_�A
AeDSG�C�E�������E �ip�Z�D-ur��2WkF�������]����X�\':�IMw=�l�p3|��H�̅�,0��*�����S� �6��Q�����)]}���f͔ =�Y�x���6Ӛ]v�k�{'t��y��í��f��Ñ�|)��q苦/�nt&𪸻�p�;M�f%6�B~?:J�jP���㽘�x���{TW��J�Mn�h��ͭ��1n�"s�:��=%ݼh��+R��ꆊ�/&��{{�&�($�N��-��0u�Ỵ�o&"�w+��
�we;x�2g�-dT��ҤC9�+��Qk��y�[�d �{�H�9(��Mʼ�aǟ���YN�I��
�3�
�����뼃�H��A͌IS�&���5C���{�㒈o��y4��A&=̯Bl�h��P0��g�M��w�mH����� &G�Ւ�lgq���I�==��c}��
�Q�Us�$EC�����z�JA�G 6��b(��$1�/���\���l�ڠ��y�����JѲ5�WE�.��w2m����H��-�`q�YG�R��K̹�Ĵ��fK��hEu�rn�w��p�M�@�P��4��F(\ ��>k����%?Pa���y$���~� v�6_K78} �p߹t&��95��' Y�5T^3Q]�y�j��؏�/�8���R\J��y��˽��b�U��is�����('�u4��'[-+@���2)}��F �i4�f��	u�;^����`��g�8n@��˿%����kG/�p4�5�S������PAP�J�����"���!�%繁�~���4�81��(Bf~�i�1�5��vǆ��&������Y)6+����Ͽ�d��R���M�H,5~1�E�o��?3AO��HO��E��lL�)�e����{�{+�sM��,t#NM�{�3�7�Xu1{"�K&�`���!���#6hwb	)W��r��T�H�"��nμ([���X.�嫆�|�G�� DEf����$�@ޒYu8�I<U+F1�I�3�+���ZR�Xp�m��I�V��&��aM����>��Qͣ��F��9L*��s-�sg��m�ǉ\��|�Q0�%~B�r���\��d�1�+:ˊV��$�h�ɢ}řUV)�?�Z6,�j�Ѡ��&�6���sf�X�9qZ��|$gS�Ļ*�7"�Jp)�/̲՘�S��k��υl�P7�;�g�&Z���ǁ\��9\Kc?��ܶc�82
�$J��c���}.��a�0k6��鼒t�`�Lx�?r�Y��a�h��A�����8�Ѕ�W��ָMs.$��U�7����� 3^O3�`U�������>��rL��Z���*}`Y����H�>I������dޞ���-լ��%y/$$���^��B�5�Uǰݯ"�h�A�l,"��A�`��li�l�?0	}KE�h�Ýp��l�AU�aa�q.W�E�dU��WV�$>���mdu��/C��(5�<%�j���:�j��@/?�����,a�?��a',�}fQ��p�r�n��Q�hN3u�P��1l\
d���4M���혁)Z˥�D���r��8f�80pK;s&FY�����`����ʭ�eD�l��t�az�]E��V̔�ŤF��c����Y\pb���偒���
uZ�s�I2�]��g�-sqo����D�K�Cc3��Le���<G�y���d���T<'OYi�fn{��
�m���42L?RX�R��!��ٰ�I�`����-B
{9ٿ-��12�'��IؤJ�r�2�]�l+^���|�4�N�d��{N�C�]�e {�2�)/(���B���U�)pD�[�aZo{i��H��v��V��1Z��7O���y��ԗ+��!r��E_=K�\�߻�0��T31�!$M���RT�b�n~�\�9�%�0����Ɨ��.hj�/����� �}�����X�~����{[�#P~�<rvy�b*�"�$���l����`��zuA�����s�i<�����{�'��ع��j�)�u�����29g���ҝU�9�	3%�n-���hH�z�D$�fOs	:'��0�8�q���,Ła`'��H-U����3ZT�߉�G�,��b��6w/��3:�z����C��F�e�� �:���o�����y�0�ov����L����h�cM�伀�����^��@���7�j��1�E�r�t�VlA�����A,��]9�5�T@�q4�R~�D�CH�ʡ���,vT�����T�#E�.�K�INw���I�WȢ����k����nu�-�p�b���6:Zy[��	�<Ӷ��b,�p ݓZѴC�Vp��ZYe\�����6AL��ֵ��(��l��
�H��e=x��MgSe�X5WD���
�������D�ˊ��O��d+�=̤{���M�U���L�z���0��-�:�����{�	���<3���ɰi��