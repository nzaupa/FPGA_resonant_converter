// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Cw3V9oh98BZi+6qExyRd0w3ieh4exjHq00YbrxH7YT+AtoLDkCzja5zZd3IvyYCgmJ/JVsZNxQuq
q9osPJtjUYW3QFrYhyKQkjGeDqL0G07jf9+6fYgI08Bn6B7nrXx5Zl4phcTsCZQcDoZhPPOXales
8k9HAHHb3iYVf+jUYYC4JXjlimIplJOiCkp1v2+OTGjmuL4szZbtDgKBf00l9QMTf9Xa3adAx/hO
NPG5R68EgthkNZWVa0TiUINHZYAf32OjLM59c2PiBqlm6QeuNMTOVXgeHjkHJf6jDMAX0iQ8i3FC
taEWDs7kNaq1CY7wa/vdY8vbVbpoYojlgiandw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9008)
vms/xrh4x5xkj+fbYwt4iiwcBWp+kgAv1YRYjXNfD1zQbxvVEr56h6fcV1alGzbfXZVdjiD7a0QG
Ibcu1YMK9lwFG22XjIY37Em28QddrberNI/AimMvVi0u0zbsAOhgAgiBs6lWrgPVcN7sGkTERacQ
WPyqzDm3c3uII7CF8Ng2/75HG4vMw+uIcsYEWefxF0BKPwFO7Ear/l4qu4O7RzJwLIMV78u5Cvo6
DLCpaBI67C1ZuZMVB58HB8CAuquQQivl8K6yqVtBnNqaITqv2rWGdmcfDzxy0IXlhPsHa0Gf78xp
utjhCeQ7kFrZsllnXMKfQQSu3y8coNoAU9U1R1g+ITUHPWd7UDJuQrWgJtUBbChnP+SmCavySXN/
odBok5w/NbCgjVoaJrjqG6ZbVzP47WXf2ivtI9YLSfyF/PCCY6nCp2GpnkmPy9okxwQ8IEQ/kOKL
bMXKEA3Qjp8Xa+W+thiFBogV7r79NQVo++brfh26ftEhGCt6wImeKpMHdVhF8BYLMAQvqm8Amt2B
XjSFYB16Bjo9kDn0XMPfF8CPk7hwrklJpVdoGK0UNBd9KjyzeEOn9D6SQIJNZbP6swLEEkBV+Guv
2XdqdUgiMC8G6CrDFfNhqig+LeBdmpX39dOdo8wLGzj0a4a/9ecVSKYu6Pzug1BHX0niCGGv6lrp
R1wll3HOdMinp+xVfI9GLN7oKhNdtUBJr1sqhVMX2SKUzjMSABMGxxb7NFG5a3TUFToi3DoOBjmQ
aGiaEcZaJ2UG0bi47pJylb1lybzR5BCncuCr3CiMXWpMvYIM6lQHtJLI5Qd1gPYR7G1RJ/qTaA5R
+9KZ8A+9n1ZJsu7zveGrmGkHthh/iW9mSduPGtnhl+oh8PIbr7C+p2+UakK0xVUzxEkAJthyYu/F
EFLZy9BYx/r2Oq7R4cPTYtRjRzhAuif38qoaRF/Xn5vRynW7/pEygc+6uYHczoB4td+Ren4YHYpv
vHfUKtBGUICXqO6EHrQ7tnReqefj5GYSGLsVm/pywP9ao3Z1STYuAPtP1oxpMpLvCsPR2qWJ9KXE
T868HD4hYW6aK14LeqPTbeVKgPWvO+2kxc1PfnzWtqYQ+ninDvRMme/FeR6AOX2ZdgdaOKWd8p1k
OIA6WwFjZpXzcQGJZYx3eul5p44bmp9bsMb+ncfS2KZIGmH0KZcgdzcGvKbiEJIdpju1YRsSp/1v
PKTyywUnLug/FJM8k/DnjgrTzv/rnP1guEtO4c6NKsjX9Q+bVdMTKbQ/1RbmssWOrsBgJS6zqAJz
14ZSogqc9SpRBbC7KpLtOb5Ip1YqNvZ6FDyuAtVDL6DORCkQJHUghKDLVZJidxTjE7oqag43iLVJ
gyYLU+Ikk/FpLhVpDO0ThOeVeCQlR/1xy5h7ixwhskFVDYh7k6WvuD06lW8w13FZ2AknDh/kHomF
zSNzr0fuoS3ESkYoiLqZDXKBQNJaVzAI3ib4MeJw8m1lnavxnUWlynyTcx6C/Sf3/gXtaUXp1g9F
e8A9Db5I9850rOFuwsgMQBLSpNt8l+TY81gbGsxE6/ATpPPk2bSY4JXNYfTPqYUR7V2tSICcQHPi
IYAnAt+3IMOby9Wevd3BZ09KokxmnTwlgTKyG6mYImehZaEQblHkpeI8pgIheK5jlUHhjXtYFZgT
ehs3FCIDKvrc3fl1RzzLIRb0GCkY8imuh4FdZUEh8Kf4RqXXOFrm22efYRyIm+bZbH1B+TwFdk9c
xGV8A4ZaA7s8ALIcPXgppCVFQmnAhsImE1W6/tpnFjgf5rOtXlxrWp3IPqE3rLvU0tQDlrT+699K
FZEgHk/xwdpbMkwYoycrj9h7Ueqb/Q/z/NMPIBy7grR1iwRCTnTpaE+m6eYEi4LMGLbCPyS4bI8G
vBWkFyKtM3rkvDD1Hyp/oDQSMY9n36Y62QX7VBRpGEaBQspBuv0gZ6wpp4f12kTENTpkppIWmg3M
bUpw559V7OgqFR26S1wpDjdsiEQeQXR5K0BuNTdJHJZA5Qf1PpsKfOjgxonvsKC2gVOC1p8I+6w6
vTfEMmz3l0x/IvUiOYs0Q0JtZcTZD5CP1pbbpy7BIrJ/r8wWrZNvSNIQcWTrL5Z73lImLQukuVgt
ahsKYXy/a/1nXn3Yx+3omW09vkSlhSeyhzODzce08fz+QuYieKwjIGUTV+pcNNerc1hkTe02AdQE
G8g08fpIiZiD0npxj4eUAIZUcjT4X04cwUCBl2b90xWx6k63yALAli3WfZTqU0+eQRmSVHrwKiDD
phFa25cwtNomSxFQtdvG2zz3twjjptbV3zirGN9k/1JULTLWNlFREzg8G2IsoGyulYX3rkBoAiOX
pIX21JlSdnPJ7daXC+N1F0FBhozcDfR+b1h68yDud41QAFG31OQJ3yCKgNDGWPaDBfakXo1OMEIE
AoYowfAK/OZ7iAZcMMGOfGIoDIScTC4NtVE0E5ACqFLomRgoucJG+uQUkHAy+jLpaKwRWPTHFd02
OZhnArchmoMgDPpU5eGQr6bxO98Q0xu0sHybnlQq6z58UKn+SqMqMbrWNi8t2AQ5TgF2CUotQdyq
MpdSKFzCrqtDa3fBICsUYp7Q3abQ+clTOhZqY24Y3ql3mQkg0u4DG3bvyxShuwx8FRokgJoDQqi4
EChQZqACG6f+Vi4kZXQxvhnKvGWtkEQVLYgQoyF0pj2MqFXMmD4fkITVao9cx/ovOgURYrBwiuNV
Ez67rEiZgWUe0+zAEYU/CwcnSiEaEkxlfuj8Q3fh7Mq+DgiZ8p/fU5Jhc6Bg3J37+xEbjsJDdUBp
jQAO1LtdnIaVUP1LjLOMg7A1ELN9wWnNodWH/uYY8Pm7NSDJ3/3NMHwWzItyawD2pVWt55lCxRUt
IK6dvI0Z7baxnMaUYf9RYK9xGejCfrjvK5RltY3Pr1S85TyEeWY3luBzv390EDzd3EXlBgaHG/ht
rQCaMGsGi+WEfMMV8QCixeo3R6J43y428MXV8JPvP1WyuV3A2qCyYaNcn4EKIzkcDDJ3YU2YbwHh
sipb+s95Mh7sUfxAHFQbxV3b/EodUT7bj8hZtiIHrCS99WWfy3M1MJjS434e70VUW2sM2ALUXife
Ub5MOR1WPpfsCSAYIODmhtJq/OYanN7i91qkc7mV0wy3IIl2ygNyagHWK7L6ixWORo9dHdOHJdqq
Dns398gFPzH/XCfX8aSynivzabYCSX1EK2Si9sH4WXxGZ6RwSBj9aF/CZiYX0k2qIA+9GIw4Mb7x
p/awc6sjHOVfzevKzPLe/yT0pg/LV5XkV8dYaVO2AwenMQ/syccmbJqE28EyZdkSvdXJWjPTYeyY
Y8XUCrKMKT8Zfsy/HPsvnsysdjqI68dr6U+pcZk2x/lcI+QEILgilZRHc6ZuEzTh0eBD2l3DKftD
RUxXsUJjkh2YdRlwDIitOFWn5szhh+ZqvcUIUaFrHDSRpC9egCN3J/NXsKfGwZEnAd2ah3UG/FAW
A/erAQkY7r8Q5KqNE6c2XIMOkZy2NHmnPggO75B2N+sO1JNJM2+3etpq9zM0kGvwNb0MbR9411YE
YESp487wuorQ8+eIAfjdqcezkiK4J5Oc/4l/0Og8xXEGGHQ05sRSuBwV8Gpmp93SQv+ADGP0uD1h
A2PBAsqMnRSB2vFIiA6cp2CrGOj9YXUBhtmlR4RrZOaLZZ+xHKhQ6T9ObvACXbwagb6Q11Iex0hQ
cH1OZ3LCuwf1QFiS0iGGZzQwnsNk7diO88ro+LsD3hrXYtYlW4UTMjzLPo5HdKpX3jBgfylVgT7S
MrlmvsaodWZ5KA4dg9wXNip9SfgFfStnsRABPcbnZovsgEtmbnT0ieRZAcVQRv8D4cVawAXZd0zG
SCYTPgw5bQlnf16rsbjU4cSqjM8eFNTuZqMz9zBV00h4fxiGeH5cvgK6U1psQVIo35fO8A49uiWs
W73oevQu5jmE6/gxFL8aItkqJgMrTF8Hm0XQ4/FMSpGbOcIN+UBjY9utCgltIe6ed1aWYUwGXd0B
AMrhVu0hKoqXSL9R2OMOt63+R7VeW30EXbdrauf4aQ1y+/tf0gHtoaBDn7PZs7w3sT3rIFF4xnhH
wdO5SCfV7zrEfvraKuqiWnxd5opmQ6fq1pFXUfC9MVb6BT2QEGyo886Hx+z4djPLZJpljhyo0RlH
7Ws9RuV7J2vr6KefUxbgm60UCjHS0xb04TAxtTXCVK9liIdOEsaKpSAE+9o6EfRNo6gioX1a2KXU
uQwR6VgV4b0gxvpunuFSrPx0Or6g6TDwB2yPptDQaI8X9homT0E5EbRDNIFh7yi0mDsvYflI+C1t
lK7hqOFOeee9XCM+eaU7P8KARihNRtgzpC5MhbyZ6O9XoR39uWeDVCv/isi5iFC7K3iUNbUuqiMi
6YY1+yelvkRTYgwsOLu6JLDekF9S47nhZwi119FLU1LGXvl273sm2DKsqXoxitM8lzVpXfdqbna1
FkMbToGh47YjJTucISuFtk8oQ/orSfuYiuTBjBmJq1+X/AFgLk+XblRAjxJQcvMFhqDy7TodrIJV
tL2v41GGMN+ZllnBuTJMRvqLeKA/mxYmE8gCso40+ZSvP+1UxCSYDk3PA+G6y7hEkSodmA4hL6D6
RanEQYR4LaARx3O0Crj0TQqqMediFrmLbjw3RvQTxSZ8+HfL4jZNxh8B3vPVeAY7LPKjHRXITm82
FSFYILfc/3t/1ET9k6/q8E6rnHP1V9MLrJY+FeyWv9MXjNRhJAy1h6ZrKA0TFFvkPSRStclSTlbf
juqyt+bmlnGUEsdB5a0RQeaZK0v2s5IEP85KCaV7I9iqk2JVIu2VjgxMNuh3kio8RrmvO/nHE5VF
Hl4KUthHm+i7jUjR/+SIhN1WdrLqHdvBB8Fgdh9FMz9AC1T2mwHIadjqZEMoTIGBVTOCyiHW3SvX
Puimbdtgrmx/fPOx1ywclha+784QtmryJAwobrr8pnHo0TdPr/Jq6bS7cr3o7PX8ryP9ncM0jKQc
2wJd6GMAXcJa5PUmlsXMSHHp3hKyI9CIb408ZXS+aG1RxKGmJm/pYA8FC6Pae5p2y+1Xiae/5n4u
Pd0j9rwQzKxx5J0p1w5L6GOzU6sGJsHs+yekR3aGtWvczk7U0iaUJ+7pzahxoMB6mOEOsvFxOsSh
6J2Eqgc1fdQP7Wa8g+xM4KQQj4nqVxG2V14FU+lpcWzE8OktqjwFd0OltbNR7l0NLHWWSjh72WXh
xi0h+mufBoYVRZneOOt6GhyRjT7f9R3VqC9ar52q0rS45FE10bdke1GBuhhrsTgnvYM/BVFpm//y
KFl8Q/t9jHYi+HbcFjt3Arsbu1dtylorw97MWEsOS0MGsmyINO5rOL8eRTRQjrlwKdMHjgSP9VGX
OyyIG/VWxrIjU5L4BNC3uqifWx7cQHKyvnxuGj2nugaOgORiE261mpTkMIfaq3+kLAaDyszDwct6
KidWp50a94Xdphh1D2wDiluhyymERmeLZ7bOfAhrI8ehS3SZfROKGR5iLI9/EE3pWa+hDs7vSXzE
tddvzlGjgZ6Sw1wrJyizS4HKkKjn/xvOu/pZDPw1Il+On9o7W9Z+h3SquNcIdBzY9d8nUtcXy1KS
1rE+abmYyYhBan5OU9l/7CUj54x3TkBDDxxAvIpCo/ndRHSdkA157naKzI3WtQWup0LXVWc9g5El
M6IZlJ8atnbgHeFv3+5nLqlMVLLRpj7CjzXU8Wxe8FBul8TusCqzg667PFUVVm+bZAnvaW20bWnY
gCVMq6rhHa4Btb9X0IYwf+eTAVcWLepSIrp+pYbCKsxFyY6h85PkDpVpn9QKf9hSn+SA7aAPJ2Wz
452bTICUsEKsYDSA9NK5o+j2tqUIrhCcAp5QcWm6dxx7sbzjRpVixG7zKiA2qiCGRCJVV80sp0Yh
dQzKn5S9+1yPOmCp7avL6PG4yb44W/qb8AEPVRhdP32flYVg+9r3dgFDrhl0ED4eyWQaLjfp4DbM
UwiseFp4wOg9l44ku1lkmpd6kLdL4L214aVCCWhhNmUtwMTzTeFmTG6hFaMnJLjakaKRABPrCP7F
xd9N+d0qGUpa+JENCz+s82s4V31VEezy5Bog1PFi+hf3U6C2W/UHTJDdVDkJJLf+qA+L5D6CNug4
18CBu2kFpuvyj0u91SKZdgFspGAVBG2ZFAi1gf6aWrbqT1GNyKF4O1x7h/FA9w1+6AstJGZAQG+E
y3zPBSxyVDMLLQnxkSdPi46psAlgBcwC6KwEfCAmcwkZudNBzTrKLUMLHdAzWI8G3mncJkwkig2X
efNRqAg+IQipIFt5+BMv2C8FPyuel0AaM2RsZuuHkEFaR4TtiHJJ9peFWRBHKfmUHj2qzUi2ccSG
O8aPGuU2emCctsAuW0gzQIJNi1+oonacrnVpR4wmASsxZuePcokkCppL1Vo1B3OH01DsO+Iysxlk
lmSnJCR+IjUeeGJpFCb5Vwv8T5V5lhBtbFXhjUFbKwSj3llVrIbfeaGYn0Z0ClvKOvwxMlt9FQCX
HrHShk2sIBWZPLXMme73IC7wxRLtEv5mvm/b+eH9FlCf8cbP3IJ2J9UmphT35SkeuVTrFRSz5NgD
fHB858aWesvAvTPOXN556sxnLUOh2KODbehFT9HyG+1UAYlpvWLvkrLDOnFERqdCr1BhZ8pupIaC
cWxBFQlNoIJICjTVWCkanYPru9ukqnUMBymWXkOsvg37N8AwiJoeWOOLeZb5DPU21rzZ35puJieK
JK0jbsvO91aWLKPfkPqIC/c5BZ/u40KecnD7vfgiPYdMTaMjcbB8nD7V8R+/pylKcxJuQtCzkzcn
7eIWTLLA7+ziVCJApXBPo2dW46Si98TmI70a9epDtXCWZKeQ9soorAHahoZyxCe6c9vJmLQvKRCF
HU+IMRIpBsziT165gTuXDZSzMvHdiuNcXVqk5SXGFj7jnAV8QXrZ4jiT4WxUfafhx+x3WwfrkC4Z
d8dA3ZwiTwrWNLlJ3eLUsGER1W1B2632B5wRsQkfcXVTpzYIdLSci8xXltBtUQocvyxEnxCSGdBu
WUIMuoCM6kLHCQKSZZt/LHVju/HHnPKj+1iFh7ns/j/4WbdGUkDamKeOc0seGoGx5QC3k64gbmic
AOYlsHihegA2eimmhQI7cvl1s72gQqP0MGoLyqlVmxlG1Z9s2uBrMNLUGJgUXiyAnK8AThrlON6w
+9Z4Pm/Uu8sMX8euOfitziZxpBMxgi/+q9jcrV+KOc58tsW+mJjXCDiy0Ok8uwVIaxC5ZCABDr2M
L5savyayTOFndaF2x0KWr+MbU8wqKBTNRr4FKo6Q4XdSLFK4c3XfCYru2oTHdO9LkPdLPTQUkjX8
xTt+jN6kUuF44M7GCw7TPqhoa/JHcXohXBzvc28CPaAMqI3OSnDwaFVPYT/7jMOAKcp8njNKLGUj
D+56cLbTZth4tSRLRQEld8mKSytE8QvAEiDeUZ/pEin0VSKeo7Ov0RAlWS7sjtkR6UGzC+AqG/kg
v7DHbS+MinMcFm75pLipnAbGn7jduBViGEY2mY+rkBmJEYgrN86wMyUb04gHDVhQOfEMkEV0HjGv
1RboEUWf4j9gerkPz1OkJ3B6fDJ78NabUnkYuaUFAjthrVv8QJUywy8m46mrsdeYf7onQWA4/8uf
19jZ3kD0PPr4eCtw44FCvhn02i/1qU4QfCewM3LDy9Adgc61rbgYcvP+UoGmaHEHJBxbaZmZqyNN
Qte6i8J7bUBSZP/papFVYnB1CQeojIvthQPdmBPIz0FTs61CDLmecxLhxMEBtR5mhPjcHZ1zQ6Vj
9ZIwdPtpOtS0/TPde8AkL7FWvWoRDKGy4vUYEjiiUtFwh+vpbeR9m1ScDMTVkCbmJcS/cU8hortQ
65+fzXmMStXlFqn66fyCfg0WxfWeQRm+c7oIgvdcpe6yog/BSpqEbQ6rQnud2p9D6C2tPlJubZ/3
FpK1vYa6OpdNRGUAfW8fmSK2Nvc/rHW63XnNNSpLCJfBdqDrcM/GllZNtGzztryqP6jsJv+1W3p2
S0HZl2wrfRU3IzSPYaZvbfJqHOctFzBLdQ0KhBcoJBSEu0GdFzbuqB5dwsDLEgQ9MQduxcFTQPsR
SNWV8MH8ermBnuwXV20gybogg2xUjeN4XtDUlYuIwyUddp1B/jIDzg4g7k88koIc6cDL/uRgUjrk
vRLz2jb+5hzOiYu5UBlbEwSCknl+fL7hfS2sC1j4iIsuBKizjSOXDllM904IfPrwLuqzxmjotB9r
0PSxiW0sj8ptOMFdlRptJ1bJ8aZMBCln/Hu5slRjWW8eh0HZEYZ8CJYeHzTEr7NQU9SAxy7rstgk
uTZikOEOeqGy3oB335EAi8p3/TSI2PbT2Vpu35WrAjrGj5YRmsq3dAhWIyFR9LLVS3SsaGfKar0l
K7bzSL/fSm2mmzT1uvCMworgkSX6D+IbuwfInGNAe8qftumwJuSZfeeWdneHmu2TaFDy9/JVft09
54r92MoxPAOWyYkmB8/Nj98bcvPy71qjGT8FZ1RwC7M1L0TIjvE8uLaVTyLIKTKfyD92nc2ly3cp
imjpJccH1C66FJEbkuF2wNYPu2F/q8L6VVTaWt3CqGiU7IOXgU2vy9D4DEvwWzfEotH7ZjatWCoi
T/YKlFFucPqhNIM/PGKm94B0Un8E4kUZAvT4cO81NQvBsJiIHQjg/326Qm0RInRu2PfB/M0WaVHY
WjRtB3S2Eaxds7z8dEGrGSGstNDhvrBNTaUrBFsMf7e5c3BwMWGbg5hfqQ7eGXWJreJoTAJNcjch
zhbJ6xnI8GAsMVafDvRNQ3Fm1v0Z/ajkslAQ3zCq9KjOYxuN1dh6k4W9lua/ydMyPPOwNqftd7qC
AmJtuqIXds3GIIoAFaS4NYVaTOi7s80SqxiYtY7MJPLq1STEzlaM5uIyfNAYlkOJ7S+10yl2nlkd
UDr5vrCXxRovRJsIppv1qU369f896GisAtTz/aV0TiWX31vpPNHsvMpHaOo95U/vWTLu1p8Wuszr
s3uYWKqlfQRB/PTmpj81Li0IzVmoSvXgpT9t78jZfPxWCqGhvIu83PwAxUwA8TBYBiub+p70vSxS
fKqVosDTyb6wv+jgZ7vHjEOmqqojlFMG5DNsCD/DCSUH3ijE1MYSvVbumpXtLBsimnuAMKBXXNjU
ZFXInrJJDP2rdKpdrIv4zJz8CHVbhlcc4P2P/Uqn/zx7ogEpnaS6ltwzv4BJAj2DJulWTkerQKQV
uf4NTdHpSyO4P1WAG7lRtkwP/Dr/E9HzP1YR4/MkwHJnmePyQldeEJRu3Q+VyUZrsH0rj0NZm/F/
LKJtcEaCoFlJ5sE2lreHvL2qPX7KNcXORrSChSZVfpn44lfSzNeHxTzZGGCvNTd/fcmgRP3kjtC0
d4pimJmFOjsW0CdR6aVA2EB/9+qdASg/vLxylFxRa+Ogr7JoKvQnEKKH0IKd5q/1XtbhZiqWUHZn
1gVEhlkmLwXFNuxUw9e9OnU2rDGJjn2brnMMEI25GX6m46hjbF8sFT9dT8vphZ3cf9L4KN6CyRXe
tQFSjKVcQg3w859AlyBpnAyTy9nL3EkszM6vbtphOZqMEwqoxZBQFhUVsbAMXL/eTVFcz/4J7SSg
bF4YrLCk6iTp5UyR8qRMsTVQ/GVlPtqzgqBoVr2cXySJxOpn/lMAT2I6FMr3vmp//gx4h11yxeeC
EABcxbGjg7+TuZemDGGxGf6zED02X5PtNLjGP+evNekU/VwK7xSXDqcUNArcP19PEvlWs1fq6pUT
Ysjhi4qYrLWzWiatG1V5GST4d3rypVNfrYr1j+ODaP4i/Jxsbo4r0MgEoCGY48iBMtidbe3Yvhbm
uSypMLO5vI9HOHf3+LWUAuPpKiUE+nvWgIDlJsmsTNKDA3v0eEPoxFbPuWiXQ7LCvKM0dntkQEoS
FT2UU1X+cfMd/iiOndKNkvy3Fy/i2XA720Ehs4JX4SXR8K+qCcYrYelDXbUIIx8I7COZ+E8OU34s
F6ofUsnoLGkh56Nzy3NmcOscPS5TvFaIH2qQeiD42zEIhBtSnL3bGVZGuGHbgYjjSKwLr/sMaHA7
i13hna7fmGcS/hlsN5baO8iCYH/XUzE79O2lNkfEoI4dqrkna8iiqDojd8EGYzuyLmr7nc/s18ce
pJblMIm1EoZBvz62DKxzxeI2QyjLJxguwGu1VmT3g4HoHLi2b7eq3HZWnGDRYpMYrhsvsAfhX11c
GktPRT4PbgdmCDJbNwYMNUA7W71NJiKA+U/2AzYLkQRncTtNthvLK9mUO/t6nthh09PqxMAjM2SQ
LaJcpb2zXGahy91BTt8fq8mNiR4gn2XbqxTlqe93UNJ9QSFBGKsppWSUqTEgS7mpufJRinDxi2CO
XyjGgAi7lFGr4QsxgmNTzWBQOX40//1lyZMPWQy4M4pBXRllvMSd87Pd27Gz61EXc2G1o4xcpMfq
b6RwoZnhjjG7hgNsDwKCYChktdWATt0MRfYzHPzCfXfx0T6GXjWYL9sbSYDppIAuOY3oTxhtO2GL
JRgAp232ywtbrUdCU8hHU86FrMfIwFlBqo5uhq3krllg/qjDabw0kc2RB+5BaotsPJvjyzLcCNca
20FpG+nPW1dCYaNzhJi3ZjIpCmlON0iqtdznA+S+tJnGfKDsftfZl7HqCHje5hrRqq4FtuV3AKJ8
KIzV68wI/XKlRyAUxVNMTi+RLod/oSys1y0+nB8LtoXtlZyt9ZwHr6wXKU0lc9Rz73MKsbMR3Eqg
TGtLXyTzFDFQWfnr7IUs+inWWQu8DZ1DYsbM/ondHImHvOen13E+8CQNoBv5/jUN7QZhR8cP7a4Q
DB5l8YToRbt+mkbkDM69HSVpIpGjE9CJpU4gNll7ac7MyAXFqmOfy6TpuqKWORRDESXhWr680GzH
UM2qBM33x/UsVcB+ZT8LkXuHiDYqJYFQ9Ev1RDRiCM43psxDbOmwMWbXayNTzZJ9uX8zwbptT+pU
QwlpR89QAKnMjokS93E5I9vEdyOqImqT5vK8rTICx7iW2AN0AkVEiPmW1NyR9zLr8OL0EEXPIJ45
e9ewU6rgJTu5Br6QLGMXPVove/u2QqW2yo+BEZJoy/Hk1QlAF9UiGALgkMKQI/nH2a3/ylG7xnk9
kQWe3CSA3MG8DJPQ/co3Ze1w3RP4fOAZJhkcDVYYi2p4njFrWgCBxFwE9NN9lHt1AbRwIwyXHRJC
fCN+2IZCjP97n4JAKYl/liEZyegQ4OcXea+4KjfCYCmksz4WCAOFfJ99K10bLStODAoOgEv9iinf
+P6VDTb3fcIPETIgjLRkWmJrYDzLOTKi+vPiqZ87DNdxvc4tazkVuaRGdLnp9ZZqZC6ATTneQXff
QRSlJySeFNfbd4kUFAjPX0TKvL4ppB32buXvVVYxtDvWRZDY4bA+4qte4kZAwWF9TkoSGncrbz6E
iDR4qqq53PzrG2hxAk1SM79FNjVIj1L7IN5OVcuPJ/qqbzBcaJlaJw4JNIBg1Q4SvzKkDIffHaHM
UuSlPkTzsbAP7trBaL1wo1r8Lx+9JS9y4VQoXZjUn6o8nppDtMvtUjW6wypLZ5HD1oXvD7NI6Bu9
9wunMrclxmvGxqGJ+7cXxsDhNXtfgjJU/OopuVlG385ey/mYxtjxy1FuK1TP0SsGz6+HboR4bC9e
hRnmUqNUhUryfUD+DDyYFQkHZJKQXmtwpf1eChKgx2mN5JBuURPm2VXESZ53OeEtx+8ol3RqhjKX
gGrG5fz2TgsPSzkLXJ9oN6dMNQnVTsaq2n8dx5N/otXDQ2u9fFDJ5s/YOxY3yg6Jq030OlmGU2IS
BZY48OwHOuVFzLU9zZUU7H62F5k/RmGlmLhzscD5TNb0U9tRrTRV6wB0cgaoF/JirwTA28mG1nGi
b0bGJDQ9QDLhlTRrLum3OyabKypfM2boPJgLFDhqgTTyjNVsrGpO0m6q7oKmumLROGzRDiXJwfH6
0zE=
`pragma protect end_protected
