// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
P3CgKCeZo4wUXEnsJnbQFRuaXVJVCVoImcB1hYlcpsLUx0Z4S79yLRr2uesbi3hdyaHIril4aD+e
qnZIavTmFx5ZkLUc+qoKa4AwuAOit/NSK9jq26ABArS8gnXu9KSbQJy4rmB+R7ZkmF30zfGppWwT
CDIVpwXyf8IDf1zTnKDp6hYczN78+lIU3hgHFkrm6QlW5uljZBe1Uze786IP3l9mndzVbWUEU2Ci
h5dDDgFCCGoXFEYC7tN7J/rtIGR9sWlRzPk47s68OQWOWtyVajGRhSRcUb7/b92y99eTtdjLpidi
/izIgV1R8Cm/Zy5Xs6e25mgfuNzbnnBAHrYw3w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17280)
cVL7QziwbzASrCM71MWkekr7PfuKD21pRI7g67EutmuKZexwi8RlYqKEXyKHXSud1BMCGtqZM5m6
XC0xujxSQw4KjV4hIb1qPPcIveL27+7HURrvzSwoCBeAk63H8rKZLDejKYe+6wS5Upz189soOeWp
MvZCY5qHEth5xwaKcwzgwobz+1MRPmG2HHKGebPiQ8Ly/3OhowSoZ2RXzI0G7yr0fcVVnp4PZdCm
LqhwwQ/xRxv58Z6wmL6bnTXbY153AJJjKisPH16hXOzdXPGYeaFYHcLrgh8hJmpD04cKH3sQ/LNp
Qv0mSHLlne9gVwuFuqx6MIb4tZVC8kcMBgD+q9mus5QYOFDbAFz71XDTZbVe5lmCl7pekHVcqzCE
nTmliaroBIxuBFKteWZLkpfM8FYUosce93zHe636f0v7S/kVt+4ji7X5eSF93uE8McPwQnxuKJ18
OOzTWe6eNFIL4VPNkDgSYbgGdcDio6Tf85jjZPnACaakPocN31LnslIV3zOcbc/BLDc1TXa9Aifm
7xQ2ExIbk3+HDAUcEkMmItJcPcaINq3pgexEZPeO7V4laKIFsFgvPCrxD1YUgw80mfll0rUwd7WJ
CWWjjWuJRaGdMd3xxK8aE642zmgPPiKMmc30ajWiAxSmnjaJLK6BexwmC7+LI0MGDSP/aZsShDI4
1Iftt6i+pG81txvLfXY8cB1z+rugX/1oshNKRINv8KYIy902swic9PQtZJODBivsdbP6ypzyX+FU
elv7LTBwemc9w+j9q3gHB7TeD+iyQMo0SnZG0IMXi0PgkcHasGcoMoY6VLQthSevCuWa3eYy1T0O
61DuEIq56q8gqRQHzwblM8x2H+iHc598T8ay2QQ38HWpz6W/bUbZIUbNjNn7wDIakQlgQQW7MWFf
5Dh6wsvHzpZyJQkeDzMr1rKBiCptzxpsoYHn2R4axV1lUo3jFnVEl6ScKctcIpbucybnOUJ83gVl
RcBwUSFytvt5MJppT6j03tcrG9I6QykI7BfP7DwvUCKX4dxwUuUOfmpAUc+qH706TozYLmLQnzkp
AB0z5N5jVjI/D6MwfEknGhi3Gr6NjKIycYzBRJ1mFJk4lsnyP3Mb+WD+s5CE8z1EFD5YB0JyQRxZ
n2DZM5VaTqO6rRs3nAUK2A/gj1Ba9m4YLcZBOenqOZ0rQjMPNMIQvdEoPpKceKGui0NCUiFFuiQj
ftHLmmNgEPEgKRd4O9zfOpiUIkzi3x+wSsK4AUJXBnGvr+p+dMdODLI0+CuuxFO12Oe7pOWUPWZs
YsY7oWEG2gHKo2QYubKKj28HMXOHphhXPivmNhSnoTXAOiUmVwLNFtxmBa54TQmjnnY9qiJmbvFq
Yin6LRnXGtr+0ftvIW1uBYq7XbRBHhMhv87xs7ecGYYLO15p3b3X5xOsqt8qKQG+zT5Sq2brPm34
MYjsWVnE569RKg5PCx9cDlh2xcak4iAqYx+lOf6qrlfog5F+x19l/ZOaW8ho9fOr6CQQ3L2WMVS+
ChbCqQ3iQ1AH572gdhMtGtOeRosJYJ5TjjXE9WaZt3GU0IYaJd71U+Oi2QGyJGmq0UxvlWAtrHvV
0qzG8JaIuZwPKoNVxui+T2kAAhzbEeypUaqZJdWxeW3kicVUGNLK/26t6iDQ7exzb+mXJ0obDmbh
ocL+6/dotfurEvd/aGvrI4LFM65mzRMPTfMbJEVsw8Y9j7JyAWl4h1vxH6PI4QkcOcVsaW0P7Sj6
hQHT3N6WZ+rgikDu7coc8ai2wSTQz1iD78RvXLKDVWHYDfMNKixLjduXZvX9zLwE8nyieYRxVuEA
IEucPdYZSjmiDhuHek9oxdHY7+lw2x6fJq3a7l0UCZ3udFqI3Kuhht7D8qcbnp6VJDrd3ZODUA5K
UO1Q1pWOBV0Pirvfcudq6LBxgfXGxVQzHRZMzKFRfOVQC3RHP2NDK8gjNavplO/IX6e+7aFDi7W/
am9N1Q5HdaMlsuQOiqgCY60+uQiS/QN2t6VQXnkahE+o1W8PrVuHEBCxgUGT99zE9KD+9qwNX3HX
eKQ/WHkSZenNA5xrufsmTe0NDQkHBwkwFYMD0beecgRs+TbuNVxf7lWIpXh02TmvBsQTDvBu3ovz
/kh0NQLmGDwH5uCgtWVdrcqW6PDniWORPyAhF4xGCQgRPrHjOdJr/M9jDp05Sl+NVncPzzedsUur
+Yg3I0pCK4YiZp6YstLPrba30aD+MGv+l9tmghHQmlCbldrNjCzzqw0uiFDd+TA6G6aMGudWNWxE
PonhG+HO7VQDGL/k2hyiQUH6oEeetBXYPp+XeQtOdyFXSV3AvODEYO5sCEIS0BFy0l0Cy55vu5Ws
4Wc/ItHA9AoeD80cq92XA1zfEJ/30+p46hkDamEWrou9e9VX/dsDFvFBp822GtjSOuHiRDXQjeUl
lsUUw9u2BKCPImxTA+T2EmpEYAT6yVtGSETRCrwkbFqxMAccWmAiDlAH20X4r4Y8f7TyhLdPW18+
PTbx2Cl0p9OUaTRfcVdqK3ESCuVOm4eSs8WrHg3oFdz5uyOvuQ8Prn+laK5JbuZpvqzYJm/jZ8Cn
6abEJsmS8KNtVgjJP/5eSrg9a+aCT1lR9QAIRaDpiMcwr5m7kratMTIyl288aEuM7k845f1HUsqE
DpM3C7LtwaWu+bsjl0shSlgTvnHpBszjfoqTWSV8tqBpy6gSBT/TGjY1K5KeRAZgdDvFBirLfCw9
voLT1wiWrSsmkY3IZhE8MLEkNS3vkvkpoQdcey2mspxEIX7qMIqx/PX+3YJO7h2RfzXRWXjR12aM
MhZ8w1gc4l3BEqn9XfI8mUDib2MF4JPu0d5pwaiCjLu9yEgR0KQFvuxcbVd5a5xgLEKQ8z14ZrrX
wme8+qnTxJpU62dbplZDWZOp2w/famWCKJbuMdufbt1cnIUbscFZEVQvDdRxgfQp5NX9VCV3tS4W
qUJ80ZXItmS1eXF160ubCd+GDse+z3NDGduE6k9WuwHejEKGhVMtxCh2DtPM+ygrW/h2To+eNGh9
n9zAcO6rm6WQEmqPa5mhOj81x5PbUTJaPRcY5qHt9qYeelHJIR3I336V+1NiiK/pecwgGwcB3qBL
23K3uEQsqH3RsYcaOEOrdl3x3UPsrCiKq0eDlXexEbTX2G/2ZoF/ywKIj/NZrAifuuuE8ISYmiga
mDdNoWPcFyOLOAPJAzREt/XuoeXEOkB6TRgBIiDMtzKR79yGW1lYkP50MCbLbOL5kLn2oShbBc8H
G4tz9kDpGw9M5WbSFJTiijwDEU46STClm3S7DB0bgi7A+KVVx+s4r0HfI9LtfQYOYKZjf19+D49J
/3ZPruR08y+Smd8KJ8FHeKUipVCiG5q5IxYSVkJF2K88aNqADjhoh52E6hDcAFgzGD3j+MCmjeJX
dZVkwcNIClpG2F7raT4g3Ju7GZpL3GXWCriF89tVSOUDySlh4Sz4d61BflOCedcdmnIELx26EOjK
YmGbOPrtvr5LZG1O+C6OXcpYUjn8LgNsmmSgUbuRdGWXUsDFVv0/6+sAVuLQClVAFdfiPJN2q2PK
foy2lFOdJ03BUDCzyHh7kTthLRDLO+RAMzr7/Tk879eEqDVeBPQR2qlwU3A4ondGBOE7AKh0tit+
jI+oV0e9FQIw1PeMrF4FhaF+hqM8O/n2PSoyKOHvztY9wiXeoYSDQvSv6HkrRR5eyKPWIc/aZqNT
fHxCpAQaZgzAGI9m3vNiJFuZnWDSS6GRCG1/RUFUwM+nZei2k5OvYeJxZf6UcjPQFdHtqbveM5RX
zEBxBoXkjKrNAoBSBOQZs6V9drtwU7fSlDTj3HElWuHDe+pJhHm02O30w6zJZj9f5E1jtX6KIy9V
NiIIEhjaen64aTDd84onTHFz1OFlp3xNSI8ytldor1R32aNF4NtRVqphat7KcUiFpCz+YWZNrP0o
UKCXZI5r0w8s5kOlYdoVQRLIZMk27wdM9+Ry92rIkZl0lZU6x6SxI7oLMyiGQqjx+y1GF8Im52cA
kj8DUwz4PImvlx8JtiZF5b/IlEZPQMlnGWCZoo/vyBlQK8zKw3kVdGVJOp8/cz8C7FH98XE7xd4N
vk8MYO74FKyZrA7jCy2Jx9PRmcHo6bvjz1cEcYM+7spOwuKdDRQKBQQ9ec6qaYHzti8mPlBIczVk
ztad4sEXztmazNw+xB0sxUK/cUrbuYwt9x0SfOllKnoyGtIPWnBc++NJoPbCf4NUWpo8t4ZnfBNP
1njlJnHQALmHnszb5xokHf2GVcQGJcMWZCdAq2T8yAWbN5O48UvC6HaGunDqMPdXDw9iWDKDnvc3
xSsf66X/fDogr4QpDc9Yb+6A9C62vzYJ9IjGhUY7f2zMO+iawxvk5K3SN0gEca+pF6K/HvijyD41
N1JbJRxdnwiAxtOwMVLPzcaWhRM4wpzKMGsZcjw4b16l+BrcoGsYWmz9BPd2IkO7XShtFMTtRT3N
5h+eToVYXdqi0+0724bBVDoOcj0xlpFub4CRQhGXxjjIxOLNJGhcgWJsU//boKPJtRt3UTbkNP8r
juGjhFhoQGvaYidlbs1q1IhQA2hLC2xoBCktj8EGW+2Eba6W2Eff9CBETRi0hm5Ax4CDkzBnC4BM
0xeSHbjpsCXegsBKsBUEWQ8GxUCKGAppr5d4sgTvXugqKEXnulRm7GmMlSxmDiJNwKwnMJ/yC1Up
8HW0JhL5epYHR/A+NyoMeTAj81Py4dBitY/S1Mmskfjc+AztyMcV/4M8LO+ljD3OiCfrcej94ulo
Y3c5i45HpnfHl0WZAEGFPtwAxH87N4gmDKq63HDnH2TEct/q8+doeSLtDtiGKkJj8pYLE0GK/p+W
B0gKY7lyo4zzx1QdpxsaVGyCEG5sBG1xjTwRkCa5vk78K+slhlfC+NMozIsRpCYXXSUOxhNoQb32
c1GrXn6gmVlTxIqHVQjsRwzaAiCbRIMTbiKTkPJqB2+7ymZ8C5uzQpCA2g+fzX9IpZhO4Famf2LP
o0B2Za5aKXuka0Dx+l29OdrC94sGMNm0EXBthsVL7/fbXOKV12oky/eGEgUQvgYLEmn+oft/UuSn
SSqceNBaYw0uiCt2IICkMVJBEx+h5gozgitPbWJ4uXpl3SgAa83hrKx/rJeq7AgNZx71kiDXL/XF
Zdgp/rMY2UPDOmPIOsVQpX40P20Isepz8LtQa4b+7GRvGwMSPSGEldlJF7BFqg4mkoQOpHDFGTJf
spEDV/Ma8Q3IlRsb1mCxGzIE6IpOVpKSC8E1iNvKnvQaOYwN9kBJjzkyi+x513I3D4cIRX5/g+kh
EYg8s+8vaJqOKk8DtxWfM53ef7t1syR+/Y8g4kr3AKd4Jhb8lZc0asVVd8kwmil7M4q5P5cj0gtB
j43DofkvGM07pMyqlHvqiv0mDIiNFLQL78O3LWLE7hxv7MiSAOk0PiAI7dvO0XYxzT0Aw3NJn9Tm
Kimyc0CBUGOGHGqNRz9A0KAkfKo0Q6xyrYVZ+PvKKCFhiN6aiTQqktfJOkLqvCvw13bMXhyC4OHf
rBkNSPvJ/hB1RYn3Ngx1EvFYDDNuNoDSRS7M8HitPX7zTgNvS7Iyw+6BNevlHgUMQkLNiD0U6ZqC
VS4PLEm7y5hW+1Lz7r6x9GynGUm2Owce9qkujaRxyvTjsm7lCQghruDz53VdlwwgZCktTvzBUoQd
IM8LMQSE3gvWBZnylBtUkz1ZHe7I0DGcm40B4FfqkREfv1Ahj8qEcUXCQeAIoIsVQDoKmGzU5TRb
GMDJlVardDfvXadf7QFJcMtU4qlbBYgAl5+6E5M3EmGyOdcTrE9T1JdVnxeruXZGJ4/uiCcqYnCa
viG6nTH9KZGLXRBWr+If9XiAu2ck+S7DR59peHRQGIcapXwqhMmxmaDt6YYXl3EukMb8Z3SAXYcM
CaTU4FmQa+k2VfzLZBQKquTcRREm73D7uEvY3aKHCAepeSM0C+4+S9Sd9O7i30co0g0aSpLtLLKu
P3ej0hDR5s6cz0FM2ExbYg4Iwm8IZe8N6FOWHJwm/AKGu/I7IdN/D63+zt6uOtZmK9fkSkK8iEM2
GP1Sq08NSKEQ3rYux9Ho1koKQiyvMJbHKNIYP2MWMY9TDCie1eN4vEF0H+tZWoay4TA+6f5wQy9+
i6rsrvmZdyKfFASgsBUmKifQ4ciMDYh3TtGNn1lgVXVB1KE53boVGwAHFXKNgTcf3yfbrMG0Kp8j
LvVGdHiWNTQsW9gJca8CoTvS1GRGyDGdVVMXnK2Aqnsn2gbdqQJD0/7baDGwRcTfKbLxQZ2UZuJt
IMNfxpLQ18StjVr5CThV6RwspFhSWRUPOwXbrx725nmYeZZJdsRh7Nft70dx2DvMTxvVjoW9y1kE
bGCwxPDCCbM9NckRwAKw7lRm2T3tnhYkEJiPnW2Ud2fgD5qB+endwLjDUwiNu/IJzJXOpDTXXiZM
f9LpicotmDcyUxAXetGORDPlsfaxisJhuAToBqR+KqN/0J5GM4k1JNPjVOM0XH0WasbKPYGB1f1X
tHc5O5++fulqDzlsKpxrikUNUfc9BlqzhoiJx6lt+AR9DLxdfTRejcm0gWMm7j1BCHManrfuo3aL
0ooqTSlwKBDH1hQY1vvuXvQV89tiUwsJPbvNXkLAeDy8969kPmDeTdp3m434uNpb+ILwthQI5lyA
/hSahg/gR+DpU57yZkbT15E1+dzAWgtj98WuJhoknHwLSXYs9eHg+mokAiyUGvSXQL3RboHCTFkN
DmxHE/YjzuR9a61oEjeKXamRntJfjRB7VqW7fbXQt086QxfCQ9OTNaPNjlQs6nxc8l0vdzuNl2IL
0nwUe0h74sMTWJpEkEuK7ryqYeqhvb7QIvwSlc0D85G2Y/xr8KlIhsUW2sWzoCzona6iVrzMPdDu
2/gp1nxYqlWIxDUIY82G9hTkdt2jBEqAhVUajHSE24ZCRUUZb6J3kX7t2i4uBoUVfmKBNxIOL4QD
NzyV+FDn6FmmTHu7bssUr9RPnuGNSRhIYbzrl2CIpUE5ivwyHwSolXDtDAfYTR5XewW2jGyxnW9Q
fhhcSpUK2ei391C2pfDrYuQqzjntzu1MPzyB75TLMflzdJpkrU9eLEIlUUJ2cU8Bi3s+hRi7msem
hz5XQBj8u81tj5WtV7mfuaLRnmJ7J2HK8vNEaHCoFhDuDcRSdAae1IX1D0wZ3QSKk2+3V+vtDxHw
dEEcpOeRZzPQSPihHwnKi4NT3bmcriTjhHsoWudYjWDsckKs6lKGM2bW3rMQ2E1K9swfVwI5cw40
HagB5KxXmSUnT9OCa5VuE4dnl68iJYaU0Av45Pw8/Q3aiv7WWnEIjrREXPAupH4vtQxy/z4wQRhi
tkUpGgx/kIov9rtSOKoSRXr40MKgP4j0lfbiw8vw77qPTvJn2inlQoYIkQ6hFrPA+Fd5MINCeFDB
L44IU/a/ZkBJaR7HX17QnmNRhINC4lCTty/aDRZEJYaww3SV2FFgwCcgul/QP3EggpQVnWQVcCPy
N6NNM30zcvqc/ITSB5Ml7MC5Np2HlUrSAMyex8DTNu9f66ecEebSiB4nS5e3X7BHMQ179JgOllsR
WwP3+Wa8lFAQNOGX8fTRpqKQKqOW7zk9drl48s5UHi8vPVUHSmPG292jz5I0242qG8HfrWFpJzvw
EHeONMAsUMuLI1lB5lb3kGrtWfs/XXs9mD+v8xBYOQQCTPiRHROQ2jaz9hgW2nheEkWV4vEZN3yk
0kEpwHI7p8jD+ApvS2AwM3VsUPohh/DLSklS/zvD3C0O43OrnfyXpaa5pvsSc2NmXI+GKHZBLENo
1qGdWC/UWjX6Z9mCmt3pRX4p/Ct6dvhCuTJIg2LCW/4HdUwQ7/s1jOeazoTHmPuXB7Wy/pGJner9
earV16TJEFyz+eq33JKJvDbROPkUA8F+uvQGn2tQohpwjAOYX51ByWeWMp1j9pxTiEiwXQCBYlXN
rnOxP1FyxAgh8KIYRAdbkjrBr4MnsFVaS4HjcZPLxlhF3063E6xPM+dKpRQMXhEukHL32k0IviIv
92/+0rqRONvlusvQJF5d3vJYnzZN2id09LAZ6+yz5FpbFQt+jVFH8dMhT1j4BZ+DWh8d5x1Zdgxp
NoJUXSdRhVCeDvIFAIseRDwv59JJzbQn7z1Onvh/T6vzt9KClccI7IiwNjMmyWAdwj0v6DYkaA00
d954rdQK2M3gwiBY68/k2SDB5yWXAJjNAVItOOypl0tbdrVVx1BN7afW8xP1ChABwv1wqNrvJxEF
7MsfLr3CDjwp40jBfIa3Rzjv1D3wuJb+MIYtbEIHqH4gOcFFwjRk7LeCSa3/ORFAp6pUlBlSHV6w
+POAVCEfGy0pWHXLX66abzM7G2YED1k1yJ5IAtCxBYMDwzphkxog1DWyD5HfaSWrmwf3KAl1WHOY
1CJ8EWSOTu9XUf1st6icvBf8kvwR2opfX856OtUJ3IFpv7PBoYxUlafl+BZGjQ4dUdkIYvxS52YG
+5kaYQmvCJrC7wJrCZQ5ZTl2PQKyUtvzuh3C//Y5QnKbHkGjAouv4tWr/XopW+05846853J0AP3p
CFwQLC6uiJ9A7PxQUGGF83CovtlKQBfpFUpO8m/v0TFPZEXKGAadzOjN3C8PtO5Mw2aCZ2zL4/rS
MWlULi+mr+HfEQRPIc+Ypvrrp0F7kmhLOylx1iR9nFMXPJFT8Bzi0VskGNyZuIP1ERAW8HfKvPpG
odOw1t3UpupR83NBPgMsfxFEn4+/TzOrX/7volc3YK+O1IjUPq6SE825ltfbvhHhdPV/nLfn6A4W
odMnjtuK2YWaTAQcQAG+e0VvBA/+GP+EMUjTlYcF+u7oTtFCUU4E9K0Zw1gOmeguY9F2ZG+Cpzr8
pi9+XPwWL3TnM4lgRvQ1mURw03/q5fIaQ31VhRO79cXNVtLJq6a7SiWghFmdJza4Q4zxdijEpg/N
CNyiNFvNewo3Lo9bx2/4jzguAkItWtVMqCSpBscxQSWVLli/yp6BMHtFqWIVrl38Mybjgit8ghSx
U1AenHhV2Gve8r5vDV5TY4c08/cWOF68TeIqVAn4y8whofAmwQ1iHgic4LGw11nXQ6usPEaWTNQQ
5rESaqsgX6SjWCPqmU36qtL1Aan15uVX/PswbDtjdWakwI7AU3hystw18KoLlxaF64bcGYBg0+0w
doFpRL/z1r8o9DOkkO9TUTSuXV2hinQCDVLSjq8vicrx5vKR7seD8DjiW/6vEh5f1lLeywsscg7H
y8QApJtlLTEg7ZOtlT3if3YRNkndDADSn9r5OqL73EfZmhEKPZ73iPX7RZLn9GMq+FdOnfL54Vr/
aOdaqXb8I8zDNHirEcr43qWj4VAhxcemg/9CgCTZ5N4PivZZnKHr8LBW5xxso/XvTrnWxAVJs4cj
lEgiHxO/VjAB153GQiwXnZrnjMQW5+gkhATkeM19S/nb/gb5aautu5dAOkUXXfM9uMZSbGpO14/w
7IT168YHCnDfDRiDcSvX2Vn3Zs7VumP9ZwkVahnB2TiwhXEp9mhgwqWFxaRm7sFnWkhGHKLrGHn+
Rrm8RU7dberKi7M+Y17ax4vcZqsldV0UK4OtigGj8g7RsfCXqqduv4Upwyohsd2vI9lGHJh0pbYN
GPJ/vsBtIG0bhDYsPd/oelZHEfYzroIgfl8S58TluDnyhO9XxIZqAb2hOekpWy1HxspGYBwmYayn
dnqviVSQ+FdifLVwKpev5HxJtNjzOmQEGyRXCsa3FD2kYNFWUZqNMULUIi6j630JWiaFRwzxrd46
L2s95K2E2wvA42V69t+v2TI/+Yy9beg8H1GoPuXlUfe5rnd7MyPXNB0A0Z4b1nWayXvQXo62iCW7
VHEdIldBBUDzu6ckLuxiVojXjWDv3jQmm1eW6H60OArmhrgqwQkc8ymRE45kMCvRc23P8WSO8Z/P
hyE8ydqbF640SUc5bd0ZK6C+zuWc5eSVw8h4tWS1xNZn2TJByXVLxTfhP9wbWbFa1W3qHlGC+k5p
yGQWfx1lkDzG6NiXjuRF2Mtm0tnpdFE+PkmZmvApFQtEkhqUiaAcUsBoRWMZ/XTR+Bhby3u1WmK/
kIXMYlCg9FOwoVxp7lEyONoDKu63WQI9QfXn6Lzx4KSf5Gocc25tbPeLlUXrOnd+a1juYw61LeDL
lnfn2iE/iIu7P1Gi+U3lMuvquSO0EFx1zmhVwEOXOSDV/GjllOb5IwhN31k5AHRXXSAzyBwwLsf3
Kjqw2GYBwKtNvnUTam/ReX9oHp2C9f6JQvXmxjpRubsN3bsyxdSqUapl8m62whKe7S2t82BaVl1b
s/+immeW9hdHI/qg5TvXJlImlaMAfd3ripGxA1SOYV/kFkiye8PHgQluXWYZT9hwIlCAxcu6GFPq
JKy9sS/U32lxXnoiNcjFlx2UkfMIULoS9VxO+wyidxIPH8+ipL/Q4WnIb1IcM9CfaV3vSkJWjXNj
ZGGGCxn353H58n6dezHESiLq61XFLdb1rAxHzsKmz7KJwYP7Lt1FAFezsYgRU3oPlR85TKlQkvuY
zQBMNNIhJ5WdNX79jIsSj8UyrdWwlAbl6eZ1dLbDGTW/IKUVfosoX1tMktbtCERMIqLdukWNnFdn
KhFxQSIrKHribsIX5IbuWz/dlo8uceLph0b+K93D6mpanS9HXP54e3vYRYYdMLfl2j6Ob0FNPOKH
SRTrRir7HXtojgUgrULOfJSNBR7ASI7EA+Dt0f/1iVXEvuhHoe/5VtWnCHtXcIG9NHYomoRXy3nI
2HOv/vjoy/OFVL6zD4urveGEgZIMb7hcBfdvQhYDSYFqaYjWdAvFGx0qm3i1j5+5htl7nO0v2n/c
zi8aWcOjBk7prikM/bQdYdbdZeXgLNj4PCITNjB5a3HpyBOp/GS3luRzC/dfRXzhIsQrXqcjyauy
coCvhRi0jk3yp/St+QEodspAziISHpM7kngJKIM203/FKmrDAaocu+bSmBSqWWbuAu3VpM0ciA+H
SF/nJKnnZL/9voB95mUBoBg9/UoDlimkNzL9zijTDSKvyD5f2gI8uYBrwVbWEqP/5gdGTl7JWu0p
hjqzM2K6Wp2PJUs4TsVbckWnUfPjeSZKnrhogi6tMQOHGlPGNzCgOiwHVCt0KN+aoJyhjn64oVj+
6jOcufPCFTI8xX3wb7HsSfGihKiGZyaLpapwvsA30Qwe3NzCjEhj/HZleY0QTINpm2AfmLOZZyjm
YhL0djRaCeG1kp0EQCwOe8pgb6NTFKLz3DsC0lLEQZP8x4dl4ez9dTbJfHeB7MqpQklOT6hTHWlP
FR3duXTD6RW0iJfabP3mCnwF88LX+jJlZAkCWEthAl60/KRK7M1841MGNXwx7xaP9DiyWQcS6mg5
nn2rEehL2LIap67vYYve6LFY6P3Nwn70kYocNl19QUsrniDcFm6EIh3A50uAx7H40ziFy2eW4Jbx
Bko+v2L3HMnvsvl+2RC87tpLrON9+Il+tjRrFsfEI9//sJH4wNcpBDaWQ6sEHpQ9WN4a7FQmCp+w
SHjIryz3IL24bxHjIbeaotUZVy1rCFRf9Vk9zAWKuwUSnHCqLZXuu7s57J14RvjafiGq8lDKwgMl
G/+YEJLjKAL7UQLIrYo4yjGlI8cNsCfQJcTNAXFwO0lEAAsktz7L1kviZzRs/6c+ym8dH/DWD76j
VYpxQ6IAhjXw8Ou23qDiPcGU74tebGUoC/zCX9te/2W01gqG4SCAtVZE/Jsm3IThARNI7VqknLHh
7bkVsSiG68XplwNaG9LeYjGCK87QFWDzKvPUzVl9uX5gpPcf+BkxzOCQ1dLzZ/rX4z+OoySuwKwL
jBZHrC/CEy+2vOOXrXQftt6F9szcD6J+IlP4prcvixWYm+5xWWov1h8V1knPmkz99aECQI0D0Gx2
UhQ1BTGImBFAiLK+iHreU6TwrHdU3jVSRaJmcZJe3cMDLJIzwnVVAP0z7LPSiC/mm2p58DSZdssW
SjUH0H4eg26NE+p6txlgwPAV4XLKXppz0jdo5KQUlkU5GfLql30JM7lR1fTzrGzKpzALA5uV/hu+
HuHvb7fWz/jXkvAqAEGw0He8M/+2gpr5Hx8UGyB0LIBNVlhQWhEtgHN7qvRNfhV2vuaeJcWKcRNB
Cr7OFHuO5uudegiy3/z1IMybo4A+yI1INvZ1cVfdj/mLaSEl2zVc3OAluwddI/5IHinNWPmcR7tY
qqO2Uou8WL1ZpT/XEd6x0IHlDtFbhrKnnsPvg3vSllQv71SMxa/2Q9zfODU5HMBDkW1zYyNbzTWd
d5xAXP1K7dqBnx1UuGe9voq6KxcZZSAChGilh8sGOktmEoaiUXwq9cFzv0/J/RlZGVJYwBQ9pYK/
9wgnQNgVA4W+RMO8lp6joJZV0ke+yT5LK+5WGO2MnNQalmtgsTv1VTSPbM/PILr06QHpBGF4eSWm
MWUM6pmU8LNzBZMzeZaKA4diDxijL35EkV1HFOOKzhL2foqIJr0cmJrOT2Z6sMaDRBHpUr3z7cgD
D/xjcWjkgv1awS6ptBVVXrYjMrpBMX1ngFZM4pqBy+h0+kUUWgl04FEcA5aS0fS0MgT7l7iArqYN
F38jIM1HUBbuOKxlJQL6QczDdwpaC+ftg4kbGRCOEgzwoyLLzAUxlEkBBkN/hZHAn/oQ1tDbfkmR
aexR4XKvFr0UntALfWHBx1locroaUojXWnPXnBH3gGXfyUuXis2WiBCu5cvK1huDn1MLjtEGX5x3
E91QXOyx2dfzpNNYKYWa4i5Ut7Xm+iv9BjMOK+aLjpTg7d0ESG8GsuGueXwZdq+kCJIau1G2WvIv
HTTnR+yP26hGZPB+uA9yGZ6zUfjLxm6CuBQaEf90UMWL7MPZQYYhGZBpGooCSOxtXmu/kRfKHUwf
z4TKJzmSbulRQs07iH3ctBgokLLgl2AaYvaNZz0pBshG+SH7itf8CRl5KEfyV2z3ddDrRE8fJzQo
zs9FgiGecEziaiakeAjSh8muKxK419bLOC+0Zq+iA6IY2rqWjRFCO/auCP9emlhwfkDQbvg+eOwu
B/m7r2Z+2znzhAEKIx/zWlv1jNgC3orn6FWGZoF+GQMuOT9FTR/t9isIJ2JAXOthcYISW3omc9F+
Zij5VWM/wXq2ETuGwrIfbAHg/BC6tveoaNHChEYT/EcrmkxtB4jfF7hTA7ziUEOOyoFwMXmZbAfE
1GfDZpOgKWiCrTZ/02uB4LpMbx3XHy+T09pAk3+TekdrelY3vdtccnbuRBaVYc5SRTWkAdHl4rPz
m3r4Vp6w7O1N8ZnuTkjTKRE2YMYhAphrhYUYyThmZYFQwbHEystigjoMK4szfgvaQQEiEJBaIelQ
3kKuSF7JkPlbriLlYYMlI9cu7CFdFgQOmLAVfjYxMwXH0XmcjbQ94ERRgMOivxOLlOcXncB/Zafx
xZPpu6knsj3PI1SknvTIW2ktUFdMGVoNa37lQdi4M2TncQheK6ChTYBuV7og2KvGuLMaUaRR3SiV
5xYyqVBrrfulEho2Jk3YeqSr1oPlwk7a15GUQCHZq1L5ZyD6SVI2gJKevncCXaKRU6iJ9J2JImWi
rQz/HqtN5rNph5U3KQ10FbxtuDEE/2QMeTt7CUh/hUgIPj+RM7/V7aVIEZw32wBRwyH/XyWOCvAh
6cczYePPFYF5GNgZpkts3vX5IwWlnxqkyqA5DK2q/a7e5nJZ1tH08mPL/t30yV1awBxBlNPxmp9R
QleC9J/ulfQu5mCTjF66UnWXEuM/brxqsSADvBDaOGmIYnE9P+5N6J/eTQkWh975SuF2U8mrBzK4
EsNsVXS9OF0vmyCqEfc823n/TSerobMt5ZnE0eP1Nep33ezCUkUrTQhceZvqGWlWSnn4EBYdZLg4
4pbfN8rBoLK2Xz7yKtH7xFLaUmTY9VPRxhtuksal9MwOPaMvJQRiSSu5K5qILnNNGFwUfmvBUSzz
3GNL2NHCz6CbcWG4SoE+1lq6Gb3vf+CfLZ2oYwdkFh8Z9BCqzX0ylAM4kZf+I53O6wBpjGpU9Yvd
Mn3KWmFLsJRcEB/aKWV5PYDhr8uJMaUs3zGAQzpVNsj2m2Cm7tQ/S9IrQDMt7xie3PYsNcPOFHsu
APkS2GISsFiadccvvGY/aiGNPPaOpQDz5NWNI+BLHBekGDTcydB0v7DqRmteaNIyj8iJozxxi88w
BT9u49VuAFd7xnMNm559grJW/N3WoqoczsMpjdfXAZrDtKMmbOszp2pJOqs2o/+c1ef/CPcZ8x2G
JLXBtsG7yVcfMgrwu9FOq0gMNYjhV1qkHpM0PKVtxyPxnQ4/kkDOVgv+nyq4ebbgrOug7DIPWG0o
x3oWKBJ99WdCgOGgqrAEX6UJ8BxfBi65pPhdsh+TzAzxeaaa+Z8KXjdu8UlqRqPDEc4FciOmDX6o
AXGRXSxTupjHgV6c1QJMKgOUtVJzEc4eZivsLOlWWLxw7tN3Y11EedlkvDm6dTEow5T9FIHdx5fL
Za0RBmNoQ77K81uxLhlMWDeyHiv+vKn0041tKTkOtUqZ2VwOuUuzJpOrLcz6LpqFeD+D34qHLQnJ
MF10cTVMNHZPmzbmNbHOvG4p+fQ3YDIfV08d91Fr60kFfgCtxAyl5jf2AJDeERWQBj6pRWKLgmfh
PV1O7xVPw6QsKv3SiBpBRHC4mtth36s+zOY8lMKgdK63S/EJdRBNOMXENmdUnLDIY3xPz/ln5Pgh
M13blp23dpKWxOzTSCmNKGt0INeAAptF6qRUVYClXqHuOT0+rsYgVexIfJDdOcOSC7bOEApaZYj0
BI1x2EB5WxoQl3pa48oyiK8Hkb5vv4RPYmoUBnCgNMVsgjpWjbOyCHV43X1s+DHgaCdCVO1+3tot
L94JS1setuaQIOlXrYbeBpk2FfUmoPBS0L1qaqLEzp10hig2o/BNo6kXWx6ZArJdqUEgDOc6L5/C
G1D2Aa1Cn8hgTc3xXTG3mqCaQOh5SElb9Vq+J/6e6McpEBUXYgY6mK4fG2gTQPAZYJFseHmBR95r
IPXmK9aiSK6zOHVTF2yU7rqSpdtV5sgjXIhAkvIZ9l2Tpp1dLbAtJXZpdL7Yr3YuoRk7egB/prfR
aE2guKAMBfkvR31483DclwFsqLyITzLApxgkS0qtukl8Vpyj3PQLQc7VmxJAilyYSCh5YW6aN9eu
J4BPHJRFEwfPRX1DvxeKWXq94XtmpbjQdeWD7YBZZEnsptv2c7kBXKZTuVSzQ/NimI4i8lVQnDhj
4BqwHWSennw+kYka2+hC2oIcSdV0kxhKzi/J/kn5r3CZtLleNjNzbxMiBifpUosWmoPQz0KRpWKL
H4AUO5Ed8puymTKNl/8TkwJTx3upgWCTel0DWw4SDg/i1ERVeOZDA4Qip2+njlzHc90Z6Z1wTUi5
u2kmBdRUIcAl/JWGPedj4Mn6zLhR4ePBnttO25W7i3YzKIkPFqxgQJ7ghJZMue/Kqxxt1jUpYRxk
9QoCVlSJx7AySYE5d7Ml4Na/iGdV7pLqKNINGc37BpNwxfjmYVr9HO744XHsjaVtQ3svuLmb7Pat
aG93Ob2XOgnVkYadCKkRIkCOn4NcjwRLsCOVVSzi1Ka36ZvtykXKMcUx+2G8t5n3mloabo9gq4Ah
cB62ZCos+lBXgv7fhH3sbas1BW4xMkfGeG3kc5EUEH2u9kc1d+yEg9/XyrNPr2y3qXfl73Pp8YAA
wZ6MiX7M+S9U27P/sNjzxipj5jp/2G5YlugoTcXb2HBTlihGgAV02/WxRWISEZZFN1uosWqKQ1bN
o2B3xJNokbacFTkuRB2Z8AgRCvTzBaggxkU1LHypwR8QyxvCVgNHEMr5ehzBOkBHZp9Cmujbtswd
cbSGMezqzHDl21PHlRBOKRCDuhiZq7CdcQkuijZk8tXmAuGffEuk8hilPArxfaLPPuM6syUQbOiL
6u+BV92z59a4u0f7c4o9W0L0zVMdYmcfN42jtDSq4BjB5GuRm+VN3oM50GID06gAJi9PRgGXu1FA
B4KFK1xeHEha/2/M0qRjIF5vpTBo7dQRPilpctr+icVEy088HuDg6HI2g6pM0aZqlMoew5PtMGzF
deKFE7QBdgyJW++lwLLn22ksNPL7o2+UdELsVVRON+OAjhW2rKcrVb+b/F+IGKsTJssrb63f1Zec
DvVQnauYL3PbBso0tzXqVV4E4wXMkB/nJdaURwRPLJKYfsdnbxoXvA9QZoH3x1vbtzchk3coBPEX
jFhBJJnIDnO8ZwW9aj+yocF7UNEh9T+Bn+6JOhJnLedNJHiPiSHjFw93aPT4PzHWKgRjifT9HrtR
XtEZdF1UXF7xW8+JRYPLWfQBuNC3FkdI3B28B34PFNtf1VsXQ2dTwh50S+cpGiNBwEKTSWI9AWDA
1Wxj3njHSvL6n1763HRSdfoBJGprY3JyMhv9AboLwrRblR2rxMfM/PAzP0BSLHnk1hb5vjG67NWP
JZyeQKBcqu7bMTHcfSZ0hmo8H06rojGnyeW7u8uqoCzP5wrZJ8IiNVOsyjc3IH/ltDJo+Z7O294T
djMP041FH3EyheW8qBXX+vNpa9RdxDJE9uGoYz3O77S+hjjZ4WRYk+GYJYcOOGJbA2IEifeQe0kt
pkHROc6OIkmVNGs8LKe/0swtjywM1t6MxNvzh+OLlYKKzH+VUMaW/n23vBsj8bTeU6K67fXIwPx+
dSuSwJdPY51kC513+RPnB4kNe/D+d2MUkR7u4RAJJ1+x8vkKTY0s9bsoEUnZ4Ie+iBWzcUK7YLPS
T0HIBDHTO7ZI08Z3rUyJQM9rvBHoYeGzz30PU1t3+inbYWMKpZoIIdP0UOrYFVWJWDAwcvB76VMp
qMrO8o7vPQLV323XAPHTH1C3x8KjGBpc5FBIYnhbgAfpHWBiuJ4VuCpbkZ9T7QFjFgpPWvqqDGiZ
yTOexUgBFAYk3ArqKlTXPzKYd9w+IR6fT7/0d1cIuHrXgeE5m0VSpF2Fo4Ls+gjGBTJphO4mfxhT
fMHMswP3FItIgsVFtrYB0XydoSXJwBjyU8FJzsOS/3eVQ2lLxr9Tcx3GPTReMF4wQEy3caLS1M5l
z/kdZOb6cw8uUKuvaEKGZgkxBUdfKj6MhDOzp8ShxERhYsX0dAw82yFrIHobMmpz7c28VJttRBJF
KfxHpGqQ3AlRkcmJurcL3vCywPSUZgw5edgvBTz7SXyQXYu4eDpTKAfHA1u95KbFim+WMK6je4TC
bclqbyr+/6NZHLgU7z6v5cZSoCJjLMIIRwpEFUwSI2kiapGdNMTddfu4MDLJGfJGgfimQUSBwIec
9BmFxenkqr6x4NnF4Dg0nt0Sz9acDux+uanOCEEXLpnH6JmXbsmMsRtyc/KM1MvYeJ0PX152hVvp
tMqNdFrZJ6ET/BY0j5uATEClhIdWEl2XOYL2Hto3mfjajw8nKSdhzL4mHYdMsFZohQWILbPSIezB
wX+uyHav/XsPB6FwniZDRBn2NXYPUxN6Qux52kPFxhmE334IHgISuSIJw3uxAPHg6E3Oqoc0a06P
bIpIeeu5avnvyctVV+AioPqmfxEZWZHdpkWErnWlaIe2yprWAs5A89NqFuCVvkMc9s8SQAGBWxvm
RiKu4WoYdokV1dYW6C2d4HR0xDwGfMI1OCc+5KKsJQLRFmmMQFSIVJeh1W46pO3VE8MBF/SBdwvv
xMrHoYXbYDi+louGdiMlnEUOYSXvbcWSWjkJUIDM+4OO1pjjOk1QfE9RYkqUREgFXkZymtZTO9aP
tf6BJAB1ekCQABTeUowd6QT9xojCtwJ6lN0ZMgocvlHL+eWfVHAdXrcbBjSqEpikWiCCHx7RlLo1
6MTFtGALh0ks21A9c3R13s2BmuOMUM7nj/41Dfcu9mCIgjmyKv/x0dbrV9STXZUz+hMKhphIy3XP
n6Mao5GgyFoGFRCef09QNaeFAGh0lRBe9FV6wznURJdJpbRDVCTyBbGMliIL6H/KyR4S67depuGL
GaC1dJTijQ2Tf+Y34hhZcjt6lUVkyQsNJDe+6OHyCFsforeDe9M1NZWI7RZ8ilmb82WyyvNFWtyj
ROwpPIc5x+sz2x7OSmOpfYb2qKZR/IaDb6tKSR9fmsyc/tde6vWW7XKPyeFrONKjGllKA5Epnyh9
ISLvf0VhaREYSIBCYGFbAavhVofKe3EMTdFqJoYRgiQjy23QwfDN5X0FfkRqTsh9qi9klegxweQP
/Y8Tzait0nI08z1kOEzUCEy+652c0466HpWnxywQrDabnoxn3LRDJpuzcVhKnL1oJhQ/8lcPAxt4
zYqJAql+w9odRCJoFsVI7d/6HaHXHaCSY8nD6dmcFlH5yrjmXbqqBbo979OvyFTp6oqYLvGmiLJD
lcKUJavim74ardnNhQGy2TpZgJccPQxZ0NII+WhsahqKdKNLglI0pcxkaf5GGtQy2YkjFofIODcB
ZBtdRTUYKUbY/lsJcInXbIUlWVlQJcUsGX1XbKLNip2saftKJZo2BbPlqRie37CxJbkB7FouD8Fl
nnTE+M1wvpYiyq2nytc0x9Gu4BjDKt8aWHIPUHtwiGWEUksTMnBRCMnqCnV/RXVV3tnn62hGSk6s
zCmGdIw9LEvpYlw8NI/CEg+MMqI7apW01deMcVLRcWy0OQGKs1ZKtpMz18bdesNo8vePPYzfUSCf
w3gmLbaaR9oWlpQXRWLMhEflO9Vxjcl9xHSHyEbgkexndX87MTFFwuj6Mnvbqp89r9kzz9UhhQS1
dKMOSvUeiH4kirKiXPYiIRfmFwd8Qo5jEZjPcu8EeexWm0isLw2mbvb872nIkshvOY7unV3fDcB9
672XTjtFjDcUHc6h6LKEka0OAS/T71z5YISKHmpHbP+1IZVFlgkeUmof/azi5DRkG4gGDidbd1lg
TuRSTGDcYPYXek7OqfR0YacFsxKPsGYlc+9Xmm0uctdT0yepeZAtaEnO6DvwhQ3fVjGoVt0jIWwu
cXy6DYjP6YIIwRj4NlP1/+0SmYmPeBKfEkIekb5r6gNPMN2+5/RY+KlvM4xDRt1lU9epgG6cPEY/
fN7mYoSg6n20xJUuDT5J3ddZSHmZh0ztHgdJ5mxIw3QfF4ajJGR66EIWxyjyrgXRKFfOUi5kop4Y
2J6ARne25doBGIhWYz2KdHkJgAkCwJp1TSmh0yoqNXqsdDiN1TEDjgdFVEH/ghgvuTRJYEzRgqoa
bY2zR2cYQV9iLo+h2hG/Ho1qMV/XWnkd2UINRCsGQKu9mZmIWoaX+QV0gtl6s+LCEvxxjuj5C8XW
5J/Ky78YOED+7bqA8bhAQIAo+WgQcsIr8OO5Bh4W2gZfbhlmFd2kK3+t78c5+FqKPpBPqb5e1ofQ
L/lOisyRMeGEjfjZm8OvfafFGtzdOKUAqS2N9yJiQBeezqG8ww5BjUmUw/Wvi4jO2YCzeCuhF+3U
aSbq7l1qj4H9L+ohqVDn33i6qvsPsuW75/kUuYfPjG+mjGxJU7C2jAiIjZqaynasYLQJBzeXQNWO
58IxaFb9KSkkXriFwm7+6d0gSoOW3WGBLLsp9YJhE52vNbDSz7PwvEp6oTlYkJsmrTmi6mrr7j1d
cVwu5V/goSJvxbLQo2QNdO/3C3i7nIPHMHqePDRuFXr/QiCF7YUswvcpQVv7vd3KPAEK2LWMEwgL
5UZwnHBl3nkxLkDhP1JqrngNSRAIqfi50OFF0XKrC0fKJQXKxLsZJMbMx5QqcvFLnmuhc6nvgyq6
c7YEm8G7uVDf1yz1sSetehXmjqZMkWRla7fHIO61DujbCCLXnTaMCvIEOuyJbfXuYFPbFSTCLtaH
ZmxzXx2+v0cEHGF9bpaVQ29/F0WtMxvyq40D7wVHl5Mop8uHAbHJCocDPozwie3ajy4c2xRiuW2D
DJfniyhCDwwbr3y5soJ9Qxv3mWBeQRF1fE3fJruGIJuOqGkfY8xZ3IgASPHOCVN3uLIwioLV+PzO
cN3fPYJBa0jnEptlS0YLZwBO8aQ6pvArJLDJEBgjdTrx4tAzTJuekG3DEWj1kpfk67tJTsZ9UaDd
sCUXRKcTWt5pQA9awVPto9+ma8NGIRGBwJ5jdW9zxHH2wV7gCak5av3aMY7RcxdRpisSZ0ocM0rX
fhf06h1KfHsPyrz4GLt771mkE696aZ8Y/UYs3ripaYnevRx1Gr3TbH4CX+9/QX5HyVANoYYFRrGp
cldGEL6VIri/hWLIGv334jG0eta6WcsuUIrBFPfA8TYFMNtHkQNCs03Vwmk2fhGEAgGpRc5syP1Q
6i7F2cbTqO3Podn0I7J0mDD79xJsKG7zQtOUaxwav9eqYELz0T7XEB2MHxFpJ+UCLtE6ASRnSHIE
2NIP2V/cJ+Tlqt6HpC8vukKDJ0a7gJlu4wtMOv5M3/VRJFGzkgtYUCZ2nEqdd1vjT1/eitvdQGD9
3w2mZXRD8TCuzPXjQNiBmxSLPEK/5G4lsPG4ydcpC0+lXExlq2+oDUDgu4BeYsq55geS42xJVn1h
KGmeHf6EEq9jIOVDdmhWLBHrppKgl/fUAu72VFhOfY+ed6L8IOFLKPCKRlbDo4D9FzhmXPopBUEh
tPdcwn6Hs+BVFhojcNvNA64fdUiyDQpXpk91YoC/OQ17tUvmx/I7JD4GC9XinJoHtotJqWW/Babu
EyYff8HqjKmolxfR2p0p006aUMXXFsGp6t33I8GrzLs1aoNr04WnWv9ILl0z8E2vD4Me9DJGI0dD
1BvIUIrtF4J8yjslRgO6sek/pmz7zBr7vxMG94sp2KyWGQtc5EjqKI+Atq1XVvGCAEa1dCpzQSdN
ufCsfrSWfQ2FO2uRVyWNPeIt97aFSfhG9+XTcHd0NUVNqQe7/4zRt6Q40ppLk0OM4NEQsZa4t0YQ
0Clf0b8ZYHiul0vVGHlc2hI2/Jeqx1MsBcQn8nFm5RazxiUpJqHe0LEWciJANcJX1+qfxgrCvRHp
uuffYZZc7c+sBP1eO+YedprNAwX6s3aCSPRk1daao3hCZc0f7OmjnZw9aDmpgvWlaFgsit9Pg8rV
VcyeLuC+TAj6C+TektNEikPvUDusZrAwiLmIEGlS/ULceb11fbStzDR6H0QP/zV6btRdUoS1LyFR
kXxQb/3lxAxW3RZgbDSqRMVXy78raePO5DFzp6Fq95W5qmSXgDX1q/FD3wvL7OZTtM0rubCOw7Yr
bnvxK9DMhG6OMH4o4v/eERe61ZLPlgSBbD9NcAhtpzjV7suKMhjhPc12z5CYasR4ds5R2JarkB5V
+OoOJiUD04SKrw2IonatLkv8vlejfUEks9gat1PM3OARNC1XoHmHv8Z2IoP4/LqAorZ3Y/WcYzRF
gfHvZW6gp7Nn3nk7v2J1lc9syWGu8RpACrE1c3fgkK+MGBRaTRCDomRJDY6bdGUGOzjB3L08sU/v
YCkim2Hmze+ICdr4F1CLXUnDQ1kP52aYFvfTo3mU1jsvCD1EzyohV3/mf55Qa1cWLu2hNzpqLWHZ
TexyXVSlI9GaaSxOEcO5RJ3E4dl7xQmNKGQPQstThQkLnvbeb6LLOT/Oh8lP5f5uChlz/pb6j+/p
iw8uc/B5BNsGk7manZUL82J5TvUKCP1eWAi5UdkpM65lOUayu2c0ZUjmAfj9RuJ71LcnoQqFg4PY
MQQ0eVsTJodq/rKY8zLnrO3uUforMjow39+0H5jYIRD1TQVV9eaUC9q+2BjjAb3Q9pfCzjmhOsgZ
RVGhbvRq+y7cvo4tTF9xG85qlBIO5ZDS00a4hIO7jiKxJfQbR4NWdIoDIzimilBeOuvEDMphgx/A
j3uUTKeJyo4YIuXv1MzqOkxBAUdEX+8sJmczDen1KXgDehVMXaS4+CwVhBkgnXfholdtIK8XDELf
uq1N6YAYLSPDYYi+Py33AaOgbg4XpzOyPDeGJrUTRq0qeOIeaQ3m+xhz0iGhYg6exs3RecCrQALw
JAq11CcRcyozqIcwTYRccLftk0ezaWDoc80D7+MHm39BRdaLUkhoUN5h8OgKjkuMzhyveBRA8kOn
P8ca+0zKMbSErdQ4HwD3GMclNwQntGDMvlz88sIVfcw0SQ6DzlvXMIAhnSW1ZteMFnC7DGSDig1Y
QYhplHupZD4iYbGELreF5mUPR5LAImBRI1e9NSxUpcs5tY3RHMibKNgj/cPNpW25+YmB4rMjTGFp
2KcThiBmt3ASQEa0DMd+SMoXRad23jPiz9p54wjLw0w8mdz01/Cgdey9SK6Aurpy2DzdK4q7xzRv
aPcCVTYOuFT7JupZ5BVl1RCIDfVXlYbOh581bSBdUU9z7VnYQ1bS/OPs1hEaRT/pHrQdI9oni1Dc
+OF/xxJQirJnlw2rrL4xmZ77tNAtIqoc8WZSITbDXeaR/WTnoxqeEFm14EqDgs02UD/M711x4Mm4
a4LWEtlOKZ5XqvfPIiGluzht35ZgsPDySh6dgA1Dat9poknjBUOVBPjFFabzM24esHTDDl7cVzge
ljI+u4gHF77/0BkqRLoJ5z+R/LwHSTSeSfEpZfQ0E5pnm9TBTxP7L03k6ZiQwf+NmZc4derRZpSk
IHUQagyHjORkmzdro7W8rwwZ1ddpr2YObprZm8p2X2e7/WXJhyNnJmrfjo/QNw5w8rXiOYXWJc9c
aWuNIRTW3sIFDgquE+thLjEkYUqg3MsbWR41ssVYy4aTq5ayj0AX2CSj2sqg9eBC7oladggmC9YP
7Leiy9SGrZAr79t+hrkel6+Epf0jLisQIUyDwgK6sXiAJTKOJ+DEPkFO2QDHJYg/md8Xg3HX+Hs4
M+9xI3Gkzu+Ht6Ancwxnme4gB55q1IvUhpNjhOMhoLUJpGOmNpEf5+8JKc2fqAAlzHqvVvF04eDt
a/lzrgvYPoHOQwDQzZzbYvn/Q20s6Q7Au0uQuObgQAsJDY/lxvMbpkpgSp/N57NpH+sNpkyC1Faw
Gb9O+WBDtd+rezRVEcNsc0MDOzqK9AxRlqd0oT+0klJGZLh0YKORvGsaocPLZbfZq5t72lKhmI5Y
2XqIoVxyghE3
`pragma protect end_protected
