// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
goVbcZDDabC28JMJv79fOVrwl1ogYusi7ElgLnLEQp9/dNywLgduaQ2usDBly7zqgZjraOPuxCm4
xZnKqBmwuOEX8Wl9Ls10faZeMu064t33yzrnk3XEeg+oqbLeZ1fkvZmiqqvUIkz06UPuZ33I+rxY
NTfbNDcwZG3HyyGf76R9NNq/JbZMuHnlXPz+8w7x+vxswN9if9M94EwbD/5W9PBU4i+8TXZn5I3q
wHQYNy9FFKg77eil/4Z7rrnb11EbKqJ0L+3eMKi/DadBLDtUnO2DJIEA2Mah1/pOAwbGnnEMrurJ
KpfM+gr5CVk8aYV8IZpcPKGkSQSaVsnea2K61Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22832)
4U5vc3v6YurVqkNKi4WU07s+r5m0tkbaB5ytxahH4ZUCn3XGcJZF+rigMkCMSgmQngTOinC1dl4c
b4PtTf8MMfcxMn4E6hIRj1xxkPTce+CPcSUxgBhNHwRj5yu0TBl0zxLFgZyI2c4oDyFthF38CRd8
jBaPlHNLTW/juTAlgGa+N+fSJxFT8mmuLNw8NOlAPJySLO4OlvIWq5c4UlV34q+sS1sWmNO6T3WZ
6jrVfHrHT86dARMsQH8yNieMVKuOA7twGFnkI9LKCzNmm+eAHu4ZoH2hpuWirgDDsFtzjO0Q8faN
sVKXBdC/k7LxRjxGmt7D+wcNTfDVGYwCD+YIiVJ+uCekypz7E5dNxWbLPmS7AlhYCA5UN/6PYD+Q
qdnjJawblWhRzYS/U8yMLvRSENz0s48zu1KuiHhwsMKmBm+AXDfqTWSJTYnkBVFXY/FJtydMGomP
C0gcizJ3AhvzFlPLzbX/4cVDncwufTUVneg7ASanbmJ2EIdNHjtYXyhyDoLZjPFVUBaxA3ukwmJ+
VrnGmhnq8lJkPcqrA3qaWGxkNn1P3eNbrHYPg+vR+QGEIqlDWJ6MFSUSzXf9zI6Bsls0Wrw2dvXV
L4PbXKRmfEGKlXgdMvG+RJ4Po7blGjsNzNkcaIjGh4oYcN48YNm92NcP/lppVfLwnQvJNFkJUvaX
5juqhKD06mP+xeOtEV8g68dhcbPPwSCQNSW6662sabdzKFCrMhmUm6Y6c0sOh0PVA27Wu0PZHsMp
wtbY/6Ut1QIrUV3ndHsXXk6Q1BZJggIRHM4CMpJhqokZpww/lHk6/inRxIdxSGsceW01aTUwL0a8
4H/nrSIAF+xn2yh7ibbhqFct2KW+XBP491QE4WVqEME3Wda3aWs4pl8wEbkyRy+0nRCqAXUV/7L7
BL/9wUXzu22wiSCDzxB7pLEex/3dbouhnUC0X/T+myoiluJdvbDJm2fHnCcLyPMKp9E8ZdLbtwWw
TH7whfD5yDR+9cqnoeB+soiQJx0DxAhy57+PixfxCYrvKNLTdPce+NM7OsebytQKr+RmAg6KBNi4
SuXyOw8oPOc2e+WcRs0D1Tlodl6QcO3Hro23B8g/a3ZTRyrGqMtXw6GCoJZiTZsAvaDRuY1B6nVz
7GxsWbvVE96RQzhYYnEHbdkoskbel0GbzQwru1MrdD+n//Gg9oMpM0dzE9XIMdD4b9ZYrx1Azwcv
fdFWZc/7E1TdQBN8fQlLGZ1pwNEjv5PrinTNmVI7+pBYgRwGj1CBZMam6znZNH+Bh0sKyo/g8Bdh
rUm2L4O2TY+2egSBsUr0la1bTyMiMfTa1+dLlyUgYtUBTBfTjWecM4OXzVXLWRMbk3EsosHlP55u
4gmB/FcdTcfefQH8iaE8z0A3IK8gDuLeAHv3ctp5PBgR60Jfx+UZhbpEvmQf1O/1P9Ay5zwB2LLa
P4YW66fXA8GgttdqeGuFe+Agabdobk/Fe4+WVfj1Vcxlgk9KgcznbVlK+kEBg8UHKzyePomnax/I
+WmCn1jeF0G0vmkgGz1Ny0QBiJY3TwbAqsi8Ur97l7NeMkxZZA0fqHj6/jv//UarNEI0ZanKU5CO
JAhwKKeDK1Hs5J1wQilO/5kqGkqfzix1G9oeO1qRn2h64IOSf5v1hTbGPhGhWVfh3tVhJYrM02FE
LElghx+Ev0CleCXkiyiJjqpJ+HElnAepfAt1g7zFNrrF4tZqcFcSjReGye1GJPL3BaRdTlQwNAPq
3kIT8lt5Y8tt0wurgQE+lcQ4132q9eSJBJ3rZx7yVCD+AguMCUt3eEK72i/bw7EA2hShHDZ4a0d0
GMxbwxQVIO5fM7X3O26/hTEOKDyXEBGOKvv76hfsRmOcT6xBvUZXHEScJNmX0yBm6L50Lmg74tP2
2V5yrBfjO2twgms77avGpfVbUnudd8HLsGLR1o/jaSkHT6aZjcneoFFp6UR5VU6a0PsaR8RCUgTX
PvLXc9uDwsU91X3mEs8QkbmSaiRymlK5J3gRKAAV71zr56Ktu4fe4d2w6EMqQK6/u/5w1OLmoe1x
nj1e4IGCleo3Mt80J7L3zVj9VbCFoaiTSFwYtW7CWPWfiHUZxEuUcB2/bHUQOsW5iTYQ5CEvljUM
PnGrSeGNvU+rEoAfuMx10lGubfdbN1YaEkc2CFQVeeP9Y6GINpFh1FPg2ytCTAhbpTYb7jsFiVTm
ShTFvn7HwwQHg7WbdptSM66leIs4K5LK9YOk+NREz+ymZBeAKoY+E6UKZqDQ5gz8ZoQ9yQaH3HBW
FJ5HGeVRTadd83rWjhm17ek0AZoSUQ1jiM0oEA8JnchrkAbnP1j30urUaZXZZZ7FK8/YD5HPJVAh
ybM5NPDP4l5TM6wZyAbzr/FB9rUC3BQ9ZUxuQ0kVFCMUukGg2iAf5dg9roLDY5TOAm1snYSmAm6J
dsJHJrhwJv9FIq0USsfrv0IuO4ZHreSjlFbq/K1czWR6k37mke8xfzrfU9viCNBFfWK0Vj2990Vp
wROqC9iJLhSHqw57C2B5m58CKL+YmJQd/Ox3uqWS0074oTLZqs8q7kj6wVVVj0zmZqX/wCYOrNpS
Ix8uKDmQaCKIs38D4xKYn86trgUYo5vvVPg+L1Nl9ggrwLupxdKJ2sc/oUbxYh8sKnS8BK8l4Qvv
AcqrxVybxq/c2lP+VQnWocQsDQmsYi1EesZpBm3n/RIulF9jMqH5Ux3OCmW6vdaNYNqnHWKEe86T
N+c9P3BP+YmlpmCXVyvtkj/6by+vI6FxKEEYCg+GzYMSGavFeyVm678FncV3L2Sg4za4trwoLU2u
STnn05PU11tWs9IKdmeEzoyC9O8eTAdfzjOY80foNrmgwaLrUmdlOvBmHlkehGkRhXlgUeafEoeY
s+LCaZHDj+nm6ZelF6e0+VERvP1YmYn/3Z7AOfnmT41REUgk6xT4S4Ew0cVjBo58Gd2wovXr609a
kNfSgO/PW/5hYxuRSeo480c+KyoqtS4oTGPd/BvzwEV933aXfAjOxHkHrTF1jZ6fDpMQLyXtPnq4
L1nff8a3b76INhG5Rt50mjBLOPa6JDzEwycK/AiyypN9rX3BzjNs1cgK1w2gWFO1pHILasOsF/Op
0TuhxUJZ1xUyA08qTNvjwcECANDzBbVZY7t35lUaXd3f0bLhuaUwrBAaypWY6fJ9Nd7o9/XzVGUz
dHaGVsJgydmiEdvluvakKIQwzuruiRACUA4PyQ9yMeUsXMjpZ3iJ1JkbFRy0yuDteH8ba/yexXzX
MJy8XNw0conOw4lZR4RS1wizu8+JHTG6mC0rOH9YN9imQ/DiWobtQqucfMfpEVDJtnxnde3Kbt29
tb55kRa34/g9XXZ459s0C1kTwjqKzXCf2cTSHM1sXOpaBHMszfeULPjUVOitRrLWoXeBo0iPZRU/
L/dkdEocmX/eWVuhQvQicquGqbL66RL25FfdWTnCrVhznTnvZqdvbBdUt5eJT2J1nr+JHSctfz/v
dtouVND4i+Y/J+z7O9s5s+7ePXwnT1Dn0ge689/1NdIfUn15hNhmYbB4qznZy+tRJO8T1wNL0Bge
e7AJMlW+ihxSBQXztU2Gf4rT76DnTq3CBXesR+oQtLG+ucoPDL6lPAy63VYhB2wY8al3rn7EBF9v
gkjJ/84O+oxDfN1+cFrSAnxRRpIcn/FuFjcT2I1LZLjDHk1AXHKQ7a/jJkIj1/7WbZhGHx9owPFw
ev571fVomaXtaUrDFPWftTsQULJIlptZK1dvM30ZnkxRMH5cmhZ//XfDGDEW8sxUVCBXmwtL6+Fx
TKq2ScebNI5JIauGJ98qPapIkRT1Z7IsafAqLSEH/rTlYwrD2VvJV1z7n/vc8o0FfWo6I2yO/v9e
689jPcKJv3S04GA15j6G8XF8ilqVNsWq1CmMvgAYgH7HgfXt25gU4MFDs1MDCieEnAw36oMiHW08
gz//aUv0W2DJwRGEWNkWtDawfLzfFEPNnsKvc6Ym5vy10hB9kWX6ZTCUu8dVGfMpMvyHbICZa5Wj
JqmF1mtJEIQ01ePpIYOZAMD37gl6b6BMZIx7p7jZx8ul2D+lFAVXISqtr6wEhGkJ4IzI6IR7dldT
E/J1/H2EjzntA0QkPagJvidJZNb0Kusn234vd85mpMzz59Fw1lU0SrRjegRni7zpZxCZfRZ33O2v
CcJGwiqs7b1bP67MtxvhZ/IqKh83zRza0e2F1lZf/fzR3YBWP5C1go5RYKnUoXv/Er65oxOXN0Qm
SNfT4xCMVtXLZprjlpPiQX8MRI5azgJIm3+6PXBBw4Y556hPK3+f2XBaLCoK7U5S2XtbOqqRBMIR
5s9BDjGNdmK9qmTexYAHhyYxqwEyu2zQqB0+Q/iP2IXRxOt7g5GIbTkLaOUpGX2K6uk6/s0dDKVQ
/E/KY/nOwLCeJxnfkADI/+dEo4eBXR3yH3ZGWORcZtsLgHjJPynxCNweTkfa9WH1ID2Akx9/g/HJ
hgD2DNezrmcMeWmAZCdictJhI6NYvvqBfcZM/u21R2M5+aAHCmM+3oGNq9OFKzsiWrf6/mJuXh1Y
94MTmXflrOeKe/f5tDR2EpxVrRt1GfspVP2yrY3hWWe5BwGp4vGutecmILIhQ85RNw1LKODa1Voi
HEAkoRO5Xmm02pz9gGclEjZkhp/SLdnGpy96lHyBYSV/HDkVZhnFVVvKAriojPeIYvQqiZQtrgtA
NCH8GcJg+0ClO/1kL2/qbFjU/pQ9ifLc3pqKFQl3cDTojyMZchKx/kCoOqBgqloujCUsOqn7ORgd
whaYSDEwVxcR8gS7nz1NODwp0FzimcNiEomZZfnU8oVfdxoxFgaK7O6fmlGsoWQmQCVtFj9kwbyI
N0+CsEHXOdYSz+Jzn9fDmuu6as9FsDIcgn9uwUbAYU7YJ926gtzU4Q+uTSEcIxsm/rbn2RQBy1zN
vG1f62Wg5QKypfQoSSKh4cP47DY6Ft5g98Zs4TVI6AmMjeKgV10dbdD1BK8GVZh2KNlAPX0kLI/F
WKQ1R3h/TfxbFZPK8sORCaBLMyxvmN91ejOXi/GIBvU8G043KufdmVU6VLNoNW7DZ2eGwgW9/6c5
AZoj26aPrvEoqVk0u2uwTiq8S4isuX7k71D51GJczKX4cGBX4GeSQHo1BKhXGavaCeLLsC5W0z1P
jEQjhTD3OMiL26fQzXOMS381jjwuDsNpXkZCDtditKKWUrM/KM8JVDrDk+9CHIAI66VWL7CEAzPe
LXktUiRNyvU6mz6n9N00uuVA50FtF8Sdlhzd0RLahH9WL9mT9erTbrG2vYR5Lav7/BSc1IRoEdSZ
BQzdRoGgy9WgPti8NHfnaFWtUYNAcu1M/HbY1mxr9jc0pDz4ch1CuFPiP4USez665O35M/VS3EfX
HaK4woGGEVa3OL3Z7Of65yQ+q9w9uH71h5NhZGZBl4ymJvdLhpmlf9IVcTf24AoPbS7eqmh1DrAJ
xzuKq4utPktak/Ad10liTHQdFOnv/8WFqi1phZWdwe3woitZqphFuSTXpTdiiX8bA+g5zYlby4NW
O0GWKEpyBhfUXsSRtCOIEVGni3+o/zGae9d6I5tupZBY/HriudPp+gNMtN4HzkqlCNJcFGcis0ih
QRn+NqM8mt+aB8PqMDvZ+TSMtrI8L3sbfYYdn8ifwwvcIqP5JtUh6RPwC4QJxIn+iFPYRP+24xwK
fxZIYYr3F3da6T1FOyUbwoUd0wFD+POpCpQG323x4uoXIq+yN5lPMMflQDdholZ9wkX2I945VcL+
lKPA4O2I9QwOCDWiA+8GRmmvrrX2etlJnExrngVWHSL6CDByw7Bg07KWFQBKGtrOEz0M8qHxotgN
iAvm1ViUKjgFO28HIbuR0Hy3PZLHW1DkTEc9D7iZ9X71lHOZdfY4Zm6U1lEvVEmHLXNt6/Cu4L/k
aZ/IFpYZWCBzzLkLGv4xfCNrVppRvZQsn2n0bnBdHvevSzMRUgoD/kkJb8WCayZrUGa4e3cgH+EK
ubE6UEeU1ASI7pXGuPaydYFaaPs8diYbKA4G3Dm7XywujK73FlXPT7hxCOocdetypfSllVowTCAK
HemwItcwUm5hnvtUQqmlq2OmszPHH0RQDQL4UCwgm+51QY6JJFFgsUZP7WL2/Oo/E0r5w6RxYQSx
k/ckIRmAi8yr5Ike5CroHVZK9DW2+++VejhqQdum2p3d6wNL8WckSe+3QROzZu7ngpgNj1sTylN3
44us4ZCDE0LZGFB36+5NeHykwx4Nn8po6+kwNdUCisJUrnz9Sw2pwqdqddToTdDsC0Zia1Dte7/3
7wmOina9aNHJux8kHIvr0+t5ThVLPIS3w9YWJVuKFzwpW2IsnC3ksbiTEhdSZfaFwzMaLwySSZEb
vEJ/gVc8xvZDp3b8kickm/qkSiDzQLFUIMkqw1yvP93KUtl8kdY5zoHRi4q5UdNb5pBNNIbRUmKd
dkNg03bsATqL1ZBqDP/6IqKPoL+o9py5qay3JNqCeEK2nBwqwWQNiV04r9MXIuRFr8pmRREUcQV2
ZRQW7pTBsQz0c//k3Gv1ztvg82c78CrFU6BI+51q7Ljfuj+cKZlmxzuCZJIDIyhhatKWw6s7K3yW
NnQ27X7ZMgZ9ykQoiS0z8BioVS9AQtRQvJyblx4zNBxmJ6qLBoNQsdbKhKzFbusQJpc3LnxXtqFd
F2NnKNHv4vghBBwGXNRg8zdYtHDZR1j/UbbSNufdWk/HL6w8RsU8AZESjavnHwZVKQ9x75Favb/4
8ffJhvY5OvwFhU7m03Gd/iIaVx5SDYgB5n86TZ2mli37Isq5PVTOq92wdf/4yoidjVoVF6CK+/OR
tirlUMtT4li0/Xh3H/VJuNy4lzr1W16sAVel39/Nibkwi43Z+uAX83hrh10iFwn6H/KcHIIlRhnA
xGdVa2YQ2zbz2TbyEv0zcG4H8g43ak65SBmNVtHsnuYlghYWM8mvRGlVBiynv1OFpWUIu8Drs6cQ
nL8XSueH+T9RgIRjEfKNZbLanwTFWfIEPdmhUGmDq8aG9orAJiJerWbCY8uS4p9IyavVHgIUA0jT
3l6OsDCnQD9kz43kKi62J6L750wGTXbhtbRznGhokdxgLQwVucoVAiQiAvG0FDvVSDQYwFZxfgMI
6ob9odaDglKbM1AQCsYxyp5IARIefqtChmsoCaC+BQBuOv+ovPpKVLrxZneF2Kq4TTWID8HZ38BD
jwkW61DthSDq834IiTgxjXTBlcYOvSDwACG3f65Wbya1lm2DniiPCrtF/r0ijCYOQQTQLw23zPz4
y5zwpvBl4GHyKJo5OKrDwBGYAAbldoJRse/uFFh6abnztafIbBYhSFjcraKQ38s5H3dQiBRRM6SQ
2V0JotM8nCnoavRMG1ICVikV3nCljIpITqDjJUwFdV16VUJQ87SqeDI82TUrBICkP1velnEjaKnA
bsshVgSqYvo3GWclKk2uSbrB/a0pqBhtVkTPxnv2RrxuMNFtGsgqsWwTmSYpFWKeXsAUFLdQoGHN
7S8IuKV85BBXysaEZkxxcdU7rY+RP3+Spw3+wQ3E/29DCu7VhVSnm2OXiuOnpk3+PyPtgr57bWk4
NpSA8pcYGRMTXZQ9o3/lC69Tlrv2wL4Or58VN+yZ0FqBtoYcJYW4RucPkFTamnZnnVZMIfgfuoqe
OAEDukTBPf06NndhgvE1YiP8wqLwEC4tHL8kLcER2DJhXe6Dp/MfJ/ZeTaAhtwkiQliqUjBvu4tk
wnmhi4eS2Hkn5HDKh8hzRcOXd18IOfgqNbl3hD10qs2CQ9EMbNv+dLDixMXbLhbRCLHDr6hKlM+G
uBLqNweUMLki1xe7fOHDpdJKlyxxphAGJUkXYAwht8FHCGdS4Wfvj7nDmhVNtZqBwvZeizzSHeui
TrbmgnPmwm6hNTqQRSL39w4p9mh1G4HmzGJlsk2Ktq3HURhq2Y6v6KPe3W2Wn4g4RI/xmbnaFe+M
IaNEOuwPcjTFxt4T0mqKPM2Hi1XEagaNz9kkmyfR+GB75sNfj3DGJiUsbvZ9pNkX4SrJ5Tzi/jAh
mmG1wjllRQbO6VX2NQoP9iLzq57nIJKVr4DK2X7U2ZY7NHbiCpfpLnNvBW68DMHldJPzTo4eB1dh
+UWno3zrGyS9PCZveSkdBzFIuGyLv1xQnCje2QDvExI9yuhGEmuc1E/YkeQZiId36ketC/Ge9ct3
+kzMurwScqye5ErEzLm2g1+EIQ7VhLB8IWH+EahraP/9gWXySR3DeSLpSUdqXaD9Yuwayeu4qKgD
00BKCRsY9KS+w+mMwt8tHbVdrKlyvTKmKMD2jhOlRqBKXmvgFs7fxr4U+kWe3gZb/kUzAD4YDBn9
jZj3NuXxf9NqR03mvEQIxepcXaOpQXtgQWhbpsFPMdVq8hYCVIavfK8UKAH/M+zjZn1DP6HrmpHI
BWSDXmrQLBGsNv5sszJnmS94nUpnungNHewrTIQzkPZt1u0EGuP9pJcGUWu9cbIMfnUpdp2ckt1r
aCiG8B1PAlEIkxhUkeeh5gAnR/MPKknUtNdeUjreakj4Vc5gax9LhUQM+Z9mxCf+VLF9IQps1g6V
HsckX7AzLZj8cWQuQicp18LRiJlFGqGACsHcitzOubJjYVoduE6CLAkjkuVHIxIYMworJP3IDBP9
L5XbDQWKHh6v/ivEstPp/GU9FyPVoRaP7U+hn9+gioVnASZegrqVMI//1k7VMaQ7yh1uy4i6KAWj
MaVNC6jzTsHA2bhtxdpS/dlm7ig3NmocxWYH7KEH26k62rDOIBneZFmNfTlkRC/1YXj3N2xKesmP
TF3NXYOFu+dDF/U1kFykD/72x2Gm2yqAY581BuB2S+nG2xMuZergv9EmPT1ya5M/oTr+JAtkigq6
K1iSQravp+IiuBnhhNz7nQaW7Y9sLLnfa3xZhvfUVkmZ7TjEVRGibMvphWF5H1uyGv6eovr++Tdq
LPpAOexeQNOeOCqiEq6cSI9fkzvsdOHKB/drMZRZs4H/Rr0RSGsO64EcsCCdyp1zMySKpOvgV+G6
XgNfKC+v4iS9zSKie4FJchd5zuCBng5xeZLDSHPqj8EOOfkw5McmSnPrxRzjxt3aNFypwjH0toE/
bvCcgngsLEIs5yI72gwJNfqA3lv4MobFu4ugg633k//a1EbUFd6YqZ/aVDjcDO8nK4vjptYzYo7d
as7hkiemK9BU9Y0Y4X6C8OpGFEAiv3/Szr5LFZj+oV6BxAHDJh4/TcIlE57eZGCy+ofl/lR+K0re
3JJLPwD2Dfa+cDXVFabdsIqcNnvVMKjysJIJtntJusnpfgzM50vTsw2Ap5f5bNvxQl87fuMkYm7E
ZJTQlK5XewCjKoLUVgUc3oY84pYkc/E4B3rkKeVBSzsShQVobRMuo/bVs63pvQCD6gZhiNDxWKEM
txsjVBty6JZVkTqERX8Z9f3T2echKppxhTCzB/g1jI1xmrIpF/MgLYojNLiQJ2y+A423Dp/OTtwx
BLJSN4MCJaazCe6er0FWYm/kVrYyvDOw0GES+rZl3/XBJFtIuscyjdaDijZy39sOUnQzXI5VRG6T
mfIx9UMS7xPCiR8EadyKsfxiBI4MYX3Ab+9rGIImOJGXSebhlscoMjFlAtFUlWjkkmLLQIvtddP1
ByiYNSCTwStL0NehZGkigvpNwZE7eA+ESLHgk0miafeyuTGXrODIs9MyacGmV7TckmksmjM3DNJF
S/r7lLrGvtJoyyhtAxiWDlwgoApgFLCwhv6+GytUkoTotmagw7+j3YAhH6XpDtlxEm/18kC46eCx
rmFgsT+cev0QJw4Lz/xgWCGy77dfLzzW86s/qFO36UUuOOBVjY5IxnN4WpDqSELSeQbjp1B37hqX
fPuUM5JnTFA5pfl0pRk5EWgxm/072OlMc6o9mAoRv34whN+WoDomTA9oN8dZlONmfu4CImG9yifI
i+154GlsICsqojQAywjqIiXqrgj/r8DytNOztGyMz03fmi8WkSyojdFs4TrXMybFvySb4buMphhL
noAhznwysXDkBMXZJ11NZG32ULsXYYAmCsyLK8WG6+bqMwWcMh32poPCRhQaz0b5pVSbipxOfK5W
89VAPuQR6g+1sBVDeRDuaglCVZiRWTcw549/dd/pEH7gA4yDUgfWdPzWfjpwPIL5mzgM7iudQZ18
3vW3wTzCc0ajy3nbptk5+iMOD/IoLJB8cSKLPIpnDjTM/omshcsz1g/XrDlpxyIfF8qDaQsW9WTI
vnwHUPTvwiWdyyUf2YHDRovMvRKhMSclTkbE8L5YCnm3NFkOToAzi2CroRqtFYE0RlFBwDioW57w
wYT0ZGREj5NWIhqMFbDN8TN8aKRLPMRkvW140PHllHZm25oWScST56Xj5sIm96Uofs+nbk3BnvSG
RzLnysHjuAHqCMsqVrs/IBPrKoGKsZ0g0wW1noz699hho1JofJqysm9sTkbMQWZk9KFGfSK+1HGd
lrYug3W1sDkKrdCSYgLks1A66d1tCdbIpTqcliJz7D6B++awZy0OAF3myJrs5lES5TWGWmCRsblf
wQ16MDhEhBb/THWwL3T7VY/W0+KmmjFYacRe7+q1Yc0ZsSd1baHTMwTb6970UHqMD0sniw+vs+lE
5MiBCpuLppOpPEpnfhxdjEyM2fjDsAW96TRiwHPE7qF7HZiUMl78c6L7hho5yM6wnI5SjoAF+w94
BSs9HSGOOZbgos5Wo6nXQtH1XkPitpywGuI+wzbarR23sJ2i8gEBwydefkRanZWNeQe6ctPIULb+
w9Oky4cfPof0+DM/X7Dh7KHR/HWs7hCyD+Ja10Pawpc3XHwUeUFgVErl/htJ2MQMTz3niImB3PO4
WcZ6v339s5NAXGI/8FI2j1sI8DVDTLo7J9LY4YqwVkD24GiX0a80GU7KSnoO5WyWICj1TPMO1ZjN
79gjNTRjhjgaEVHlikj44AQm8nCevk/11O7aBqT31VwMtSrke147aGfBxiZZ8Mcms6AvjYVatYHZ
29uEvVf3jgRLkprBI048PUDOnEHwHGZa20dj2NfbvmdngOOJn8nXjjy2eZUqYYAhXeArCYHfvFR5
DCF9KAkpbqMsHqsN/3v7leFp/BqAw5h3RfNeFizVa2Hf3ja9BCeHWyhhkckyJfpP+E7ogllfixeF
8mUl3eoVVcK9PBRiK45yxHiQG+mlTU3yZ6aHAUqxfRat8Dz+UdNr1HSpC4aO27t/qGQIkCVYRNdI
r4/p/y8gtjXCzSQDRa8ohxY/SHWayPkSrk1oHPG3GmOTTjTBlFu6cV72zK7WXz9aOPms5MN6J3u8
jQ9UjQett97yFZBtsrZUo5lU9bLNDD+y6V19UtHJodjElmEE+5zHMOsz+xUkKi8TM11Qt4GbE4NS
RWXzzA74Gg6ljHKnmcboIeY2V9XnhyY4ScC7hvBNCs4GIto1ZRmGih/BHkxTIa3Qr8tpyJJgPWnD
6A97q/faDAgcWdu22J8lw7iQ2J5XWFg4QdBLF39RvxE/PWFzyW6kxRrLYavzavX5LyUbzsixaCfO
mVMB/KeuGnsl8cHwx8UYLootbeCDk1TxH5ObYgDsGCJtYX/0strx/I6/jb6cDjmL358wHuK6w0kp
4BuOvRjGxYfSBh0k3se0fIC64i/8L1D/jHg077DZlxi5xi4eaI0Wu7/7HnVpPgcfAUCOEU7V7SpZ
/SbjNtJFCquZCK3pQruc+KyeVRZDN+WUV72TLOfrKeE4Xo/bpNNPu7oeKVnhogzcwOtjm2WSS0yy
IVczt77cvlXBXxAO0NFuKf5lmEqrtPQ+VpW4dLHrFYdZKrTEXzQFsO/nO/EmVR5RhST2LbPVlWzV
HlpEkGbREyNbJQ76lLOAHVu+7G6Hu6WgFQ6aTJLw7z4zu2YQoHD9rqRae0i5qIGN1pnFMoG4bb0q
N642t7JyQHxwM18zgl8nC3kwFnUiS11atMZGGmAdsnQpXPPjaaypIatVlyttdyzV+g8A8F1OPkVc
7r4pzAohUp6uXsXrvmsGGohIeYqBUwwVvGHGORWD9UxYEa2dz/2Cp+cGgRVisQf7ggWA64+SBgd0
TM3AJ57FNJUKFlIMQcQ1tLAsjI74XDP7g0CwG6zpTrqIYgv/bXRkbCArLgYugXXrbZwlARy6ELEs
arGdUedJQ85n8vA9zH6iLBGR2RTTje+nZq+3j2sWYAC1JZQzJs18hKKQymRR04PJEr1gQC5wv/32
TAj3L/kT0UuUYI4x2+G3T0HF6fwgES7ZCikpdmrNCre4QBNP4+ZUW0mlVPdd1Mo9K90tGP4cFgEB
pmN2RDzps+UebUS04Qv1wuTBx3LfU+D8bt1LvRx4wzFWWlRYVTzXoxXz1OLjYJiIkmKq7T+42QAt
1loWgUXdEYzF6Cnr/e17qp8HHjh/z8y9ZMe4P9ppJMc3yNtRqv5OnCMnHCMh9uU/7UrxOiZwrsu7
/7XbAGp1P/qhmCPlIBGDmljrH73CSy2RFADJm+g1xcVFS4JlBipeFp9SMdj2TAhmH04WWhaPw9gv
Foqny7fF7IREaGtxzcZ390lQssoeqdNGrq2BqpB2CgSoU8Xc/FDsfsz+89VxK+9OdSva+xZyfq9K
1+/i123Oyao6UJSCH/wwITKJzSYoAQB+5FurHHD/KEV50RHY7aiop49b97dv7XJ9BirxDiLAKHMd
U9YeE5koaABxAVKuyhua1rSVdu/pZnNJ/MNZNH8/VFcXNI78CkBM6MIhBbkQywGp4ON/R9bLyuI0
rFDnSbByV5WkpAgvJQP09YkmybBW1wkjrFOLyJfenpWIDb9YapGDbP+c2hY9+jX+3Pn+3xY9PINR
brQw4a6Jqr5izCNRpDNA4LuhCmmcHUXeJQ6K+apN+tzs11RBoGMssw+K6sLoh8/oO7hX2Xv8x7b3
+5Vis/WD1dI0RE94Iu7GRslFqjqsv+5R27yYNAdV9TvM7ixl0jN+VvXVZtcjdr32MPhbKVY98Kmh
jDVZ5NCxdC3qO43ei+I+t1E/t4aejf7ZXGcXrboSrSmEh664/FLaf1KJ2gaxLnhav95bC9Y4Ew2S
dXBaH1GEON++aBlZrboorjClBKtRHooK+xmSbWled5675LZblceiIWcWznWa0okwmydf2B+QbdNZ
z42wGM0cOw+KiZIbFxZq3XqFDy4vo5jS/tS7/Jjy88Qsv3Q+KHn1Jioft7k4K3ygynhap2wTsLhf
Esw/TsR4OuUHLIYICMJSwuvnULVE/nW8pxfdoVpM1KRhtKpXFjrlyLRrckgXzTzhG/UmazVIe7lZ
kHdCVvZd1guYNrpJnbTb2Nz5F4lPffDFrYwTSnHwiRhhAkB/xVP4NtfZmLq2GDmI9jYXngejkwHF
z/eShSIeJXjy1h97j29rninpitWjZoVy4eQTbOlJSMcPw+qX4J4qy+iyS9BdkmQN7AIp4jNzbeXo
DD8JVknAxAPfAHymAgWQQTrDzST9kuLFnBcKFA2UJ4a0E5tmdw+5Ti20iYDM1mi23xA/7oO9lCzk
QVH0DcQOApjerYq0PKKLiVGNhZMxkYklbe81emGdl3GQ2yqUVae8bY3KkrbwyDwzEJ8p2vM+tfGh
wT1CasT3qQqZU9WkR+N8L2tqGkSYLz3Mo/vb15ukf8rYm4iZRBwLPtQXohnbWKcxIk73ylvzX+75
6z9Ub4KNG1WcvHmy7IsPPJswFS72PiOeqbxO9OW+PaYSMlTjsX+WB/BNZwHh/HyCrUJazcWr+65E
clef8pWIl4iPNQm3RRJUr1s4Ptw5Puy+oC0MVkYkYI1S+HbvQAEYBcc7FQHHV6pne8CujZVZtc1g
/NUMurmslf0dWNbemQs6YVWLt5QUVeDeEXdY9sDX4sIkOqJiRhW23aMkLGdl35vQ4vYa9Ns6pqzi
lppfuU+5X/ovamALbhHRzonPihrn5lcZjlm9ygSPmem1lGnbGqGYpziBAdd/YnNpbH3kaHw5BOhG
0z/xxRBjRPzBgxvSxC/whzKbbJhYJDkNX3RdMRj6mpjn9zl8+RQhz19meOQxvp2U2U427tE7cF9I
cpFQeVlfsiXmfHls2sos8eNGL3tHKXYB2cNRolZrdSJsloXaLbgLSSj3WRqj93piA8v6r2Jeur1F
R3s3Z8fSVKLSijiB4L3CE2ebvHnGHJIACBmox7Ow9KYxWR261VZU7n/FByWdEw199zx1tG/YiNTB
ovNorlGoW3SHbXwd4QCpQH5jlWv7rkM04u76PHa1Rook+RbOexVeszOkiSg/zwkepcm/MEtUlEC1
lLNnb3sBvqmxKSyiHAQX93Ii7I09poPLKwEr22zyRsxMFLVw2lVO0WXo2Cu+S3pQWabyGKgMjJZK
o1G3uDXvWtfoNRLBreoAku3oXQT1ECGpzGEYwbMSD2KoXJz9zi4maUOnXRYNpSzboSdIIhqfyzqq
qv4GSJ5DioCuQ1g6h4st5UxVNEJAnRNoJgwuSZurYW55sHRhweva2FkhgBJ3ZQkiCV/TIuNrNeI2
s/wbn8LWbHEYYfbfd/p9JCDEwMgTBvJ7LIUS4EguVzY509BB2cEhMb/DINyNYWezXY4+ClKwiKu/
Im2Q07VZG2nLavOfhYyQtbpT0WRE9BSA4vLeQGSR1b2ACewV9/6uSwCKIqbSRV20mF+sH3LiOXYa
CXf9ae7TXzmz/j9BJHAp9hwZ9mRSR01xF7kLUf8cH0cQpU7fUkQbOg1JsAoP5V9qUkMJulWQKclV
OIi8AGPeiaUhLHPDV2c490uiOOFHpYSDjS+T2xfGGzlKiSXIooFQGhdi090XAzGBSZyLGB+cYcTg
/5dns3julO1f2V8kj7w5eulkdzt2G8FEBpOSppm9mtZv1u4Z045q4s+MW/XCvBdMYhsdxClDnkww
1of/yTlTI0mrK6LXRfWdcKHz5d4icEsMgn8/474zluUm4DtlDrx37huYkQD8sXJM4D6ZvntZuPmb
LOg0lLDH7Scrc4+61EWhTMNpn/ZJI8HSTvsiT+VUzy9upJQ27J6A25T9Y41GXY17JWmcAB1r7nO7
QG2Bi3ksEPoroXNetmuOw2Kun1g1q4eZ6XlGEpzOibPSww5tbR2fWaTREjMaLRs+S2rPiW8Ra28e
4w00qLnkd46lCSbefDu6aQqkVIQxW/+6eU0uM5RcnyKCGIblo+r1g+gp67hGZbDtIC5a2ZCmgFR/
9+2sH5jYKI8n9hIZ+iQzIiqff7ddSLxzJykEJJtz6ddEBnDprsBUG7CdKZOEQAXRFDDClmeq/YzA
6bYlQxAMSW6uoCWPEKacJQYDAWhQKTnkO1N3sHw5R2O4MOfQ08z2GQf0AOUgugUiyUcbaeQNqGJ1
CvNzJIXla0Je2qm6me74VVj7EJ0Z6AimB7wX+dj3NMugk4jU1uAcG8gmCsB2EfkecN8UQDNcPOMO
OqaCQKKYPJ1DcjTxbsZzrWKVJdp+pksLw16Yf4n7ObkyYqF8pLjWoryb5PLpYYaWOi7ies3BJUDD
ML6Dg6qvHbARgyq7+wFXSAi0ApOFHScmYgQb2kbceOYGAm6RFkZzOntm/5VVryCQkKL2CM7exfKM
u2d2Dq5F6Vmco4ghbdvu0gu/t2PCIoW9HZ4yHknQZMigtlUBk5SkeOypf1v45g7ka3S0XVyqaYy+
NTDKVkkdk5mRcFnI7k+I+J/FFB7EW0CBv+D36StSV8Aa5+4l6NRsMKxMYf3oBCNssWCwntzSqxZ6
RPk4+sJ2FXLmoxaLR63P9OuvKwSakXJQTKl0jm0T2T8vslHVNHzVtQEUWRSADBEV6IEWGqp3Hzy9
XFF17sMV9uoyW8QDJVj8h+kalWh68Me26fOUkXCa99DIm0Igp1X4gqWfXSR23kSC265faHtHVHBm
xnbk1IxMdxZcI9yb9En2S31YZ4T81DU4dAzbUCOIqH0ucw/3zG0JvumX67IDaXl1osRyAk922phZ
k1PE0tq46DPCQxHMPlGAX5DkYM+u0RqbOzUF4b4lO/6HnIN7koqPkfntO1gv+yHlpg+nyxSLcdde
q3tZZgdwne0TafOBP0Z4noVFuoCOt1q0wKO1/qhleayxE1CXMt1t4Nh5pmc1w8jPZg/Bs5qHG7v2
BeyCtgUsYjZUqU6zfSC7UisdkviRZn11la23Rg4UqyuHUjukQO9QAy91qxsI83+LvA8LP9v0tCPJ
VxoTrNEHq8uq0fUP2LW8P9cmp+ufrF7+CPXs4ynuAmh5PRjZOhqxeW6/3o/dnt4WgvkhRyvHP4WV
yLxFDsKlKdbW/gvpKKMWzvkGbrnlY7rdeclHAa/XX191JKEDHYnegaQ/rtJLbaiosULCU+BlX4wf
9xz4IdSE19ANpQQ0NXPFCgsR6ZsBzlnC88DJ3pcgY86c5ruzaZU1QiVbWGpxdLG9H1e5MLVdYPDQ
COlWtOucg4mQoakDJvR/976KI/kK9sRjKWX2bm6EgmYBba4tIrGEU5dmnVpvPHNjO9NYmKKwjBH2
PU0NvWedeCK/XsAwyM10/ZhVL7Sw63w9S/maO9tTbyjxNRILsAxgPrCnY7bpFsSppDaoSpehyyCh
/dZ1ZPdhCj0UWMDidxt/AG1tSS3g9t1l8zv8pl8xwKeCV/0G2pMwLH07kwPZKt1b6DhUqx8ytgb6
2z7EjPRSsCHecT0jA16UUAtyzQR4G2GU5b/NsJh2GhUmMXMot/J+S3ohfEO3aqAyYbDiVCZ0JRj5
BQhTChaUjZwT5ma6ODLiMpYfOJuhbJiDD8WOO9Y7P4BEXO5KxcxQNbJrk1dK5x/yOWeepEg3bAUW
2yYl4Ekem1uyxTN0crVtnp4OAsM5QTZeOUEmrtbj9Y2RAFWkBmhtX12qHPDOBz7BZP02nD9tItkU
Yg5GEDWZoVPKBPPkw317ln/cpIaA1IUu1q68kZU7Jr0AF71IcOYGbC9sueGtqf/nr2Q/9ZK1WRZA
I+CL9gRki0TcGAzKOzvKn4WBBfBcllFt6XAqAaba2JpNTXCAysy3qMKXiu9ZW/mG6HFlVfBJgHYj
gyUU4mEx5wrLrtrEu7zd06MgOBIL4rHDp/8OEyn944Rpc7pAXKfdGyVpao63BNOTfUM9yMi1dPL4
Y+zXJHsNx3ocqyLNzsFFqPqE1Sy5+h+3haFPgbtLr09sjj+RhRIj00AO6/tLzfR9SiN2GMmbNL8U
IOf/OTyC8prqx5F5urUhdfOnArL7ImSL6u5kI9l/jiuqHyhPVRCXsVoW9Csjth1h9NQRR0QvlKQG
TLQy+HANrZPUwjxu8ek6keTcPexvGl5L4uaRwdSRemwrtpmMsWt8xMqOaidrzQwHfMWFpuCp16bC
V7OdiBBws/8gBytbeEdi2R6E8BCfTTNEeOWcG4EtMO5Q16KGOVQKXaQCSJEeb8IbOCHwrbP356Gw
Bh3ZJam37h5pE8TR7AaibHlAGB2NxVAKIfqY8k6kVgxMB/WjdgHAtFkxisn6WWnhfkHMFbQ8qoBA
JxHR45A6Ri7KN57qUf36+Kp6dKJk/BWkJsAfQeNR/PGexhb4JJtAyYjuZv+aQ+SrMl+1ofhFMsXG
QAw6Qa5NXelWQkvEXGm/S8YRKPNvD33XLSgPD7f1OXNlvLpSsn57RDJNzL9hqvGJa2fCE9/8ECoK
oHJ1O+rYJm0dWjtjgEyO3Zfj2626ZtU+4nC7eCtSG0tTTjD23A0zgsk0XANnTlmA/BVMzrVw7Un6
vjfOT25d2C9M/VEgsTe47ckB3kJWdjs+QkhmGJGgUCwAQHppPqUFxMvmJBh8+ETTR6RopXtKWJ4N
7DMR7yjxtCJR7nwXApulcjWJi8KNyPc2lxp2JhQ27ATZu7ADxIXaT6Og0EStqtVbX8AjIXXA6yOi
jaC4q5sysxHqZzUCJ9uwVXR2XPJFWMBp4T9ezNXeyfE65JtsTg/rhScaBCoEda1N90yreoPiVZXx
nuIgpeMp6+7BPzk28CqyqShanQ64BJN4KXUGzgIXJ5Ya8NOv9dsmHmvPxmz+cwQr06efaGQZ9Pyf
6/fk4suz59s0sCG2M8I++oTcEGTLUffknUrMrmobfzyGbW9pIAILrD8YsBSd50lvsBylswbU7w11
L9/FK0ClWZ9yadDk9KXNsDAmW2cFJcblz2sPsgETT8TZ60KptGhUJqo/xumaOoKSIf+i2FTOSB6w
QJy/mXwt6wppSh63VlAYNYduBou3hWz4z0qjHPpYkHw+WxofL40fg2+nfgrW+sSMnnmxeiRiYDNt
/dS6EUHPnJxhuZfrQjOB8c3Y8lQVaoLN7zl0ROu0pWbJC8v0RpjtsbiDDifHHEVlkJSDy8ocwpC0
1qbA6+724i9Q15fHX6OfSCdQoGYyyuILVWZXa0KL+nGKKhteHnnFTrQRdf4QakQ8l3/hhlaor4Kb
fnjatc5k/67w44kKlzM/IQt2sL7mAcYyXC0PTby+0X+OI8JgsvxOs2f9EQ9ADRlwYclzRKaBJl0m
EbgP5xgs7jq+NYk1/wGy1XdeY2FaqJ6dQtNcUqgREOpfQLwm9bB8FrU0eWSy0PNQXbF2JnsSlCuu
a0Nj+DvKxNZ9ttRRV5trtMilemtYOtB8YIkBq4G30W85PWppsJb0RkEzCqj0m2D9aiHYFtzTWIQx
L30r24kn/16iBndL69M+/rIfh50kq1PVU1X4ms8Dnj2HCG436BH7q6N0ON2VjQD++96UBDEKwDie
YHB3YJUTNisj/CJAivQ7Wx8cHfXtQNwcW0sgsQHcn59YAxqwLtR3bXGZ//J6u/URkf3sB+UCttWI
kLzwkLwq4jZrxJlpUtOrCkArH835n2x6kpcUt8Zn1lVraUmRn8w7xjKx3CHEH7BT++7n5S3cydXF
VvvwasAWXcTyUFIpFVKft4NpllXa9bWbDcd+o4sciglYsj2xzL5Mwcn+bFBayG/AtJWx5YcVelHK
lcdI/LhNclQjS0EmiQYcOwJqzZdNfAeEWtBQOzid3vExXWN9GC09J0nhIh1vTekuOkioLChONJo+
T5ZHYbFYe6jfUyCRkr0m8Z4subZdCf3gByWUuzGF5KVqSWXSAzUUNUScwWvB9vju/Z2lX/o84Tr+
gRm+laCeoJnni8IKiY8Y5Lq6VcDdDhBTQ2rQfEygByCyIo86Qm+x31oZ6+MzFK2kK0/xfWSMF7j7
2EbhKXmArvQHk+OsZblOx0wSwD2dxZsg2OqZPPNKtqrdXQGCuJsm76eW+rDiU9zwXsKEqUkdqS+j
PLmCnzkRQaj48IILA+YaxrR5sTTU23Xrc/ouf7dwzAd+9YLWdwRV5uMZNtASLLMjv5lxWmoUtv+2
aZ5sGW5t0UJaMec99kETDwEh4+unF8YOeAFx/Fjrx080HpQbEd9YchK5EnbI2/cdrTT5AhfdfNnG
BKe/+tIiqYVBj7lSOWfOLpJGnIHJ1yzxHs4YxUG1ov9hEwn8A3vXI7Kfjy5A5+ajN5R7MavpIvRO
Z6UWVxouIgx2kDSj7NBMm8lKai8Nd+2gIMDLV7fZZSKTTzyGiq1OwbVVnpW2MELjKigMwDhXISeO
HUEHojVY/zoQ4pl3At9CnzQk9jagtkAqt3I63X1wEcYb094nl1/n0c6MVma8GpSqtITcAKNvuAgy
cFMDJuaLTyFzp0LoQtw130J3W8zUH7O3twpcGY+dZGoYf3BFzluRgzK9LM3Xeq3dPQkezmAKyBzg
2d80VO+aQOKva4gusw0t0WJ93DSZRK/yHcxE8NkvBZYMd8StRdJLT+V9BfLNPF8O9T/2jk571yxb
eyW6DL9J0/fq2XCLM3CG+eOt9lMcf8Q9Twcv2qqxA229RdRvj6wwxKWR2YJeo813IJHwYI/QUe2O
PHwxpqqB3JQz80s3Ex3Z9cyz7hfVKrR8dSOmZyGCV91oydHb65RnfEL5rR9VjstEZglJP3yMgYLQ
Lp1Ezj7JANXg/6LS+6WxaD3i3vfa/4LnvDxTAw3W1HmBUho/P+Rq+3y0LiVXZt0dcK42OuiRfCCX
lQi8nAWOH2AUHsVrPrNv/CeAHIRFnWmJyJHu2mM1Otegw2U1tajolpYvT5Mqf38Y2J13PqO7Ctpp
8R3gfA/WlO2cybI08HJLcz5joyX9C+p8oPC4NtBTbt0BXTeUCqAYyMAwTDDcFPAxicJ5bX+1PDnq
PRNiw7s3Hs5T6vuZ3C5joFlcFgUguuXH/2jevLud5uMGxEtKJ2/sA8/BahqsGVA0TCoNt2vyJ/LA
QnPxAaLwZcRFKZMgdtt4scI6ukHpJ51dk819HoK1REy6tbFnEZ+aPckOPPBNr6RsXhi8XqJu3/Sx
86aLZJYY5aI95qKuTgyQlnDvqwCrIiPWYF8M3JyjZ5TJfSFOFvjjr+Qthr5a7zQqdTrGHOmlRNxq
z9Z8qKxRD+2Xl+Xd68d+wPK8IKZktPumnecLt8EEyGbtH9XJ2u/HQIQ6iwOSVmyQtSaOlI5s0Vvl
DoxijTbLw7xGxR5cZSuYabuHBd1InRks0y3Q+FE5nnfDRPQtW5v2xmwPtB3ArD/Rbx7brj44Ia9/
XFC32r0MYhm49nscggzfDg2LDO+q/mx5897ms77F77czAJ6MXe7i+jemmJ2a599fa1P+xLwMJm4z
CmE5ued5xinSXwyp/0n84A/+3u5rjE+fuRgvdCbKyvCQNMeyoqlUczSdLdC/VZdlVHd4UPqr5zGK
uAB9C3/8zeMNszVDdBi/3zZXGySRAMmxdF38FODZGDpeazEzpW1wtCh0l+kalaINEt5mWiyJQz/Y
GbCoiM0rRpGJEsf60/YRJiM9Y2wv2fQ1lweHJJzeVkl7hIBkkyZbrp37wXEgEwjiMWnyDqrJDVOB
qq1rQaoiQq5J1+e/maEYC9p2JHMSR7gPmYDtHg9tJqOQr0Rn6TDXTwBKYLhd2mW/ACo70/Ul5Q3H
upN+6GfeOvNqvvrnzh3KD+8LWIiRVaS/Y0HF8uYEpuh0cxvS8Ddq/4KPjJyoW1GBVyKfe8Z3v58G
9c9WNDciG7Yo0kQc0CO/XB0IOa6OCGhPuqgJaj3zdM3Fo2KduEziUrdVhIUg9woCf88Q67AI+qR2
L0ddoA4aIlj8MlTwELx9k3+QeBy4HR8Ozn85/QZ4ctdhqPTLDHYUhXru7FHOM6Vc+/2GUOn59ZFy
tBZjn4E71YyzQSlBp4njtNntuBcqYzjuUm3cXbIsDYXkebhDKra01nfY3cji4qOfeEXodojrtA0J
cCv66OLNkd2QMq5+pQFhSIqVIbakVrmz0jOA+EyRibPTya3l4uSCXSh51DkrOD42md5ApTHgSxT5
igsuuTa0Hx0MAyNx1gg1JTzrKBLPZsSZ+uWSOT+Ury7EYbspt5hCd5MIOEki58qorPwU+KkWNexo
n9+zkxF0Vhn78xqyQVqQddKLmDgnwvm3zjmWRtaO9C0oPksyNTOIco+YWbluif9Ads7t2AJX+85L
60Gc4rsTL36hhwqBWBJsx2jteY1C701UnGOm8V2SZJfZJ+glZb0K/un+acX4/FpMpdeDdYxON6cf
k/4biZFFlhmgTuBi24fDuuPN8tD6tYKJp4JuFWqpSUN4/8fX9MIh2/6/YNZwzWBZUa85Ucq0mXcg
KvDR05pqTczV+/2T/UT4sibJm4gNi8i3B7tcYXD9oi7ZN7k26pBmhzOC03Bx6iul4S6KroPiScdf
hELpyKHOkMTKzyYfJkm8TLZvjaZatm7GoPKbWn6WxAY1dk4mMifabuNC1qyIYf5vTqww/0OZDxDa
vOlnF4x/jXJa/2pKL6xljJPMYX0xw81WPbxHBYY7uA1m523ZXcHoyUyYJvO0PGeC2VjHtLj76VVw
tvvBMfhax3YmOR7Tx9IVH76F97pmCSErfrBI+hyAmEj4vF0Stjtji6ASH4VHIFsTlf4Vru8BH3Bo
xFTEIkFWuDv62BASliGl7iaq7ZvA9WCyu7ax4sh+JXxZ2EnAncIOtOAE59pL/YbBbOHD8iVyIYyj
ZJZdqEGx6Fz9wxIwOCln6+aKjTanmVN4Uq5Q39l8GF5+WNO2wS2jeW2uir9gHsq361iyQa3NV9In
LErOChtb0qTV16SziRtxNanNwA1MU5L0F/RUaBlNEB67GTUcNIq5zUC/a1M8gN1RAy6oyJxDbZ2l
5xd15dliYNsJ/qopYxeU/9jwCiE9ZMTeV1zVCnbwEqf8LgVhx+ormPQlASakW0KNGSxwEgEi9cRV
Sw8gmxdR8yOvN/xBi+95kJBMwNIFSmvsIntjfg1ymC+s9NCjQpDFVxl9as9b3+hJJUKCh+bitFYV
mjnnh77INAx/T6NKScvDt8ycrIq3l92cWTfVO11e3/x2vE89F4++8mLThydslsydRqRjGrWcqYDR
WZ6mzLM3BivRzmxH5JH4SDRlYEO/ggUnJU8C171D6NACLpGss8gsVFqcmoit3w+5T33TY6qtxpdG
AvIKcN1e1CQ8qOooGdxDGiJgpey4K8duW3VWULPzD6bQQtS8O6zTnmIkbKda6GG1xkck1jnZHEbi
HMhGFZApChgm1Ukws3iwHP0mo5m9vXQtH1DAwVr8Ow6gPl/cdd65e8+vgP3strmY8arRjG5TZX4k
0MveKD8EwimZJp3ZKXcwP5Xr6U44842ME0GwQ5k2WajoPtnfzGqcPjn+bgSW6Ca8ABNt5X0nFwWX
MyDPFOVVqA3vhr8L4jtznyflgRC/36ABpHERU97sRvmxHwgFfCscSwWI651VwHbTJWtNjDlNgySJ
k2dWZU1zNkkOAFCNpjRN34nWc3wLkCmhsaPQLtf9ZCBejn/BDSh3XGNrCZEY6VrTJ7UDMr+jv+TU
zflS7U+Yb5uIdqRfs3y3Oj9SGc0OJxBcyrII1qmCBjtSUPRGnVJEcYN6uyUwMfloBRoQK44vlPE2
lVr4Z41PHDUFWAwWJd/9qMNSxcKvmLemXZjhD8HHX4N7KfasVrZIzILYBxm6d783Ji+5qm8lGV4l
31hx84KmPbhfwsm7+sSqKBdB2aUDoL96zzDljiYXwembOfq6b9UCB3AoinJSO0O6hwKnyYP1ODdg
TetGcQB8+ZJ2uUfeuBySUnTeNGzsjU7ln2gvuC06DAzif65CnkUSp8VDEpXdIQWT6VwSXcatQbk2
CJKMUtRDFQh0FavUCkyfpPf6Ry8KIV/btc+sPXqzEKsYbFPMzcF0yKXVGr+hcpon5hanJoOvmOXH
91m5ZJlFvjajAgryo2/FmsP50dnGshY41ABBayzbiIMpfme1tVNm72YDEykBD9mfcPtCWKI/cTGW
qvndLX1VsjLlx5ZZzpw9xb5BctaRCH6elOvEbEWAf67K6pZqESjb79A1a9O/whtZEuzgik0NIcVx
GtJ1bnmVhKpjRaVUkmAgcmZQ0G4pFT9ARZ29a2+iOmtu6Y3UPvRehiHlviHwdCcE2pSiki3uj7O3
21wKZZ6+zwYCSkrCrFDCjhxfU1xYbZhaWlfVL8NiBDFJAuw6PVDv/PgUVhCq2Z7iPBPboUglpYnl
KznpBcc/1nIWDlT2Lf0FQMfrRXsFRqV05VzumCLciVNglsw4N2TGhGvCK51luEY2D9nAtvnbg+d1
PTa2bclF14P39NZD0aINzQ8jde9HZFDmZuUHMAYs8qQEl+Y7v0IAQIU8fQwsephVF/4/BG2Hq5tO
WX75c09CKEsYRtgas8VWNqenl60aNh5BUXfHI9XXVswdsu85t+2rlKuU6+Z32lMe5X974psqUcLT
EKGWNnHSF/DbfuGH8rRdieDKsBTucafkF8mcpXBpIjMnfMp6iCMIHt2iJCGIckIlqQqDQqe6auRD
Ze6wEMHy2uM2YYcSZ4DglcPeHAHItLiV+4jonAYzEmIJ4k+cCh/uXVVvvIs7DbZQkwtGHVv+Hss3
/is0oxr+ZhmtfQ82Xb3TdRMnlH3D9OL0B0lkahFKTZC74oMmtIrJTzE89vloJiv44i7u26oqQ9d7
XB1QJPAQDdmKZWs3mCRDOP9Qgy1DanQzCql+AK9zrScaGEMLKI7nXlTJzu8gCZNRiJLOZGlpDvY7
rFfHvSeYR/Fq6UiI+ImMJSsnxcFNsVkPQQ7ISCwyHoTg1Lp7Je8ypEnCMJVqWMsjpem/4SwrjUHY
0LU7YQxJnZgJhTqTuVza6qCj7w0Nxa/CiSNeiBu2luypJWAGn0s5EOi47fHjI/rQV09n3EQowGPu
14ji1N6LJg2L+vVNCYb1H3pvWe2SfmzqmNrOmv+3Rr78oKksxm0GEynt3uBdP9KTysNDmMgbIw6y
E9UMO1YXjO+dWmohCR/L3ntSw9S4HbbRhrTQXTA0UEhXrqYymIyQAfZI7DvAn+DooqNNOFfcgZi/
Ds4Lv+OD6XUUspHNNav6g+DPbzI9uUVEtqeFRHnpCDHr+2nbifEzpEh1vYHAc9sKs5YdCrTKjpXH
XRdj8CLFyJLtsgJS8h0kl69fNDxKCEWuSkHxiN88Y2ux7spIY9HWeRND10hTEG7IAk6vR8m5MdFS
FrPxUzw/3tlTNCOHDFAC1x9w6Z5V/QfV0TQVVZFG9RlCLUaJ1rnpnwBdIlyE44flS0VN8CNQ/eoQ
WcTWNsn0k4+VrqDeL1kRbi7d9jeSwN5lxWe+VFW8+aUL4sQxlWxWYGI43h44i4ITSIGL1gfukJq/
FgR5+Kpar8xzh2G7B6/ndn9wPPuWbP319CLv34QSHDKw6kPDQXcUg2XNqtgl/qn72fBhrshe+saT
tUZNLoPv4ftHlvuaHAsEW5MY1bROKpFd30Ft55NhmU+k1AJPCq8GMFsBbIJFW95yfqCiWT8s/sUO
7R2wDNFkFpO3UyzyAHV1/Dfdngwj1FzXx9RFcrBTW4yhWPxirPZJrMNQ+eZKmrpo9y0yj0P8kDtv
XsT0HVx2oH33mUVaUtdzQN4ul7fHQIPW6yF/rQKbtDF2j72iWerO0cTNZGIeON+QhA1nia5iDekR
Bh0oQvMpOpzeY0I/+A18SuTF6vD+Ctmd+j+djTj1IxCakuivIsxChl5uLZX6AyBpc0mZUnNdcYKK
t9DLyIxJYvU/gYS0MGGrimkDWprschchDBzlluxaPwrxgRDyPJBXkkotpkHBcxz7x3x7oia0x3CG
jQUZ3ciMxXULE78xO0HJF33zfF8dj2pfwGo8w1hoWL0//AW5AT9BkrRURzY0kv3b6VP+CEJFS1fM
EWWnVQTi+HSJnW1Lhj44/NHMUpE7Jr3wIRFT91N5u/VBIG6YcFoPSd26KtnVhghNXnc/BeVrhy2o
fAhheFgVdHO+b4WQ4J0zoHGb0Xxa7pTUBWbmOSUOD3tWE1ypG4hOnUZn0Hmdx8jHAtIzNycxEgmT
lMNy2qPHniNpnjfu9VL68m/OFm7htRTgbFSAxYaXX4xG6K8LtT9e2lfPOyfQAid8MNmN+88TGTcW
NlBNEricdrphl/bkrp1HEqzZqvMG8JNzvRkbzgiAPr5OMuTNKq8V8hLSS79PCiiRhFSmi+EpMcxT
GD3SOGxjFYZf8mlQEvfojmwSiL3BWzk6CZYPe/J5R6SHDr/Fs+tqJjFrVi6TmeTXw8kenX7zf8Me
5FwU8gRMDM0857cPgOe3erecFNst1EGV5Ba25IbeXCNNgoyA/00FYeLLBskF/MD9qc2e+oM1s6Eh
jrl7y9BF7ymz1P/Y0Hq7bS9JWrdviGDGrgy4YpWCHmPfsuU7i/FKSvgHiL5oeonxj4u1bkGbpLvE
PxzpF1vh6cewRUkvBxU5SiUIn/qxscMgCHuPMqnhwYjNtX6Cgot+btH3fv1Guw+5iCLL12ikd5l+
2A+eYvipPAf+fCdK9PJrOkMFx2f1iafXnaqE8y+tT6WsZkZN1l1BXRX379Rl0NamYPe0kAoGSnih
Z/v7Rovjmou72qCMchZw0cWH5TqPrGiyt3hWC8FzS4Jp+vJfjQNyRq+jbRNtAMZ98PgoJ1LKSL2I
9lhOTahPcvUCdTjTKYE6InPUn/JS4xZddSFN57T7wryuWWQ8/HTfipGUzrKEYJ/IPSvdqkhKEtfZ
/WVxnwbBDmH8Q90UQ1PWzupLI5rRaY/FUGuDF3GDR3hGozUapXiJU2fEAcm2SA5ZWSf5/+AvoOi2
fvrxXSNsL/yVmC4sJGgxEzXfKJBnk9blwBC/unTm7yBQ3yYgUxZBvEdAD5i3L//aoNfqxbSY0RSc
lw7YhbBsudwgy0LNFLghl7nMtSJ98pY8anGBW1NruLWfXvI10QfKQSlyo9LW3xxHK731hhsrdc0H
NmlaiggQxkMipqRoM5CMgRKuIuQwx3/U9Gakrl4S/66QaPPyotOM3oFveF6QhB7U6ZuZA1BY81to
37Uhk9mQkIzCTb7oFKYJddHz0imEpB6oeojNjtpKwJWoErhbVX23bu2FN2s4WMOGhJ686gwg4b9S
WLIMKd3MIk77dR5pSk1zVJwpupPr+azY5M4m+19Q5J+4UNeAmMOcDqY7u0sFWhZRSSAkEbNkswsj
NwOZwRfegaOcgbl+xKzxc+q/aVTDbz0s5pV2NL3j+XBsJ5THQBeRTXBZE/B/V1E8znh0K8DT0HBB
LIvumZLQCkl9BNHcGxAk+Dp75f3Lnd4ABDWQpT80f4UtHYO+cjWa095PkQiQeG83fcwbFZNkbmbz
gYw3yQldOSKHFZJtph7icMJNP+pNDdZID7OLvt4BGGU8gmMQ39eYrWFwbufKTFeLO5gV9LQncA8e
A/NlGgTcBWfFFJcuwzj8iLHftOWPpneS0fmGxh0qMM2QgtExUQjVtzuwUKP3F5ziy94t8Qn+J/LD
5wPvNaJ2wM1ax72uk4RUfBz1xdbjqYlciNfX4OkMS9+j5cjwTcHJJtNdIa1Krh5ef2yOdDBMkUzQ
ye2zUzAUuEwtqnx3N4LN5BdUFH9obLRj7E7nCCnnBf/d2s+51TKSz1VLboE+q+dMA/J59AKxz/mw
0CsUmDtgVFbmojefpZi7oj8RNFE8I8a8xjg8hBQtXPip45znt/6pwXPgWIWZeQMiMB63XoUJxf2H
X0tTo+bkphQIpQbyBn0FNlnX+Xs5MFH4v2YwdqENAoqlcxjD0yUTl8GVsqSp7deVWBNyKqc+lNu5
YSsdx1WK525Z/TuD1J43luITMUaTzc9bU/iIjHo7QGPXirRmwbAweHC4zc0bB4hnznwnnXq4lCNC
AnFd0mW2CA+oK4WY66EgL1nWNAqAVlXwyr9oU3ysZDc/On5S7G0oK97bUQKCcCeWjwj5G/pLF0dg
EKs38azTfJRLxRkrsohKVaZibwAgGyXByjJQ2KlWdB1wivkxbDP2IVnVSoxa7h9gvMeR+OGEUKlc
VTsr4hk1aVIj8Prlvqs5ePkYHES1fVqRaA4pk/m14i90y9sZNS6KHYlqOjHQCrQPSraLpBlyfpHI
fVukplW5o8cjSYKlgSnn58sXqgIkbwFG7/QVb1l5oH3U1DLkSGyfEZzev2qkURhGj7D6JEFoM63O
NLQQHSVrF4CPi68resanXWW22OqigjgBiAh0wcR9XaK4TyjE800Sk/UX55iVe8RyeQCLTrzIsejQ
NowdHMep4bc/zMeWmSib7VkqIq6/oSQpWPfwCs73KJOgvo6BXThMlTOJ9RwBgA6jJKiaNnxHPWUV
qDX9oSohAMOUhGNmuPRPN1xsn/2bTwIxXnmkmWyGBSwvpWF/0I+M3ffjJQ3EVTSINFOsXLhDFw7x
Hf/V2JbqjTVrQf3klWu8WPUoz+JU3f6y0exMEcA5aKWPIi//dJTPhvV3JAYfl1LPSGN3V5W5v9M8
Ne7mLGCOo42aZyAQHOcUgfYXGeFqDGob2EzMSBww5fC9M26xpe/8JPFZvDfclGadrPVYKdK04T2n
L3F5eycmcXpI27+MHaqO4a9SMZ/gc9ExAn9NT8HjOb55kVxLbJ/rwkfCdm9SXdaDIZfr3XEq19n+
1Mz+fFPLnFOELDBjm74ATH8HtD9VCQFZ1qtVAoY07QlwLkw6PsTgDMQiZlZMEscengAsUp1EXaDl
TXBwlg+Uy3s2l1Lv2WQaqFzF+uZop74urUKApcKRsE3c02ToTnBax5zVQrvvI/VPVbUt8rVQAxqI
r9CjMRx47vMeKvG4sBaN+WJwQUatibMx20Kr8S+ElUL/f4knOBJ5oaXkv/JACmCnutYCfsA+Wzqa
BubPe8CHQhbNym9g7BlGyH6Q34Xl20J8pO0hw8r+bc87PDXavF4yMN0FY3I6c8qFCiOSCJH4U02L
f/yi9yRAla1QUD86wUgZi5UX4VEUzPivpe7GwjSm7tMADw9KBerpXU+bhH0vFH+0vnbt+5Eqruu5
tUxKLIPgQLhT/GIdWfhNTx/PcoFKK40xbbhZOos3kG7j0R7k0lyb6t42nUd8YzqACdt84IlX76ih
XLciP5K6BgOlrjNer1h1FI1D3PLsz0vH34INY3iVEFroB0tf8UMmwp77eBTOqulPIllJJmlmI+aV
HvbUPgRhUgY4kgeFMVoBayJl2VtZX3TGApmznVo4/eU42PRnW+rMg2XRXAgP4bRB2Dm+LlkhU25q
NWQH3gSuPgSi07rJMOs75ILLJgaNYpgeUQTop5yo6QotdHK/MTTWyyM5xR6ZdtRP4Se9Q/waENXw
K4gctNia1FI0y5vuI85tm5f8eMOrA5dfmdbnk6pxpgDc72h26yMkglFYRH2MYUPyT67R4C8Sq+Ai
8H6ydN8pconoauwaCW06U+RCZ7dYTvmSs+VnMuIGHbic9yBHFcA9yQmmd5PLRKwS2OG+YadojXws
i48G5gQAm2RvgM1x2k0cUzobL33NU6FYP6tLfnR2binoyEuQkgxwxd/55lEh7BsfWl9XCSROxi3+
yJzTWQGlmDmf3MVYLuK0iiKGB8ALfE/haE7N49oMJnwRUK/yk6pxUq2pySMakOzkZZzZBa24qy9K
37gmT+WJSyaNAew7ZwrtDjNn/w7B/rOGHe3RtCBAYG0KDZSZjgNdd7z7VbFg/re7RIDwB3Xnnh9S
X4g9VIzfIWL9R+GJ3ZwUDqNj989sMNhp0/hLC965iKITI7Qli1XmeFQ6VAZevnHnFaei5uwmwj/1
sUqE0abPb+22ygNuUneL7dmhFSpp89VgcPJ+m95iD+nhKncLhjxq3wnxmQ6mFOQTAbLoY+2nDq4/
K1iyN9xJkWteyZGZerpKK58dru97WfqwnMpiG41tyBqjprWM1K6cx1yL4pOktXJLcOx8b2qZPiFl
W8/93yvbhLHbBMH1kYOdRtg+EeNc/7uQ4wKQFUjuQ8tzMLKYrbt3Po4bmZsN32RFyZKTeJbBCZV1
EzcE7ZIfsoQD0x0JdMytnqYGjYk4ZGen9b0mlBgCshJ4xzFa0LbJrQZ/aNPBUvwcFFd2g169qksK
SH6BnAYbW/rxNEIY/fAHxDMVa/8HeX723jNY57XTX1/THBlC+wx34yuzTmA1X/FdOj7tzCd+y9I+
67PkyOkoxTx/uARaG1x3cpchtYEPvPNgRlBg/MBQKWPz8jerN4bt0Uh8PTDjhHpq/wvas8Fi5FzL
ZgvOKzFKqSgHr1jvrc5lidqYtd+7vSww/nVkHZm4wvSFI69vLLdscZidWVopCkw9hosk+PKkEu7B
YuUB+yifLaqTZQxCXSDlz3kVqH4+LCQzaHn+kF71YKh7tpPhqgQlyBIwDFNWCMrVOZjVv+eM2Nvz
4sPrAXfPiOMI0dlXL8ZyBOBElEpfKgh0O9g0fWj5WkX1Kfqj6i+sZmWaD4BVXBk2sZKnb7edWe2g
ehShD049MZazYQj0wvfic7loSuAAtMI2KbCWgHKdgOkOVh20meghfTfF3cGsrtVJb9vgfTSP3eaT
DXDc2LPzKaGVRFSNJXJxB3EU7mCW6JzjP8HhAnEUHQ3nZqLeatp1qjis/D4tp8GeVweROf3Ft9EB
5UMXr9OkOSp+/ptNqbBX3SRCj9/6DI9uMZhHNAMAjxSp1bmMVBk8wfjISQvEaH6qioj+KA4lP3+e
Hu0xBOTQ/zY/4gvKa6MMq9lxAVyX8CM0+HHJB7d+PPkpvpK395yyJCDvlEtJ5CjEl91TcBx9N7/R
RQOnMUVwZ77KiQ2bF4ss5yZDpXIwI+ewMVIa4M6rIj1yaRSWyndxtzFH9QDN4Sigg87MF7hUGCnl
oVh7rR8Fpyt5zdobTKFDF0eTD1aAmzKm/NqMsSlZogtsWavgLi4EgLoQaC66A7PjRDLqSCtlb/CA
wA65pBijtO5OV8FArix2cBA73EyjGih4tLKhKtLhiEU6K35qEePnx4hSN/rQ8+Oa8+OYKZiwDOld
xIbGZQ2CmUd0xb5wWVJxkIB5+MTfr6LLKM+/MmkGviXUDOHpsPoU5ssvdwlMQeoFlMo831BKSZYN
pSkGvrLTN/WncnLkKKpcBzBrZfNFpKTyLyoj90i0hiUmYG7WcYHijdRQ9YXuhy38Lz+iknWZo20r
0r+0yps0RzH9o/MXoNQjepyx/PiQl5KdV0DokP1VsEc=
`pragma protect end_protected
