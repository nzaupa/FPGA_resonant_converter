��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_�����Ξ����$�n�?��3���~��2�j
��n�"�4�	f,	�p{e�C!(t^M�G&B� �h���C�{�TV4�6�!��z��?&s��(LW�t:��K+͖a���Yו���]+5O��
!�����`
�(d��-�c8u�I�jR��OCդ&��j�Sh��|��w�q����`g?������O��aom��D�I�4��O(�h�pR��B+�n���~dӷy�.tr_]���}�iy�(�� �k#�Z���Y��/�[���z�N��{&���C(��h�\���+��@ZE( �;�0A�+�L� *���X���I�1Q°�/x�
���P&yIN���U��m�2���
�=�J~������LSx H��O���ǋ��sf*���{&ItЪ�5�.[�xL�:����#YF�t��*��X7 ��W�m�MP>l5ۈD��1"�/������ks�����,���v\������ f<���LU�"����g�-���<�
����X��LG��iB]��c��hf�ղ�4�����G��-]��/w�M��J�uۖ��
:<��<Np̓�XAN��d_g0l�-Ô�m+N�^�X^?���A�hd 7�=�k6�͵YZ
��t�׸��?lYr����H	���Ѕt��44�z��U��Ma;�~�j��a���^.E���s8ЈF��_%��}�Vۨ��@�׹K�����AcǛ\>]�\?��aU�7i���~�k2zy��5!�IR5�hό󟐍��,���q!A,�=O��nI�(���󳥈
�c�f@���>���S�y�*�$�ؚ�|@V���l��L�+5�(^͘Y�pC�Mjs̭��ۺ�D%K���2�Y��`%g��8�c؜����َ�=�c�m {��cf`�{����f�Q�@�*-g��3q�'��z��!;�.���Ա�޽w�&��A��T����mV7���l�J��3�r���ͶV	p��4��=.�����w�Rx���LN��7�Q�f�8�_��#YS��u�B�������Eso��A� b|�@:p�&*�6�5-2���3�:6�����"Hi[�X�JM�	�¨��A������r �w��#ܛ}����AA�ΫQJ�?Z����`r
S��&��?������D-�Lx��vZ�'MYM2c�����s��U�*��R������vRv*²�����'�� ���S���?�N��c�Nђ"����팀�Q��������L�~(b>ʶ�ztf��C���C�Wm�|�����[����F'H�ӓ���)'/�7ڡ�ץ3J셄��.�3����;��";$�ap��3��_�l����5�zԼ2hWH�C�9�l�D����׶<$�-�PX;��:����QR%W�n�_�]�v�XŹߣ/.-)!��p�o��)3zН0'�����F�=Z_#�~�+�w�P����3��Y�t�8�×�<έiyv�B(���L�Oc�S�悡O���O�d��D�W6�?�wy�T;�oc���g �S7
��Aڐz����CcT���	:%����1���ޮ������_˶��+���G Qet�Ύ��MؤHH���K?�}�K�Î;m�_�`�`���` �kw��Y�TqQ��^��Or6��97�8^�u�_Y�nP��ôOO��1!�rj�d����I��F�V����wYM�kF���8�܂��?_
�^���=>}7uﯦ$�;��{�Ǝ�X.��!����۶	�
u��Pщ�D�\Q����mAN�`C�G=�_s��/�얯�n�usUɆ?��p1O�>H��g���`l4�j�	�A8�v�>��2�� l�ڗ�5��Dv�{��=��ujO�����oJ��`�����e�DA�bݚ��lM��MC���hާ���%?&�����z%eݧ���ZB���7�7�zk�q%��HT��?�#0�W�-���-
Ȓ�x�P\��6�����LǶ�v��6��T���@����0�л�SB�MWU��s�@!u�G���OC7`9���a��R➦�1[_Hq7�oH
:
Ԡ�zw��4u�����@g^Oݐ�k�Ʋ4}>���m�_7�7��YA�Kg���{b�ϗH�If����VQ�(p�4�Q{!I�r"�0b|2E�4R
d�!$��8����`�?fS���Ѓ�t9{p3��@-��X���I6�j_�����J���m��r,B e������PThMb��Z�2IX�D{��w���3H�����$�����G'k�jϡ{q��ç3��Va�[�0v�#�E�J䠙9�9�Nk�d�~��F�4>WbƤ��i+~az��/��0-��I(�rMb���\x�K��J��B�����.ؑ���W\�_%�*(�k`K��e��O$9QSLQS���ZgXnv\��1���Ä���~F�%������i�HCkhG����u ��d���}��΁�y�B�M�6�⭓>�O��{�$��%w�x(:;� N�q7��Xe6�B�aqC �dM��)	�(ҹ ����[��;���CGn�:_��m��(�Rjy(K��Z�urm�Ax4���X��f�Q�X��Rc@�}FU�x���T�SHL'H~]��%:��G8���nmr�[Gm7J��w�#A��*�
�x���w��5��'9��G���۟i�s�y7����V����e�t�kPG�3�	��TZ�v�>�I�bG	^�|VJ$�He�
��L	�
�ӥ�e�X��f����p.�3/I��L����L��ш 2�k7���4�g��Sɾ٭�Ր�ֿ�<�3�R���9��*h-�3���	�m4�c#����4g�fܫ�=Ԍ?{;v@��M�;�"��5�����X��b�����0
�2��N%Kj�=9��y�V�!g�P\`yEY �?�(Z1��3�Q647>3�:
�٘�ù�pлK�3'�,�X�D$��YB�HB��J[�S^��nL����=����]���d�(�/����ؠ�}�����./�"��G:r��2�y�Y�/�9��y#2Q	��J��EENNC��u�)��ɔ�7�V�F6q%���q�3�����z�Jk�R�aˏv�����ڌ��?�f��cA ?j�ƪԂK6�Z�!>w�C�	��8#�c��q|3:�G{��Ҽy�>�jI���{{��9��{*e	�֑��D�ݞVbc���>8hf�h%��$"�g�����	�CY#B�:���7dxv�p�$�����Z�����p�	����s���sÂb3V�pP���1hj�<w�{PkCl�n+�p����IR����OXM�j�۬d%��ژ���KN$�o�6�+U�c���&��0vJ6����e��!���@3	ݲl��//M���6�_Wg�ê�X�al+G��<�.�eB���O*h�[Q�#�N<���CT���Od��|����T���νa7<x'1dk	�#)?R��G�k�}�AY� ����hP^�
�n|��1.�E�J��0삤1L;�Y�fK�t�s���6gf��%��� ��)g�!����Fr�)W�	{�G��1Ԛ���V����>���КԼ}�jw�q>����)&T��	f��"���{��*B���ys?v�Y��.��UN�d�޺��?'uZ�XL���8�����	�~/�Lr�!��dޖ�$ʅ���~�^2Kg���Z���3�;a:QvG����Szp�N��=��W$�[n����d�zm��{1�}O�b�>AV�ͨ�BSn~Oglf��o	����T��操Qd-�Z/;,^����)�d��Y�䫹:�i�twY���1�/u�&�j�54���`}����ۉt"��yP#�4����n��&��!�~߄��:&&獭�0�:Tz��I�� ��� ��t0�����Y��ǫ-�N����¸s�m�����/�5���lv#P� �h���%(]s�(j\QZ�yی~e m]���)��,oG�y.L.P�ש�b�vuW6}�3 �����X<�����f����	H��V#}���ʒ�VٿK�%E�$2	h[�K��ny�Yy��6_%���#jw<Q������~�|�����0�{ +;��!��Q3�C��񨝉`����EV��E\�hxW�!&G�ez/��b�!ОB��й�c�@@�i���MCü��V0&����f�|99�<V"���m�뿙Qm�3��8�H�߷�~' o&N��\����n-h������d+�6�=a�ӌ��X�aZB'�o��L���ܥ���=u��$�>s��<.c:���]�u͆�^7ɂ�@k���9�)@�#X��4�%���j�(��i�vͣxꅄ���fO�%�Hq ��D�k���ꤼ��1s"�/�P9fw�{�n�����X�H��Q��1+#M&�#��+�f�tQ0W	��W`�]�\��\`*i�Ċq�2�H��߆;����5v]c��׎u�7���j15Ϝ��4�Ј�S4��O{~�ܺ}a��Q�3��P�?��2��в��Ģ_�OH�5K�(6)��fl�GI	����ٟ��B}�^����XssL��	�vZD�xC�A�K|��[S�b���
�]=W�%��;A�l�{�>�-��lNN��L��,��\��!��E��~V5�ex��SI��@� b��㧵����6¢[�ɠq�ė�| ��ڍP��l��ϔY)������]�j����43;�?�y9�r=[�96�'5�����&9�j�R�8
)��+.�,0R���s�	�&,��dux�	�B�%%{��*ߡ�e�q���gB% �, ΁8G���.w��n�����0|����㴮Kk���(W�j�b#J�m��~��s����/�'�/�RS8`��Ȓ 7��>d���Qc�\
��Ȃ�O5�CDJ'��x�cr�p�A�����c��c����F��;������-�8�fm���I�r�Y"v�ZP�W1�G���Nʚ_s&#!�+�X���y���_T6�+� ��ԧ�� ~�$	$PP����#Ԟ�l.�!T�.T]c����˦�8�Y���8C2(����ϑn*�&�Y��`�}��*hZ&]Ki��)t���h�0����YE�ta�je5:�#]�%j��~���l@��u�eR��&�e����kM˝䵂��l�>C��,��X��fj�T�?�Ε�M�����0d�*)��s�� i�ç���V̂CX�<�?�͕9X��:�[������5��|j{\D�\nm��D�'��]f��N�2L��^�,P��n-��en�Ȩc/�����i��A��lUX-5����V��jUpK��|�<7r6hlf�;�P*��7��Ѷ�N�}�FƱ��@�Øְ����׊B��a��\= L�V�*U���j}1������F��e٠�ڑI�MfL%k�.
��Q��|�;p�	��;k���'+�{ݝR�}�*�jl�L�g�N�/W%I�6F`_	�,��hLȈJ`��Q$�G��2��7�g����끼���f��`����(�v�Rc5���_)6S���x?�m��>|�pb���oZϊNb�'eQ���X�'Է�<�R@`��8a��]�*a�З� #�$�3����`|��.}@�f��L����Ьț�G	W�������q�����̍�-jW��bM�|��(�.A�1��ҭ���;���n�b� 6���g�J;���Kr��e��W��x���wr����q�������%���AݯJ_���D�|�Ъ��y=0���y6�Ao2�Z(�/��_�xk"l�(0	,��ВZ�y�c��Jg�_	�`ˤ>�K�]�25��Ur���9�n�G����W~�!���{v<���@<el��8wm�L�EنFk\
x� �#r�#����PhϚ#m1��ݗz��'8�#����.X�r�����.�~Llc¡:^}E��߆!�ޥQ���S>�_������%�ͬ���D�ɪ��ō�/��k��Y-1N���שC)��+Pa���e�᷹P���iPv&����!���s����ʾ����\m���[�x�Sv����r�U�x=\��|�)�|��[QcH�O���$�u*�{
���������-�߷V��k�W�{����o�������q29e�`7�	��)Lq�-��� ���(�����c�Cy�|�9F";�p�e�����}(oA���W{���~�#0�XF�3�nen{�Г*up�v�o�%������H*�c.h�H������A(s�
��_�����?1$�ضCr�@��A� hZ,Q:���]��=��"�w����As��1JdC!iK�~ѓ�~���Mvd.E�_�A�~��w�"Y����e|��x��8ͣ���'떁�3���������^�hɧ�n�,��r�����|۸��cn��T�V�ţ^����
���_y��Mk�"G�-d;�/&�:�V!cDK��m���s�1E���7G�]�c}�Ta��a��/�H������MM�G��A-�4s�V*�TDJS��|�)�\�l��q7S8�N���EFvEB�`9^D�rh<M')B�[�'�悛X��zc����,j;78hpGI����
Щ1��/�i�֜��Ƌ��.�V�zL��;D��</|�����i�������?|�'��J�m�ƔI�hl��tF�z�f$����ϒgp���%����A�NB�/2>q1R�֚����V����I�r�%��U�WRA���q��"�4\y��N�P��t�K]�M�B�;q狕?���%�)�u���!>��A���Ԇ v����,:>������ޚ��iq�kI�����}��s�72��̠�4�'�"��u&��Z"b��B����YՑZҜ�l��xWW��)°�����[�f��PQ)y�q��-b�<\Ef҅��wf��N�㙭n��Ne�J�Z��PSY�3կL�FxN�Sd���O%i�"x�3�
E_��r��A�EA�t�m:��{H��=#��Jj�M��Z�V��Z-������?|E�\��a���{�n�Nu\o�.�nw�t��&�t�
L{`SpX]��{�m�C��|�����#�<��P��f����)�Ĺ����`�VGE�J*�c��	j��c�~�����������׸�0�-�Ou�!G�yw��E��)�q�������s���"�kZeX=��QB�x�E+�,�O��N��rvH�ټ�:"P��ķ�r1��H����t/ʔ?�O�H1�O�oq�ZS�S�P)���=��i�6�rSt���'�6^���{+�`Q?r��
J�C����z=�k�,��f(Ѩ1�Wg1g�`^���m���,a�v����'eGh�m���I�����<Y��8˲l@J����V4���=�
	����g�H��"��q���������^q�U}V�1��4H67(�w�c��\	ӟ�6��Z��� �B4a����ʹ�x���sei�u_��,����KS<�)���i��9�"����!a��v��q�HAZjQ([yy��\�����̡}�`9eqn 5� 7}fXyv����S�P����襷U�l�Q\��ƃ'����[qa���0��F��Ak/�2�CP%1Gk�B���qԤ�jɘ��{~Z\��eԆ�-�b�H\�@Љ�Y�n��JY�����������s���B��9´J�_��uV��;z�ڹ��:r��x^ ^,Z%G���pf��ն��@ϋ{(���Ӌ�%��:��r����/��W�6u��9�2z|r�N�쎗����d�b|Jy��tu�N��b^�Hp��y��T��}"$�S�ĺ!gvwo�y����#�1ʺ��Rɉ��F5�Ԑ#��*�ϟ[z
n�����o�EI�����눽3���q��bG�޼�@�CƱ�]8'�P�<���v��dZ,)E�>DN�z�@*��]ʂ\���a5�Ph/�)�|�t,�^a�m5N70ogP�#(��Gg�N���3��v�Re���{!{V�[�����_��/�>�
W�����%~�}���T��3������Tf��n?�/Y�
�"׉a|�]¸Z&uO��h'����<L~2:����o`�ϵ��y:+	��=���B�����`q��Ƿg���d�9}nʻ}���4jǛ�gP�Pq+|7�녅<9<6����+����$����6�KQ
��_��E�ɥ�����8����5΂8�_{�У�
0�ꌀ-�H`�����M��l��P�Kȫ��,�����*��O�8�����9�k�c,V˹�[\F'���_�ŀ��Fk�:�T��V$��ƨt�����n�j�E�NHx?���!�K g��F�)h!�-G�uښ�f��W�Ɠ�MD�z�N5"l�}ꗼ�`2��9q�Yn^�����
�x��ِ�'���6z^q@,����yVo�É۔�r�O�_�S{s.��㳦=�d�z��K���e2����M�B�B����Uo���*��Y�����je���}�$�5�v�=�������ߞ9�WP�O=)E�V�t��C�>2�vlA��5�=xh��.�ܥ�S[C^�H�g��{������gg�s.�1M�N�ߣ��
��MW,�§BC�{u��D ���FC�-�ŗ�NZ˙-���0j��u(XqֆI�E�*��S������bJHf������0�&3{d֔����:3�����pW�IGP�����
�	+p��)쉱���~E-�� ������%�-�$Xy����6�%�j<}<XT�"(�����;l��񏃤(ӭE�Yeo�l��8��g|Y��*�;h xx<�,��
��ʑ@�Pc�m�P�H�f~�.)��W�o�h����~�F|��lq�Z�����[p��M%p���M��1=������1ъ/���@��C�*Z`��f���n>W|��99�~�h�/�9`5���m�rԁd��)�@�v�8���8�7�=o4�e�Hd�Ry]=�L\AF17��Â����u.ω�]��%H��^d{<d�����m��b�0�{ ne�(�,������[�l͡��9�Y����w�i9����x%t���.�	�u?�]����9���h�����_`%��;��G3z��H�Jɢ4����R���E��]�Lc����VG�xGOڜ�
�!�#��x6.k�%��t^��v���+�!��=���S�`���Y���ċ#��b�x(S*�~�3���B;����Z�O�E ���=c����������h���ln^q&í��3�K�����axC��{�S����b�മֱ���j���$pv�
��pf���vS�g�� �%�`MTm�X���Tn+->m��]��A5��F��;�Q�I��*ʲ�"j��e���y|�)q�QQ]V��PS	;KYbn
�fo Ԝ?Ц@Ȭv�0�̙D]y�e���Gd�
��A����d�BO~��Hy/���6Y���=F�`'jx��f6�%u��^��.�����vq��z�D����~� O�����	��0IU{�nA�����N]kk"�BE�Cnpa�ƈ✳J��@
��O/��0�<�r����7�=~mD)���'c��i��f짅mÀ]1~�V~�`�s��Rp�%
�x�Y7̾��P�z�N�%?���_5np�FwTiF6��a����VJY�⍝��-{�[v1�YO
�[�3B,��W�u�Hb~n�o�(4̡E�Q����LM9�Szu|���|t�	�˶��$b8� �������GU䮡C�g�OQk@-���$�\Q��0�����Ԉ�4��~T��J���o+�a�>C��ջE��ݻ��j�x�EkD|P&��`��bߟ��5.7�c٦'�ybe�?@��L��u�-�H�_�#�o�F������D��[6>Y\�'�M���~/�q� Y�}`���	#�q�xȘ{�mSG{ʍm�#l8{�=�]��ć���);w��h�ȡ�P� �����j�*�������-��Y��E�i�uH�#0YPĄ���*�����`�����25��{� 3M޴��d]�-?�W�H��6�(��^�DN�Y]�D~���x(#�_6�b��9��p����8�3�%%�	8:�ߣЯ�C�(n��s�)�2�1����7�i?0��>[����.F�Bk?��(�����W�0��܀�>L3C������,K�(t���� <�q�s=X�y 3��Y�>�^N�?�P�,n4H���l�a%�v�)����V����'4�`�����Y�c !p�8j����S�"��S�Y���>n�{�1�tE������S൱wQ��y3�������T/<V�N6T���|L����u�`2�p�`2gB}5���<���Rg=��U��#����g�����=���R���P��oq�VHl�,e;�'ת��J-_�nTw����`�������?�p*tw��^t���R0�0��O�@�\�X�� ��?*u��z'�.��f椟l�i� ���;�SDL�^	�Q����� ^Da���G��c��Ŀ�Y�+�UE� ��/_p��m���ֽ8e��� �!�d$_�Vb3��֨TMO�Xy:	��0�?$o%�8C6.Q��,AKH�"��|NI�Avl�Ls  +�1�!�&�`��ͷ|��1�j/���]�J|��[i̋�}�y��`��)*wgz\o���&qe�@���|������7R�|���+��$��Ʈ0D�4s�U��a���a��1��>���L�,���������%X}깔v�-fΕF)��a+Y\�&fl^�ޥ�Nt�5D�ikp��� ,F�a��G�Hp h?W\�ԺҧD��f�8R [I���cgC�"�ϩ�xmJ��pZ���0�g�?|��>�Ӏ~в�
~��V��_���~`�]��RR��&�u�TRtsr��|n`�r�Ԇ��*eY#��A� �yp��+��[/�|`��
�,����l�=���`o��}}[.B�Aw�Y��F�i5�!M]��?�Y�jZw}^v�x�~7�+�(K�3��� f�~�Ƀ9����z�{��z���qՐ����fx��X"��o"�g5�	D�55O��y8����m��N�G�c�Ηn��)���w\G ���_�ɍ0�%��{˓J�����]�\*Ya	�6x���7�.�?�@�X[��y�����TOg_X>���C�#��r��\
e����%M��ݫ����qy{g�K�q���.��Ѵ
����M��K6혡�܂���<�q��No����SwŞ�6��	��Q�����{�X��w�/ų�pKF�zE8�a�}�#������?ڹu=/�}�HQ�3�.�9 Zr!Qj&,�F��T_�*V���X���97�����,CP�"�M8	�>NwX�񑘖��LZ�E�E�G��OL^��~��9 {Og�5M:�-�J���]?��C"��G����[[�ϥf�\�L?�}�\4c��D�83�$]6f�&�����d���u��3�І`�a^�mWԩxҐ5_���6|-����D?�
����� |ʩI<�HE��
�V�=���9�66��/��8-a��_��{ �r��ίU�#l1�p�O}[�<m���vˑ�]��^�;Ƃx-�D���l�o��-��<5c�Uq�i�2�r�Jo���.t�P��T�`-���B�3�?����/l>��@�����m��a|���
�7.0�=��b�KLp
�M���R��L񄍐>`�?���`_��	;ҤZ�:Y��%{@�Z����G�O�K�y(؆8��X��	4?.�r�}/2F��?X	mZ6i�	C��������D��n�[^ݠ��Y�� \��njVpR���ݨ�zA��0@�b�.FJ�7�
_��/z�7߶4H0��*I��6�ӊ"�][~'ԑ_�	�-[�)5h�y:+<*R�:4]�Whvڼ����f��KzJZ��8���["���0��E�`���"ۏCp���:�dl�vK�3&>G�L�K�v�]�Wi"�����c��tn��QT%@�t�{l���Dߧ�hDm��D"�A`�������O�*+6�|��7� �gz$#X@H��.Z�: #��A���G�OͰk�u���dȸ.��+V!���\�� -�
�i��8IP�8B��m73��G�$l@�yU�PA�4�➮���G����r��w��s���@K����0f���~���@+&�uB�7�L���ѯ�BM�w�k����{��O��2]�:�:�1߂[>��W��>�(Y.�
��{[�X����RJP�}���w ��r#B�SwpI�jY���t�wt��1|-` �p_���쒒����#�>>���6��¿4��|� ��(�bI�0��
�<N��԰8��hZ	��n,�� �"a�y���p.)t�d0��':� ykX�+ȇ�Ś�%��~��X*����.�L1�+V���V}Y��{�S��㔱k��*'v�P��~V�Abd�_���8�0�kr��Ho�z�KВ�-��V���H�)��x��z89'�kj�1t>�
���!�Vf�~���}����0�/|u���q�r��AT҂%�����V;!.vVX*�Q�#��r�ZY����j�è�Gfz��`��>��ȗ������M��}e���ჷ6�^�X�� ��84\�R�Ϟ�e�����և�m#��p0���N�D��l{��,�}�mAk�@sh��&D���c�=U�4�T�T"'V��RW6P5 �{�}u�>.5�;D]���[AC~�j���J�]����D_��zt����GC�RԄH��:7���=��v���gsƿ���a|�T;1�B{�W�Ki��E�Aatkt'�����$ʵ���U��#D]�#��$��Y��!�>�x��#�~��\���e�r��7���&�6��zfR��9�H�ueHo��ڈ�P@�Kg�y��|)]���7_,+��=ӲuD�����~3Pv>�UD%��Z���2���ʩ{an�}z�Yq�(**c�^���d{�d�d���)Hpݦ����h�X�a�]�����lTI�v��?M[F&R��;:z�����nN��7����]Q�y�y{Q�����Ȉ\G���)�Lt����'DD�M�:�vD9r:&SV<-[0���[Z�W���Bu�>�*�Wa�8a�5=ܮO	��R����I]�Q9���61���B��	��Ǐ.��-�:.u���&�z�X�[��a����Q�U���kӓ�e�<1�|kV����P^�a|e���ipVo�R_<dż�1B:�3P��^_��<
�P`��S������K�^��	~���_IT+�TO�U������E�~��10�#��U� �v����R��&F��<@������c�u�������+?�R�o�zF��)FP��vp!����$zT��Zw�~c��WO�t����n�^���48�R����z�!`���&̔���Ña�zͻ���זv�J*?`w����9D����.���`�A�a�ze�������+�K2i��c�⡵��fd�1;$˨�=��Y�ea	�����ח�����7"��Ig��"��O����_��Sox-�[�
��=FF����;>}T�o���$Nλ\fձO����`ܘ1�F��K<�g�y��Mh�Y�	�= lr�Ι�$�t��9I�7��r���k�>B��8&�j���J���Zߌ�*�x�T7d�8+25=w�Ʀ�oJ	3&�O�OКR��8�D�G�J�O4�>�W�Z��B YR�����6W�2au��R�Yi��?��Z��¯�����B�1"tWE0���tm������O��)��)%X�vM)�ޫ�pHFJLs���	�cD~/�����<�7m~Ç�		x��J�J�E˜�(}�g����lڡ�S�U��\{=�1a8`�?g�D��z�v���R /m�fh�
kV'V��̈�.U�$�K����}o����������VAHT��v�o��9�F`ȳ]��:�%hqQZQ�z�D�E2D�����Ð�$�]��?R��<Ty�b'�)iE�?��+����|h�������Ξ��_��W��ǂ��z���dE�����@^=~~�F݋�l���K�6sYc1��a�w�|\EZNn���ֱ�}� �X>� /u	�
vՖ*X��p�]��fe�,��(�	��yQ�_��[��
}σΐ�����f�7�w�!7	������&
X��![�N[�y���,�D��t>�9���	�p�O�f�U� $��@N�UVo)�tt0~d���)�X�ޤ�8���L�EȮ�����Y�[�C��	��3܆r?P�M+�L�]�ق^]�E*X	U�B��JQD� �g�/�aI)i
[�M�M��GؼX0�B��d��W� #e�`��"lC�&Y�0n��=SI�����@�cH���W�*VZ��[���\0��eo�Ż�I�Ei�N�p�bi�Ű1HP|"��c��2���E������$h>T�C-%"�;I�+b�k:�Iֳ�q3(>q��.�O�J�?
w�?e�r�C������i���k��>~1���R�?d�[2j�1,�]�и�ˊ�B��`"�����4���D�z?�X@��]�@Bϳvz �pDFsd�]Ȯ�0���?r���ڱ���ݟE�ƿ�h��И�'+7�Ve�5�!�@���XL�W�zo��g�b�ş�?�@�;��%���6կ?�r����p.Ͼ�6��̦�,�����"�Ս�� ���X@�I/iMAN���`eƩ��w��$b�k��k�[�^zm�(�W-��Mȕ%��1��� ������L��q���|���v����D�|���!�����-mPnٝ���__��@%����v�'j�R��qzcj�*��Q���b6JC��?3���{�����HQ,��t�M�	'yc}s��)m�ɣQ�r�� ����Г�e�hwd3ev��7�;��ӹ�~g�N�$��|���l��](=�?���t����}�ț���"C
�γ���1�v��< JO�c��i��l���.��k���	�1�
��]�.��(+���Si�����О�z&�s��C��G��s3��3
�$=�U2X�b���Ė�BH��*7J@�����;�/�n�����E2�����V�J���M��Ȯ�G�Au�V4ׄ���meb2������ZGZ�(=� S�٪(��Q�.���VZ^��.N�I>6���K�k����ނ��ZY]�n�o1mIuù"�к�Vsa�F�����4�Pb��W��W�`]��2�hdF"�KM��6�h�����2}���B�С��<�q=�|q�F#QrTz!�hapyG:�&}T}:�|�űyR�+`%��@�H�?y���@iM0���¥�Mz۷Yg��!~؉c���ج��]��F�'KL�5���S�L�?t�m���o�Ҍ �|�U�[k=N����f�)�lq����{����x��y��B@���~KY>
PT���'�Y��K.�t"T���5�&7�G�� ����H.��%��}U���'�d�$./�,�7Fպ_�FX5���*��|	��V�F�3;Z$��)C�c�Ur�֛����j�Y:��C���c���y��/~&����+���2䀇�%KWGl+�p��
������q�i��x�
wE<�fM��D�n�c�{O�n������cL�r��jǰ`8SX�rn��|�XY3;�(0���s`��}YW'��h�z�3!i��0�S��m�*Jv�Q�U��8h��E�\�Pl�H�Iȍ'P�3�s��%�9�%�7Nj��5���MT����+n��i�(���W�v������|N��3DJ���y�+��;�N��R,�2�aH��V0'������#o\�i	h�`_\38�	�&Н�a_�K˄°s��9�ì�f�;���'q�X�$n��Cؾ,) bo�b'[�iǽ��t*��62h��7��Q����`�F��,DP֐��(@�m]����9=�n�v���B�É��z�@��=ٰ�ީ/5 Z�ƶ���v�M�0���ᧁSq�'1�9�*mT���n�7���\�:��Z�D��,l_m0`�t���1�)����k#v� 0d�q��Y��0�-W�QT�=��u���n�F�#�.Fo?��(�͍K�l�C�S�0�?�5-bos�MO� ��ʿ]�h����6�J�Ү4ګ��ގ`1ܼG:b�X(�Wz������!#K'�h�K6*Qa�l�*�6/X��X
Xk��+hR}�8��qVx�e�`h>�!��Q���ܩW�nW��GїО!� �葙\�@]u���Qf:�;.l��$JT@f~a�A)��?�n�����^%;PJ�o�=����v��7+JS���ysώ��ƴ�q��[�rd6��1ө§`x�a��n�4[QE��[;\�I�1��%�o�R+�7�rz�d�$Z�}� A?�Ca���N�������F�`Q���7q��t���ۢxJЋ��"�U��1x�ȴ+��i�[�t��d?�d�f\��B��w��$_9	�2SĮ\HV��SA�mHL�]K ��g�>���E�n�qb��U����Y���X�%�o��fH��q�����~���1v�ţZNG$����(l��)�"na؝�#�l�1j���(�_g]K��sl��vpZ��R�ҨUR��")�R���*�47��X��P��x�~W�7�����A�>�m��a&��Ủ*�z�Q1�8�0���8,�Z��-��;|�Z��o��WK��f�Q����\�������<k@��g��}C9�?��`�MH+nu�	�{��r��F9�{�;At���7�d�SoC/�~���,q��1Hie��]e�����Wg�qm�Ps{%i|������|�v���V�v;������q�1�ԫ0���:�j����*`.칢��F\v(+�_r�n���Ɩ��Ί�R�a�?6;�蟭e�N��ɚ �@w5��NU�z��bZ��A��ụ�1`Vj9�1^򪒄�Xo���60�e�_�H����<�"���ʟek���yU{wpid� ���KZ�i��]�����0U�a�����fmBW'�X�������d����GIh;��f+�ɟ�ӽ�,��z�y�$^��*��>
FB��/�|AEF����S_�Z( }L�~m�Q�m��&���~v]>9���S9hz�u?���S�+r4���e����D6MZ�g�ͪT�3ա�����[d�]�Y�S"�/���`	� �8xތv�=�I���#L�PHE���	�{K0�e�ٮZ��5��CP���<�3���A��jQnM�ji1>Rʳ
��+>���S���,�J�e��@�z�G&�6Yzb������;�p�Ʉ�9y�##Jy�j�eC�hP 9hWs� ��0+*azsވB��,�4�����U`�k	7��<�'7�5�)����V�h�ﾊ������@G��3r_�T�=bK�ZF����jWׇ��lW5�[�t��<а��鏺2O�D_�O�aZ
˒O���`!*9�^D��	Y�-XG�;��f������E���w� %��$����z���~^�́��\՝����@;W�@���W�=�?�h_O(9^`v���A\2�2��7�	�j0L�JHE�Ax�C�g�i]�@�-6�'hh�����~�8�7:,!�{�%`m���U7L丗/O'�)��wF;Fyb+��&L��M�_N�&SB��+��&!���=����Z�1�CȏsR�x�����Ou�£�}�Ȯ�!	�l|����w�H�����DN���B�JL���7ƌ�А)&��?����KE&�7/���Ub>iE�>
�a=��[.�;m�I�E2zL� !V������ƿx�3��}�u�N�Ó��T�H�Z��(����+I�YFU�F�
.P_�ںf�@wE�v��օ�HdM�ˌ��ڧ�\<�y]lƛ�t�"��W[ȗ0�0�f��.�J� `���+<Ʋ�g��b?�.�aMӧ���9V
�Y�V�b�Ws�lKGzWb��&�^�?�s��JD������l����!�)`[�<�J#A��5������7�1@�.dRB.9_M�I�h_�\�_��iTnԔ��9�5�M��>*�f�:���p�}-�!h�pc�E=�t?tr��p15�����Sg������@  ��$뎛A����#d<u����P\s�];Ё|��{��#dL��ʑ���f�k:���:B���4�����(�xDX�a�'[�*�������:~`�L�)�uG�gVݸ�B�?LL���oj����U8�\G�,D�x��~��е���K;����UO��7�L�6��Y�x	��ML�#�0h�O����~|;�W�y0� �sY�^��
H CE�}�* F�lw���ӷc���9���xr׏#��'?��,�{�D��.<�P�ׇ�C�)|YN�I�M�!t|܏F���mK���rJ1�h#[�i��V0�@C$�XQ{|ҌLu��Y�����ټ����	R�T��[k�i�&��VV��O\4E�nXVnF��!�'�/�H.E������pN���ب��uZ�\Y*ѱSH��(�D��1٭N���y��&f�{¥�P=V�퀼�jVZ��\��);0�pwU�"~��KC�$%X�:Ғ�bj�e'��v�H�u�C5��_�e��+c�Pڇr�om�iN�-�������t�3�gk(�����V�۱�&�I���S���/M�4L���V9��]�;`� �Nb3����0���`|-����|v>���`��x��]a����X�����+X�`rY���UO��;��K�B(���\���];Z�)�<�Z�J*�V�	8M�ҙ��:������ZM~%�[��V�V�dǾ���ou���,N|Q�O(�>����	I[��>
�0����m��b�����{���<8�<�\/���45����Y+e1W��}�u�%*v�W�w�3�<��CX(0�����I���\������E$�M�6z��~PqW�>�e	L�Ls,�8S�|�$,��A��]���>��\v/z����R�0���f.k���*I��a��XK����N�gk�u`h���