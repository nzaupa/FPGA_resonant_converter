-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AWaSu1T2nhjtR0wdOEI5J7JtPYrJo6LtSxW+2RgwBqsdpgu6iDiJMv2RvFxY2HE/b3shqk8hBRhj
RgaxAlbbIjVDUJKHF+AmBeZZd7P0KM2yjyRtbzotv59lo6wYFynheDSoVqKKZEdoKWd+rrNNZlf0
EBWrjeQErZotwbfFiJaSm7ZxDC8foWg/b1VRg6ImtZZvl3QLpsdWWCixGcFh4kFQq6yIWvrf06zX
l6Rp8jOKtvEuGRXzGhblWdeaVr4ZGATwYOh25vanoZ06ldNKioQcTcdbhNbQ33hnrMX3CmVrJxUW
1/zrz7LRX7AMt9PtXB789KR0XI4hscPGyyz2Aw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5328)
`protect data_block
IJRJr2smxd5rDsrHRN5I28RzGfiZiXWYGU+aDu45/ky87n6yy0S3dGMFmMa1Kj+M6eTTLJd93nqh
bHCIZ6Q5JKcUboJakMueKcUBQjw4zMkp5mplPSSWdDhwKFOU3JkTIW5nHi19+ne3otQw7Ea15a/o
JM3Q60K3lo54US3eXPuWITTCtCl8Z4FMITTxEsXaNe/TXNs1XxyTJ0rps9t6O3O/V3chGKJVn4ed
pyDsbuPTNwKd/9xNLmVGcnugGTSm0+anVydoyUI7LI3jNsxQ8CDoALn2TiQwPaVHMHrkiGLPfGwt
lUlwuSH9irHMYVFMN2aTxEtyKHNvjTyw6nq89el6e1NCnFnDnTx0A5IQydSnVoIiFhdTX/pArTfY
WkCTHCcKH/5bCKH2A+1rO2k4TPwrupHD6xTJnmF28uVMFzW74QIo7dX9VoOUzI52k1LXLHLnpoFb
JAeVKZXlqPxYTnctPVTH4nl71V+k0/Y3OvCdoYz03I8mMZDQK6BepoXnNOrUzdWJEFkbyoqv7k6b
lK6HGd+RgklMbq1TNwLmw04YFG3S1ReB44RuuIxDgWpTdW3GELPsZUfbIOIFt1SssrcFo2TSTeMA
xSMhGhauDwc4avuPeS9rjyhta3tlJhirTmzrcACPndM9BW7TgWmS3auSY8GRyi6G3Wao9HrjbsXj
OaAdG1h2VyKgBtHbQHbIqvPI23D/3EXTEQKTRy7GaFIIp9a0w5urlqXm/cjzpfxZej90aDb69Q8i
8JIm9VdvCB/OWwxNId/y+0/LfV+rSElFX3AA4T/kYcvRBfmX9gqWiW8pzMdM9Y4RNt/ywsTmr76U
MSmSKEqq0f8oCP956Bb/TVXIGfMN3lN+ZM/0h0iNW5Uv0WP2K3Vkvw2MziNGOq7aaumnatKgjc3x
lIldBHdivAyoVZ3HGHPr5V5I3x8VeSlSIHili08DQ0rP4pz8Q2kbrDFjpMTMPaTUdYIKacCWjSkO
YbVzLeAjhw4tVAG4cad4jjjUlFELXJ/Kj5ix5N3k0MQamOs2bDPs6UsNRwV/YOIUwiuRMI87eWYT
K05vjCRXTAMCsoIoLJCVWyCKjwTcUXhxAIPF027PfQ7G2w8IP7cMefU/W3CuWgJY2VABIPLCNjp/
gZ1+qnfmiNw81KcU/nnUzj6uF0rp90+10dgKrQarRb2a++CO3FwOqYVEyFr3cYwGWQr/MC1SPTVV
0sjhVoQNBMQN6i11/u8GVaijANzhGgAb+ZTd4bKRijsbfQG/+6HCpDO6awK1Nv+U2KpZiJAV8pd4
COum8VwUwsoV8al26sNnoWWmSdeLQADznsbhxvgPom2aqiQVw/dxXQjGKO7awGSgZBQtbRZVP3L9
KfB7FBrnZkeYXyylrM9biroYUeKPXWsaEGT9bV3erQEDvM5C7x8pfwCwSbFJXinlgUUAG4CMv4To
OKtTv0HMxSEwRC7Ns93GZzGfsWGVGRJFygZ5/IZxWNfZiu1F4PIVf/qnU+HCIyO2qQeBr8Q4xqmZ
UBWBN6pJgnVy90LzoHqvPveQf1v3pTU0ymK+2+VfjO38a/EMM5rdl3mhtuspNe3Chqizgi0A1IyO
g2wLkKVE7+Y4CQqY+yqm1UY5N+9/alfxHEFbBs/FsWAoQxknmOliH1ifDXNDPfOmnjrVKMm49GKE
srJKDsK2mYbp0ANovJ4LDk3QBix9EH1bVaSim45hXVTz6cwiZF9HPptnk8ApBmNetDOKjG245Wjr
Sp8F5Z8uQmKN/HQ4WJzAqB5wDMLLS1wgr5PDUE7SpFl3WSCeIPRwpCaIMJxdlJTqw6FPZqvP/BGz
+mh3qii5rV+ecuQ1+9aLDCqUO0Ax/Mmg5Bs1VN2vCvad52GLQ0sRfXexV6Hr2tNy0PQGNsUI+Tvr
Jn0aiwv+/0JMY9z+4rJrrxlK4uru4sPVXtFiWl/5FS1fOIm+4F9wcfro1tMMDVT3BRiiQ4+/c6Me
g6HqXk3kOLhz0rUQh+/zqOLxMsIjqfyLrWzim8FejLqrdrvHGwR/Yswe6g61Tad1IPYsP3nWTjer
Rzm0/lNMBSJH6Q50modgu5ObMVgO9/WLbDduSfEuP8iSRdZcmJ/QLkUe59V3IQ6quDV1sgbZvoea
OX/oYjvmvKILdU5jn3x763D6pLQSx7RxyL2yiZ1h/8ZQ8bjZlYYn2nER4D00hREnJE2+lK4FgEoi
q3e598+yHp+HsjHpwM/DabCG/EG2DWVII6pCLCp6EwP0YTVcguqwAQeRNtLiLEUwaJsj1MqW/7xM
pDofb/azejS+PyEmPpskeclZsMvFZIpl0iLyd7LPYKRuSOoUUpGbIYM5rr5b31xHH7kray0VE+PT
dGRiHNHTgIfQOwHDujZlLyYFz0P8/hxJHw91jDcYzO7eMM5zgZ4qbfPkH/O5J0701Cy6PWIcvx7B
gPH4krngzsNpPn1x36GzCQ9pvw1IG23kKtxBillmq0MQpx4i287h96KdbsdJkNZcMgJmDgezHM9R
1bR0KF0RGxRxepDme1eaAVqSskT5In0cAH2nysBEzFgLxqDLFG2W+F5cz9trdTZxZhpuFVNLzmO8
W0S5sJIe+PvC6LNiMdyLCtS8Uh8kG1bCW+IiVFeNut6nDLSig8wB/PwX5YJu/Q38hu0khncIopxn
DhY4JZ0sM1nO0Nd20pYAMdrFyIqBA3QzuBF7SCRbVYV9iN9+IOHkS98ijBP4u+zj1+ZaYzDuWAvX
IFq/JLAe/htP4uxqzmQwsGzqsuOFKLh8O5V3xnFIFkl8hYaKgulIvUYh9FV67ygTDcAUWfdnW1Ck
t9fEd85SDPTw4YB5FTbCWa+/LlpfK6w1vmC31XuLIJDDUCc7H7T88ayBPXHiCSLwtfRBbZqBhafK
BNpXR5NOPi42Gh59aPGRejLs+Q5d+9UHhSnhYWCs1cgpjKQt3Er2ScEzqtKWW381gMOYwyLXbT7H
mx+dfxjc8+XdTbiMdUmRZjsdg2HeqYtzCJOZWILpDlWyVWwZBC4NdW+R14M0LKD7L/xY+KfH37gW
rg0HmffkpLdzus4m/txmjqWu6j012X3ORxxNH6M554DObivyWdrLDuicsaKM2nq0eGTIE6oYUCE/
+NjET9bB9Y9AqZ4uDpvlMNENxOFGQkzeaA11dv7mG95C3A4taJV+ZNHhvoXqfvGJ/M0Ps3fhVIG/
Y4J2/9BDI41kZrghb+cLLtoZgV1u/hm5ZHAYW+oCvqdZ5nLWp2ZOn4mkJkfgUQCkAIqIvy/IigSY
xW0oreAB92AeOMjDF3vryO/12YUF3widMfLWH1HYrrGCzSj7QHoZLov44BHsEkzUy7p/pwtLo1BX
BtLrU6VAlwOQYUQ6ii4zoGW1RtuiK4xhUxX6PmB2F6t/pERNNppB9bLWgqynKalGwibhj2Ztj9Pj
ot5CeM7GTnCHIXca2BK5CHxQnivUVOdDpbueNITR5NqitZuexArww+FzUDYHFfDzfrtVw5Ge7G2G
jLC1ZaQEER2toGfSE4pJXaPJT7RfSf8evFB8ncIGsJ5tyupCnpk4Arrrae47SwS91gFJxUJKhdIV
IupCGUJuXTvemgo9zrw4VfAQCPCMfoVlHTnvFa3Y4L+VxYDAtDmuGRq4NL9AFp1lGyqipIiUt1W5
qmSJ/JgehUedpagMyZ+rSv+BUj+2xUfeUfeDbWDDxaLC+9nT6E+ErTLFA3LFqdwDuautc5J+myV4
iM+3Uhhrr4bmTxukPm4bKUaz5gLaF2gmcAc/X+VhRsN5a0QxNIooGEe3/gn4at8XC/+mNff4C+zZ
scuu5Z6JivfuIWj26e0tMTekixdGYr20+0Iu8zXYga/REcK+f55KIisC37AyJcD1fPBc+reKg+fF
ZSI/JGmFqgYAiOptubNvg3UjfIn6X1melUpzaUCqMzq2xMiSs9TyMov3Oa33w5thhoyKzjy0lugk
8XYo2F51enyF/X2Dr8CtXMGwADCRfgRZNgEMIb5av/yeAVAZRcQbS+p6B5nbEJRMzm0ULHLu0OG+
2FDPQVVkBJ7MGUr98a7W09rYClBXTXi3z/5tix14zkzrz/IRleamF7KbNNJj/i2lLyxpDPTNb6Jn
HuW33Is4bGC/fpzqh3jrhpJHNX8TBU1ZbjSHn5OFjFKepONlCqX6ePu6tSB9UFZIQXpv+Wo+GWeV
67lfGfMou0oIxDdDcYFKnTLh5C2MNqmsHhBdFfNvBZK+wU5HPIDQ6OpDA2YYEI1+ZEH+cjoI3Azg
bMcZgz3HcRDLXsRuON6VefR4B+SpjCCpF1WKtktNa8Ztklukm/CLEYV+pwBxacItI2XArKv+PtHr
yqleNLuTZ2EGST8l/80HaixFsNPxTI0M2ndR2WeL+cSW58CQSp+dXBZ+Mbsr+1cswSrEDT5mmspY
mJQ35IY2lO2ilDD3oME6jcBWnTFMtq+2C0P4sd28qWYX0M6yQnJzmvkJ6Xo4nOI4w74LkUApi9p8
8hmqXOZJkias9feHg1t4duB/JW4z/ZDrWsTtgY8sFUo+A+g6aYBq7IFlo+5u9OF7EeS9VXOby5vB
F9gkVbcS9wGzBtVmHNZHPdn1QUXBeJfIhs8RTNSkNnGguH7wGB5WMVtbcmpqAyxE2CvempM8li0X
g45M6ZtvqN39WgcNjRt+67iq86ZryMUsSOo5JlsFjnOfS2IP/yHZt7likhA8aiZAhKdEHGQCt331
zXvRchBEmj7t0Zz+rFNDcvHcwPUjCKcUEW7zEWOY2KkGuhG0DmO3E7MHEand785BVsKQc9S0xxvx
ZDBQrRkEiEXXr07RB4lahKmICO0w/AEDRkOUwsVFb/MtJQ7THnicR8GPCNDZYT+kohBhvFRUDDVc
w9sdt9zsYZdJ4g+03A+p1eK3jhgtllKr4xq0S/49b+XcV3lqfsbablHB7hA59KCemNgtC82bjxDO
rXPvLmZUpLK5SK+axuPsjIe0VQLE4GPvh3zGmwJPF1DsyK8Rx/Ws2zlo52gu5c+6cWFZwmmRlCyZ
u1bFCgVE0BcLKH24Ct4Okz2+kcVL19dWIjPgIu0bqeFq0+MBI9VBDHmj7VS0hxXn4jPyQjZeJVMo
dww0fZGV0neZBgkIFoE3o6cHFQZaA4eZUFPHsIZA6NxN+AxJfhMvAsBPsMzzUnwbHWlUUsIb1aSv
Sd5rIottyvLyZ2V1E+tDnql2G96LtNqcZ+4mFAIo9pLPxw8PGqDpH32tmQiCdH1eQ6Jr+ChKmKGX
IlhPSEyD43RnoSf2H3Bkrf+LL9FSOauQag0aFLQFlr5UwAwlV35H8yzswPK1Qn+OCKMbS8i6Z1wv
BAvwW918TWZ/vTO2ZLRnSQ8shKLD1LEDt7XuMIqt6qhc4JzA6errmtrQillmDbG6+lWY+tUP33bs
6KeSeN1tzGVolrBj1xR31Z/+sThLYPTWnbW0QjtSCtramwVKpVDGr39ytH5zpcetJrUlglNfj6y8
q9+uttViFwKJxpRkS35PFsxG/f3yZL+bw16OnnLFPKv/E+GkeOD/sWvG9YytUaSMyhj2+Vno1meU
87UjMd+WvwqdiMrqKKL5Tm2AfHghUFpY3b+5skNvxMLKqVOydJQsVKQLcROWY8bJ1+pZbo9fqa40
dy0rJ6cufgaWAVAw8SLlOxjNVGKltST8s8sEcsNRKHWd+chFF3VEOO7/gHx+cP9ahAH/e9eaOde0
6kSJP+qGRkUsgFZT1y1rsBWHlVsqoMhxavFHpiXa1usKd9qtFvLaGbtgaLZ4L4Wzokh+T8Y3twCM
m9I4wuOPWk0uvb83O9s+GNE+tRMxwutdzYwm28WGGPJlRbt7Qp9Iv6RvqAAOl+eN2TghA/hCIIZ+
2Q0ppInSkQz83oScP4Q6k4yVzQRXmsRwACp7enTJk6azwa1+30C4SqCkmO5D+MOpe+MZQ6PLY0C0
PL3c7r1EctBD4CmwmlHiRdhyjYegM0fgYutJYuu7jAu+h5KEbnfiSQDk3TjFBKEprOiKWK9otX7m
Fys0NhPB0YJxL5WLL2cXKP8FX0JBiD6JxX62Nw3r6r96iVvu42bJ3M5S65IZiQsTiSkZ3aq6wpYy
vCLpKi36j6nT19O2euX1z9NJ5zq4pMakYitn5b7oc2QYYa9Cf6efLPuCsIxsJ0tDHCUDQ1zC2M4V
y9lzr+9+EOUmRV2N0NYYflzwHvPv0RJybwjJCF5c/6tJZwm1bChIh6BGEqK8QcaJAPGa4QjPRocn
s12fRJMtstdKjAAgamSgqX7kFizFZ4nzVSydhGfowvZxwZaliDGwQPfI9Xw6vIcY2lwYB7dPQMTQ
hYDa5P33cIvzI1Tx4T8hBrmedjeO5vGCb9TOFxh5vPu5q0VsUp9dr8o6xVVWCnEEc8ljmXx6uyTW
LZKsxVJvxILjuWn4Tg6kOrOZJmSWS4zl/uTnZfaqdaJIHDo/oP/uRTBMimKOKGaiL4cSrA8FOD3q
7nCqhBZaAlbbXMHYObrSO/3biTkVFVmDBeyvF1dJCWcOrLlm1goGwstbwmOt/QeY76kqTVZrhwRJ
Y7AYvisQi+BrxDeXRLvvqn5Q1sH4tou6REceGoTa58uRW8OfkWhMf4Tx38IlPM0hssisj5hKxUbD
57+x41yeO4Zf31Yd6cwfNIFRkpe2IKThIs3XLt6A6XLrCojWYvV8tO6SWx5f0wsB3/isc96D8sFd
hGh55squify5GW+dysTQZUQr91fjbs+/oeBE0BL8eh6JriHMJWEWrwHjxW4XO5n7QdtsgpDC0qnZ
w+FaJLMdBbAGeTFWWYCgyY/ggJAUkZOAQAC71WRNP46j+OZ0/1Ky6lida0KRQIpA2tFpSQSoOE/E
JKm26/uvZJM5Gi4G+5LUVCUb1yWvu6EZmdNMOUByPHMU6fju8xka5L8yj6dFTMvOTX6fMMx4lc5C
z9XDvxsJ5ZV60KQCaXQHXQe0CwGz33M6E8AHKMrRw0fAOIox5+P1DME4919KD2fX+qT+sOblQ+ws
t1yIBgrQDh9OaWsWccSd7z6jhCkaQv+TeBVloHVd03Wq1v5ZmH3JKi4vngKu2UNx+Cy1DMB8HdwY
UeStJAoUmoLUXWhlWBQBBsfOZWmn3R6lJ1aY
`protect end_protected
