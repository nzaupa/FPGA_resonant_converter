// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
AASkGnlK6aZBgeowr72ucGupkGDhqb/51wYIf3LH2aheuoPL07i1F5dprnoxfEgCnIrwym37Ofac
49gnkaCa+xSik2BmHdhN7QFrmZZFtEquqmLHN4kUC0G3kO8qaWCd1hEL6IeM54CnBg2wixaRVx46
d+O65a7spLRxSMoL/eaMYXc9XSZfRDDaNBCiS6/9E63MH/6vur5Y3q8detylBshNxtjgtL9TFkw1
IjCcdMIcJ8i2gI/UPZscycP0Io7ft9Jl+L6j6JGLZJwvgmGXtqoif7PyPrCjY2NS1MI4M5X+1UXA
5YpItalY+KTA5i0b/c5goRoGQBYYKavyDdQWww==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2960)
IJEHYVkjtuQBhsn633ov+HzjnEEUlq2KwebtVpRBer+SmFKKsBiyelAl3Fs+i+h8dMbe1er8yJov
lByz3K+A2ihkjR2sfbIXxzuxtO6NyVnCZjEnOoP8hkDczj9xMiZ6mCmOLiKhqSP2ON3aa1DQhasG
KOzStrfKNePM+nKJkJz43GI6XNPKDreBfXpLUrGg3NgPfZaSTb11KBL2icjjCRhtSoF/kLs07TzT
tbNdVA7hubO6Y2pfkOV+qH0RnGbblzoQ6S/l9Bq7p3qTsEkcJQ2MNuQ9yrf1KQDD04eNs95LTbKF
OZmY+T+ewefT/Yi+sBdB6kXSKFtkSrvsm7M5+yrv04+J3219QjhQMQmURvlCsNBzHP3C15b/JTFs
6ZPk2eSRyY32nFiByhiR7t7D0k9/fFZLOwvSUq4lhjnre65uesWXbgqV5FZIWhCFEOxBE6X93NuB
4JlM8hCu0/HPvbY0AIrVAnGKLdlMbv9sFGvGLqTON1MLa1ievwkcNWzgYCSUDueyKXWx0WJ2by3T
N7dL4S47vuAh/goi6lhiWcvVFZi8ue3dznew/90ZzfykQW/Qr3xDDx6BYO8FCnbQB25Ibibu9fb6
fu86zdFtOaPdoqJ3M2OELFVq+TjCjVGOir6BljE7kp//JR1/Sr6zImxc7dmFPdfRwVTbNVEXKdcX
2Aa5WZz6XZu7OHbp0KJsg3z5i1Nuv0LL89d62dVsNIzLGVA011jDK7IfLYXJlZCZjH744oiAUAs1
D17L2LRUaSz9fPHguYLLWs2YHLa6r4oNDoy7GeoSqo2+y5X015d6UWi+J5LvHX1wJcVgdCIFsZ5Z
vB7kWzjCvN6KaFJ1CQfQbqpHuvQIgy9XrIrQ6QNu3Y10PQvxxp8l5ktvcFocTz5NFqIgK3RD8Qyi
50+qYZkX6FZcDaAwukaXiceMUA9MjIxgllHT7Q00+JeD+gZy2VOpHL18HaQloNZsqtfaM1mdISfI
wcgJCIzbCpUzsCBkN0fS7k7BYVKytafM2Fy5RovAUlnIjuOWdeKl3bGw+jnG6mgtg3wNP3+HFs3x
OJ/4BZ7JVTpDu5nrsVEXKdhmImQzOGRBv7notF9ng87cEDsX5uBYuNTrRLX2arssQeoMCdzx5pFT
5ZnEdGYDTlj3eHthkFMUruhxjEuAjI31wkKwISixSo1MRkJgDK/t1tiRMY4Az46MBxmEZqMxUCYW
xLQNKjK07GM2PzVOk0KjHdH0NaJgIaQRX86ejqfIVc8vLaKqIogXDfXfVdEknojDpkXjlXfiDcwx
dZH5yWPDZrk7MYKg+9HHxSqsH1r6wzXTZ2tSA/cIvTKSj1GwSb7gFcQfzhigSncamfr33V8TPPNT
P3OBuWcoptzLIITFHKBkbw08biyaceFLLeZdtvuZtjv7F6FYI9nkbc00cABpZrWY8TCrBfszO/Ln
XF97Gl3ZpL+jf14NihWYq8o5rEG0cRL7tGF5YJ7P2L4ryLVExfxJ6S58kwgaYMXXRfWAV+rp6qRC
yvs5epQWs2jOq1mjF/sqV0GxxXx1irVpxqTC1TkKUesU32qMUBDeMx1fUICNuB3xklrfql62zOlD
mfKlb9ch6DNc2DtSNFetAsXWRYJ41fMl9PwYyYe+EHe673Sgd1dagQshXmZ8dtM9H/BSb4W+2Xs6
CMEqHXKRnqTJPjlVu6Foab7k4cm8uMmow4YakmYDPIvRVuB6E0x2WDiXC2DFKLl9LQDXQZ7oC9JI
up33XZjrNhM8Ur8oPTscWWwcAzupWauj+eWZs+MnCqbnEvobig0XDyxFSW+AAob9WCGFJXYdSzy9
+0OsiTBc3ILJVsle1NV5x5FCagsBtQNKTSyu66inl0M7ltuQm5cuskGVkWwLLzSzf3oih/tLyerG
oBUQH+ZyeqabV09nMThi0zVDoldV0LNlcdPlReC6UHwQcbt/Jaoa8STBFxaQjF8WLnY9qz8FqLMk
rUbd9SeGLZ7sSxLjYX6wDdfpgVqNh5gvFKDlk505o8u2GoReZsdo/foOB4xdLuen0BoZwhVpJTGL
bvwbE3oX2niWxZNvuCZvQTsLWnG5lRkz4mh0sPxxMyzOHUcKeGsK6gR3T5LThHTr9LCNKxlNfHcs
RDcmtWP2xz0y6zuh0PN2cnoFcG7dGZ2m6vWWE+Qb+aMziIZJd1K1ibEVFZ+kiMu0iXYOfTTHPy0i
V42AdOr3KuuTgGA29/yIV05a8QhJ/YEPMBjKiVo4tCtnbUsl1Nk3fiIH4muIZUelgDGeJ7CzzFqx
g54IwVkJwHh876gBc91u279SoKaB9AOfhDpZs8U5aLp5kbKMCl9H8w645f18mt/Li+hhoLfi+R/b
noo0TwYxbEJF43sTA9nNl817ZglsoVW798gWzcmo22AdNR8KO4XYy3n8vZqMdhOQZPayG6mdTEtA
R/iFNX9nBb6Ntaod/t1AEddAJ/PQ+9rPlHgQus2k35W/kAM+dZ4Wvix0KkS38vbOajvtN5cIU5jD
bWoSzMT27bmuOlOI34cAb5fdleoinLPh9EwgnE73jhFgOtUIDS/I+BKHuoEI3QtVSYZ+V9ivJKGH
8Nr1RAIpeOoaLZ+lKnhr+nvIW5Pkxe933pH2rpSDYUl27sS/YsDhuerEk1F61ipSnoSDHcGoRuAT
6MWGoD0yQ3pL3D/6b3FYjsZVU/4Pt2vVWqSVjb8VPmMPa7SFw0B1/7m96oEIyusuXGidOgcsdEG1
opPE+q1pFBhUEpjt9mYoE8lpJFQI9sYMHpiP82P6TvQDT1DW4LHYnWkxBV46xnUImtlXGdYD/xJv
8JNZtlmKt6t3mI3GQd33ynuOeEIOlSGVLS9zEyYQ3M4X/UykTNH2WoFgbssPUlFeXY+qm6judnQ3
TWXMGZQ+0oaPRF/tTqszUlg/1kIsS0Kq0T/oCXdK6gj29kXMEaTo+vYbh9//MFzutxj9kU/FqF+8
iAR1skCjkercIYDR1uqmB6Nk7bngaddglZ0BA2FJoTubBMoq1B301IrJSJ3WaCfyBH/Hj+7Srkq2
rg7Iwlnzy3KNkaevvCTZ60AaTgrDbs6E8wYrjIasYxyvQDEYrcP/zb5vzOunFZ2vwcWoc+Zkp6at
29FOrOH7fEYqgsK2OpW3Nbdhr/OoEAfTZRDX05TGJKv+9U2HFVhzTYIv2Sm2cizFQBr33yL+jUpU
iZ+2kB/x58zZELYAFFIMckHuXu8maHt89ztutQ9db8RCsRo5hPK8V0teZQOT9+be+prlvLgQqWiQ
Ql/5M4JbsnyDoJku7qNCwibGwBZM8eW7xfyWWZPJBr3+6PusNb91sbLJg813M/7RKNacvaLm+aUF
VoclIFVjRpfaS7tDb+GELa8+dYn3Vd7jysoJCnhxfpevNaRBYtShvzZ1ZjHgSkVTHpyvGukCSA/N
CthxG3J5ElMldncqtcmtbgFNA/UM2fLXj4Nubtdz/wQSLtPpjtLQu/kVOeRKXWYzermZGZIhYetF
UiI+U8+FBSzP0haDW6JdmiyE8zFC2oVkEQCDyYbheoXoItPbSv9zT8rscAFh8y1xdHpsFxAiGQib
6OysFN0ZJFGQVkUGK/X4oxaxnUSVm7+mgyJsgurWPv+tBKe5BoubLH4Xp4bW4OzRym6xyf9D2Xyu
ZQ+SPRybyG2VcMC58lsr5AL2Et1qPaaP4Rjw3CeSJALnbBkt4ghaG20694hcKmB6rWzajh/11Amp
vwBCuNRN+RQAn1gQIrxh0Ef3IwhndaSIESoC8azpnDbMdVdYoLCB5JjjvcYalTklk9vcO2ZR/jWV
HBuxxCHFDrIWja434Jt06lCDRC1w/e8rZFHFhiS2ZA/wVzRNsliZEx4RTZs//KfCLxglTLd8Z5uN
CtBIdirzi3wjEDLRai56JI6GE/HjPbwJ0zBs/cO5tbJS9LFJGnQmz6zv+LV4h5xtrKUiLYo=
`pragma protect end_protected
