-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IGWLwhMIxOck6AlEYB5xQrS5rxCsRJfirkRSEN2mxcqyzxVYL1nm7fFM5/zJNz2Lm045Jc/fUTvG
VYp1ia1eVzajEAJ2xkk60jwrmL/x74kDoxBMGdaFnHTrKqZubRx86NyzlGRN2OqHGiyBoz6BlFVm
2AlZMHGoCGfURTNi49P4mBECek/ZDbkoQuNeuziXjeuwNHv2u9+TE1byheZXpNFK/muXWYLW0P2D
C92zyyTIlQhEPuomi3PknMCRIJrmhI0FIIW3AuUyxdCWpW84cQWCUS4hPKedufjxHLLp1nVgEQ3W
lMM5RMYKJ7BggTp/oVCq7R4hbuUjIYWKh+IeSw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8560)
`protect data_block
wRI/keCarZ0T9WQUISshzFhZFmDPlgmGb0cV5GegRoK/XYTUGftIijwAZzZ04tJ54VggTbKjcqP7
HzXvAtWhhVDV9lWm7vBVY8f710U9u2QweHuLBWCl5+7xGWvWLxjHxL+BbA/unnNi24ecydeyfu/H
0gJ27OfD8YhfYejsTZxByJp3UtPkZvUY1MnyqZwXPxmJNk+ct9yxcQ8uC+DqopmPrhbXqV6qeOLp
zgTbWW8Dn8sP9rI5K9bll+g+Kv/SG5C6swKKXRsrXnu167BeSuSn8Z5sWhnZ/z42vP4uXDjHShhm
qIP9b+VDpAiNrBK9tbb4Cn+S7H6IxaqwL0hP0phPhZj12cBgI8Pe0PJI5FoOd/qWjs19ajZ4GgTo
zZROg0PzIZ3u2B2iX0dW8KgDpvaHVjJPvK5D1kf6ZVxQRLd6XQwqXkLF2xXFuLRht4L1XwzIgI2J
zLyqJxSAHmlGJrUSAD6bc61clVh0hRcAByAU4GuB+SypYbaSwS5oBrmCHBi/KjRVHdPRYXEAtvjL
33HCfT/QW5xljOSP/xlls5rfSBmARHg0yJzW+wXlrVYBFmAficNfKtWcWnKbEDLq3qxiJY+2wScc
aOeiZ10zPHFeZi9g+ioAHGM7TQilN45By1m+74HkRfs52N/rUp7CnGm/OcPJHQ63aE1fFUrrg10h
xh5mKfVn+HKdtqDkGIaTG0C+T1vIbD6BIeBYI0ph9MnCD38E7bKjJiaXvEwRYsabQXqLnc+CyZ54
5FMbXZ6g1OehUQLPrseog6ghFq3g+vTKGgqM+8giTqYCWBP2xkUKcbgCqZWInRz22En6aeAZzCHa
8wpUfMURtHDIo5BB8WIZA9UkbJSc99ZAFzOtwNCamXqHbce8CNWUWih6ycwZABy/7HmEu3v1Y21E
GQ2v5ng6/3gjFJCDe5x+hfe5RjkOpkeyh7TNXpjxefRvUnGkYNAnc9JbJ40597Lb9wDiEDVbvfsP
qah3kRHey4+SITpm84hchG63alAoTOSKkvDgIacjiTlVoku63yzYfd2s688Zh3hTGCPEJI0MnwcL
F2WOM5bzIjHSKqe+49yyl8NH0yZ+nIDofavNnzZ26w1xBqZx6Emu3DKVgw+S6qs64e3sVpAqPgeG
J8PIkul3R2HeC8k0757jD4TS+dDCciemdQwTUEn9Qai1AygLqdYWXh3TTJ+FjRg7EMwQnaC+Xaxa
aM9f1vfXrNjHKsvOK+M0ZlOhx4EC0JRYgb93HMd2V589HcX3gOwUD1dFImA9/Lvu0nEr+3v7LaCe
OLH5lhdxDzhXpcQdqDBpZA7v8A4PDO152ieN2aEgQXV0cD+JsjlgoJnCSLrU1ndpKUCt45sVtPHq
gjQRHfl5Nev1ytRkl16fPnYimm9cn+aWVu9ksTXtMkUk5DF4X0yXuO5X5QXmEIf4jZ63VwTukN1+
X9RHqltQoAGYGMH64qdHbFV+n3mt6XAYndWQ1Cb1pEvN9XWl6x0iFehBnQ8wXyq+KeYqxEfSisum
CM0bQQMrrotoQ17sM+ql8iwKcPdEsdgy1Y5WMkKNmVeBMpi0oz4jHVBf2ll6toOnlqzr1QSK17bY
ClvW+FQlo/Plf55w+Tdl8tlk7Q/wtzcto42so47eWM0K+YMf/EzGw0hlQJMwGDQMS477czdysubB
TkGDZqfwHWz/Ps0t26MT5YbAR8QzznXx7rGQDU7rXlH19IJGHE6urNzDhQGkHUeo9ceeqnbMWvk3
eIKHUMsCFugkCDgOVoq0ISwuyiADwk1Uv54dsHmun/ZZ0TG9n/9y/26OLm/pzWL79fNOd4w8tlEQ
hSODLjO8VMPNi1mtx/BdtevOsE6oyCmptXrH8dAu36/X8MqRqhedMqlcMAFWNicWSITrU8oxrZPE
hpvfZH1arbOf3Kadao6IR0BccNrFkGiXrjD35bKFZoYrECOC+iGv57ToOxZuGcvB1Pb3A4SIKE2j
ZV5wnu1vbo0TDKUPjxLWp/hZ3epnjo5JYNwlxKIO9QLmS3qWqjXOkSJ8677hkGffzwVG3qkAxhAi
6MItcQO/HechgBqNLDflAr1WUMHaTtpUNTOdCtbDH81s+MoCPMJgpvw74jMx8OQSGlyqWmqSvckt
1jCovx6UnlgPddMe1ryFN+oCTHCNUoW7H2PcA1WflwwqXG2XcFqB/p7wffYdhziHevPViAv9f9QE
iNdFcPh50FmafV7Tgg8LabRnlgnrKs4RrnPe+ZjxUYg32G3aKJjv1MKb3FjSSn7Rk0XaRER9mMQ2
h+URXhFrqL24WtFmUkbGOoAO8a0CKFcr1wFmlruPuWa5da7+btbosLVTgJ3pVEvQXRB0W3LSktNR
2Q032S/l4JfoIg32ziGx/+kYl0/9/tvFodaBLxRZQVNxuIWrmUzR1GPkSH+4dwLGFf+Li6Op73ll
c/3pFLH7ufBCARlcZdlSrHOtE4UsOCqOsYaU0O3YLmlb5X540ZA9igvHsw5WhTiwvrlncrqvrqbM
KxRz0Qx+jzAhZ1iz0aNprfYk9rOZ2FCNk4JGvn6vG9qj1/YT5T3mdM/pI9HiF9lwyrzH4C/pMbgw
ZL18dV86hO0MTYrISbbLPsAkqDI1SJXKeE4lN5lVmuI6lM7SEIGu1N+VqRHsrJyMg1S7oP79mzGI
p7s5SnEkVp0BUesvxpITurvmtsJatiG9YMFEXK22dL9+nV1PjoBfxo51682zbp+Eu/P+EiA5+PAa
fezpQ9AwpkKfOgH9HdMleM5NpMJwB9oOwkWHaqNrsQcCVsqZMrCDlMEW4URbV2t1IJvgE6gkHMf+
+rwjwMn2LmnJOTFMuahAUnLoYp8H/Wjk8tBcm/n9cwe+2d1/+lSyXLN7Bh7p2Zy1cO7ZeQyojhHO
CEGkdr8YayRprsTtZVHPFK3iaKSQSI8KZAe+hBbBZnVZ4AxBXSC27QBfHz4MOfMlqvgaidlp3PKS
YGqM3hxochdGn0gWQT+Uliw91bL8xTQ75TIq+aBiiw2AiYfT9wmtiL0wPBPkBcU92fjx0STH1gMe
5HNOuxH0iDh7oW1Oq4XdMxzPQotSYeNb+7Yes2v4Kb/5c1iaF2a5ZwrfLxa8PQRGkmg7MUbSee/a
DltlMnbQjvkoh9mHuAXPnUsA0bmupIrgPh5ihrH4ie6oP8r6CYNfdtu4yiA0xQc6vnQEM6axA+Gp
m7CLwIx8ipsUAAecH5MJZNaOOzoiMiQx2OPoQeEI8lv0IG3b0bdYfMLkq7LvLuzhmIPQpKhsIAJO
VbJBtR3g1Wx35/PkKdKstFAZICbvcxrAR2kzaZSjTN7n0tVqKPzW0YIq0Tqx6N8d3uayUPOv7XST
l2pcW1tZh1m++9uqFciZjCj1JS0xBHSXDtP+DrzxTVp+kEqu6dzOZY+imfgo6J+KGZw/L5Q1ObKC
1/Ppqpf9II3e8eTb/aIRTQSIcKHvUziEaB/PCzzttFD3oeJSKNkgKVRhVzAC6aTZ8IgS8FRUPz2n
oA9ICeS5/n1BApOhE6UiU3GMSCMeoWhBGjWKMTSXxYSTRqC+Y0mcEoAbZ0otSO+E6fQv9GTYmRhP
v76DVIarw8gYWxjg3YZ5eyDcgZsapPJnE+BwWMoAixEh9uMtcXZGUgu4/p/TBEJNFCVN3h1d0uUB
6Hb7yyLiuppUT/U9EhbzfNZBkODtfR6hnWG5qQ20O2X9Oiwz9s70jFuj3LnH9kC1WUJ9qB5lrlWq
BByEcRp/8anQ2jjXGu/gupOIivxQFnnc2a4+SUNBv6qlS4nwmTqRIeyFU5DZ17lYOx6Lj1OkFd3v
myL1NhZmdsjhm8K9A+JCW0PVYuQQ6gGw3M+Qd4uFB7334UTEFvsH9eNMA3L14FEBLoqYq+TSQV+W
sd3ArcHBcJSwpZcXCsfeNRvYIKpGfyyAW1gxWhSdCv1qYGTXN1d+FNHtpnvz28up44riYfzZg7Qn
XG9BagFpcWdpqHVFEEfRK25ROTHnptjuJ6zPgHPOVVYGJE2GOszPvhDa+bRaStaMVdCR+CRsHX3N
tqaSUxpCJ2VZfoNB2HvVOu9eEJVR5Beh0M5dzsbalKdutxLhzDNgclP2UJHYdUFGBRav1t7utAKa
JxretKlfuBwPXPnGfeFQKX/XRT2nQvJozIr8ehmdAyqDM4HY/6auKl63dqTbeAPjoIlvdJQRzdkU
ZsXYROK6RDv5hOvE2QiPOyLC9XKAys472Dg2u1wmd9CWdTpaWuhtVohvgAwW7SlT1eoUz7vwqsib
jcdns+bSDLVkP6Yba0Yx81YXN1mLHPtLOxKv+eLVvmKBu6dypCNDVOHNXB0Sprxzps6jCYWw2OaN
BgPIqaWmSZsrST1wAVlMrgWmZjvyTC6MT+dDTO8imeDRftHNrEUl85aUISoLXz3vL/IzDGITfbUR
JWDk5YWvelZUdWSATwgyY/mjrZh2IP7gYGSb6t7zbvESNPAYq2FbzTvkgYVK2UK6cH0TLBaEuqfR
vvCUsrn2CVoeP82qTntOEaES0F1kSv+JiA4IBkpWl3cuzYmxuMAoQCPUzLLjQXmjE0mCjQiSjwO8
OgMrcZ4kjrNKtJuxQjVVYEyZ6JZX8iVix1uwTnIX8mjIWecYSGQYDTLak114E8yLrsOPBqYpMomC
GaAKz5QGXVh+JsQ7vVskiosryGh/fpe88JMsKrGtUY4TkoTs0cj+ngKuzxZrVLt6M449h6u+nDmH
UYSDQjtuO01NFXJglnpN79zTUMtNDRH54qkv+GNU4sCfh1B4BFd5RLg0Dqgs+iHw2WLFAPWlg6Ci
C7E2ehnw611qmE7P4OrSSyAqBQmyUkWVwB/tmIq+2N6Z2vlq7QjDUijDe/pm0CurfNg435GmV2K2
ns5amgnT4bxjfzozsGfGISMq3CUs1XzmfpzOO1Uv2pIea7I1GK7JV81oqpjVhM5OKuY5NGvMGpMR
Bxovl7Zta7nX7WFKDCNXmZrufiGU9AGX9H7KO56U5JW2HtreSIgEeN+Y3YoGV5/jC8ipZ/2sbNwt
VhTrduXwNqgYywG3IAP5Vg0i4db6rICtsI3bOUoljItfWkyujjrNyo6e5UEbMXj8nR26iCj9hwqV
0KeH0QqmsrYm5LAz8LPN9EaS+JEWtFt7ZQ2czi1oof1CfnZWGJI0vjojMtTeq02uBpSnzR1R0YyK
Sxde1RStQ18Imwx0aKPfjbkqk9Os8nsvAaUsitKH8gbAPrKoK3e63Em3FWAkR71Wip6LACoWeQlW
0210XgA262dVCGAE16+Xu/rAugiQhbQK+yhpPAZEDFxPUcLxSiwUzfm4kEU5P8X5LUqs4eiNOx+O
BjLus7M9YgzZQklbpSGcwP6jY514YKgnNl0+y/128VjzW9epj8pyDxHOTe37HwNp29U1NCMTNSjw
e+dEIPwXCDqY57ZaNNEpS1QdmoY0klF1z1WzbhMF5FhRb+RwkoEbVcWlGY0a2qLxBDmqFye+8hVL
ZXoGRq9E7XkjU26IqFwR9XPG6ymPJc1hPYlPxbxQ01tJa+90+z93QpCEX4SJRLxeHXBdmnTWzh48
dT+UjZoyVa4CSw1IVmtKflp+/oOp314EvV+D1v8iJ365qAr4MAZlxXgOZ0wxtUXJmidwt5PgDFCS
8A81s6WKp0BPSlOP2BRmdb3sWwEDGquSE38WUh/DiM1DuX4CSGOKmoeWMb5APUBC26/A30EnG/xe
CfBnQgO+avPlLc6ZNyZ/zi+4gLukcOpAhjYoPbTwdILIXRgrFKmN5KA6jWHusc9QeDKprPXP0MYO
5SNtOnJRArikv0ED65/brqM4XuCh+bgdVm6p6ILt5w+UI3Dohyn88cD6n2Ti0lAwf8JxC3ihJSTk
KmikFXNJNDod2qg6rs/CabYLCsICsWrPR3PbyTXyA7ZqYDsqs8qC+nRG8Qz1NxOnSraHd8hzooj7
BfZOIA51w1dEnNdHQ+TFDi7TiVoCAW9IuPS2UnZhSfbu/fGJCp+sxAiVPXi/9Dk38sG/eekbiHOm
rEbkjjg4H6hhcqW+UeKXFfYx67D5ZGotaN7KsmIQ969JkspR+lMCNml7WxpfrZz0z+KtW9OGmd9u
rv7p9URg5ya/gPzGRgPswqDXnUlJupAH55NMBAmDOUc79a/nxQKxE4Pvt3YxbcuK57IKhstSBKAf
2VzGvRJBXQeN1OfCPhrXEyMH3gfhuIscpPWpHe5JPXH6XqfMhYCU5hrjQycu81OG/wC6obEkcQyC
0QA2Gjz4y9BKLql6W0HNuCmIG4QGYNsSab4U5pThwAR8OjwS/Jk7UCzMI3pTHx96g2UR0AJXfhb+
Jzi5vlg8Yt0b71hrqlFMz6kxzDkPOfqu8wsGKoA+zLU42oXPGuirdq1skxnf0uVjC88ZsWvYhNAz
xZP1zxMVZ/bD9567A0Hz2SrI4pudbUKzPfO3A+uo7anXEiK0ZgH5CSbQpRnYeSqLl2QNWFftwZgR
4lXskQ+udGHoRrHqKOe+kS/z1P5gJgm4iVpZgBK6pGgK5TviOp4SD+1zXWYi20VXt4w/xHmhNztM
3hO/ZbwUqOJh/P85oBqHEUpffSCx7mm+bkg3lMkLZ+pXrRw65jkIrM+um3EncrSosczJp9CBhvQa
vrkIRbKQDtkVwx30fcnvpGowf8vxpTecOFHo+KbItf88abJ/EVAMJ5sVxIYN2q5B/yjU/31truwZ
cp+usJMm09Si8JGselOFw8bK374zfITHJB41czFqP5/SKntT3rdXNL7NET/7aruoZ6T0L1R15FYT
33YsBIB8ehanxWuoxNEe6OUCCeG5KwHpZ+01hPAXlHNEu2dArThK3UvqAJAMDb6TPUr7276XzabW
LqeGC5/EexPRheapgu2LmtSS6R/HiAoDjzogvVy+raFgFTHBVnEP67Oje8fnv/bzigvh6BBKSAFg
rR6A7jc5CyBpXx6nN4lQDcTgKfA4CI95M9vejcfVfON06UFXjvoRSUPSPH8cfocEar9feJMPGfcF
JH9HMuFY8d+37Ac4vRaeSS1Ei/K8v4mIhsRQiSCLFuErXBSmitxquE4LARy8nA2ICNXcX+zS4txx
j4W6aahx7JJ9YyoXGL+9fXCQdN9gu+HI+n7t6qWbv7w4H8838OoTmBP2t2RXwQEhIjHVYPfzTK0r
ad1S6o3OzTZkjrkFDXdGjboFQPSyxLIPMnc5F65SMwYKkahYi13zvr1QWi1Av38DvkSinCXPTvfr
wmvGqs5YEKikU3mhmQ3kLxydEIFz/l9+nRVcbFzeCVGJm2xAMX2Oyz0oeG/SZOukL1YkSP5GIGj8
s6z6v3GnXIL5/+mnlBaR8QueJA6JbX2ZjGXQzVkGUbHfnV0Wb83UrvBBmPGCcY5v5OONynquXvmq
46U/f1zrStGZ/cjFOr+yc7MGEYu4PrazRu/u7ENwpblX125OCW9q5bOvl3cBIS5RuOxvOFvY3ADH
3VZlZz0yA/JrRkhJ+vDBZnf7S6vmyg+sdGpsUCDAf+oQm+/SKNncLy6exTf6QK8pY7vZ9My6NL+D
ZtwtXLhJqpjIb/tFAVtTEa2+G5OL2JGG9f93jWeXwBn+dy3mMjkppxTAXu/Z56O0M/q1crr9b8/x
WsEMAA92biydqAE/vuepYXuXGm2BjXRBvN1ZNPbOslmTHKhVCJGJOj48JSH/gD2YKEWu6G4mbwlX
RjUG/hlWMKtoOhQwYLc9gXQ6u+/GF1XNpOf71StqSwHUEpOsHa8xDNiy/dhHrMmGUJqqaSEUl824
6uXDwQ1bwZbQ9gD9bGmfN4EiWZ5GlJilGVTmtD6JBCKOZRHZ4vgkmx6PAEtZOIQY9dcQ+qhkvrkN
vBFk3WwD3YRLmgwoJ7uwnrTgG7jW+Sb0IXEYH3jYJ8O9Np7IacVadU7weeZ2a+/X3vozvlc4G9iD
k/4CW4SW6xgykH5qTafqQIHclfAU1eem7FBC+QnXZGtiJXXOpOXz9hbJDBKyoVFmP/JFbUhTPu03
CVGR2/s39gaAgHCopHQElfTDfF122O3+qspbgJFhN2rJH3pIlB7zNZz0sfpV931FEuIeNdQNdohZ
U+/CEpxvDsWhZ8M9TzGq/vW5hMq4rxSmubp/BeMEhVWH4XaekYvWl/UAb+oI+WlFFsA06eFStqjL
5stSOT9ZSOy5NlK6srzaFyn1wPDTtckLrXJvTewOkXPmB+RjnLkbkIa2DerjhHdkmY4iWqI8PsLJ
VESIUjK66MvB+aVSiy9WhlpU5PUx/Zo4iBP7L60gRKjTXf+ixpFXRh1FTOlK54TtdVfJTBdlUwfo
UgMLgKjbBrfT04R6nm3nlQEOTLLr0WU0Azfs5sB14Hp3Gazyae15l6kkGvE5aTgYYIQr0VzKfExG
RJHtZ6UuwW1R9pa+gxDzgq4H0OYikiyHvpsKNQS6vwe18U+nhfGttk+VbctgX9hTL6MiIJs93bu1
7DGVa326Lkus1qB8f/pgihS2uM0grP9ki1CGvOvC168uwfPHXksZTtUGIt8qKbEUCerTHgHXcHXj
erxE66zLsbF59aWguQ9BdU4X4YWjsGDudw785X6dPrEFuCnXTI2pBOi5bjlN3UlWQ32opb1pHTh5
dh+oXkqP+R72Wr7JCao8ojocSncgA0vZOzHwrZ5a30xdTdq5F2iVCCE2VdLulbyzMDgrf64iEw+F
t7OxHNHh+uJv8nD0hDzf61SyARkhoYxy7dtxa7eeS3A0Rp84PAwqTICV1eq1kRZOYduXfbmnnv4L
jtkuvjcnR1FTOI3nUn+daK5y9Wyemj7ResVKj1+zSMtxOaJ6jQXAN/0n8vDTy7HTer4MppL6GFcw
pmyiwNIWqFS35yeyr7+IJDWIhSQJnyqkvtrBwWZZRAIL+ox+qCyhP3vdbY0VWpNZe5CjsnDtwGT1
HvsyUjZ89EUxhzIKLDQxNsv0UpMU9HiXGpEYwHiifNfLfLbLSpxmR3YF5H/77MUOtVRUQ5u6kTM1
hRF9jrYTVgyx0w9piVIGJeFpqz5rAirhAPd5z/g3DbOpmbuxt8wbeJ0K4O23FILh18hndVGWYMUp
MMH5VbywzPSNpqa1KsGrHDxSbMvOw+injgAyZPF3w5FmW0o+F/tPm5u9y4urwGEowyeC15z9cj+d
A2a9SNBWyZHAjeomk0ajfp2GNbci8hEeDiACaPGcgHVDEgUaABCCskmLrQA6itjXhTeQlzzy7vM7
csnybSWoaoEMUexL/s3j+lgbq24Hh3JYoYepluhayI3Gp3AQ4rmoEmUugcn3Ov9N0KO1+NQiMIbX
JdkVjcIUXIpUPA8vvVW1KC9kr3pM3XWOG9Hlv3xoIPaTxkvKxSpcDucIPXxHYuJOr/iWg8GqiR9b
uPxLySbaSUESLfJaKSIPPVzucSOtDD6Qc54i4VdtkRourPiJqx4wqrqKFNWjOAGdHK+eVpz2t0No
WCp3LC05UW2Jr/3Z/t/e29KlqmI4eL9aZFjWfxRT45xWIUAB7GMVFnfdh2opHDptKLXOaTLqSxXy
esvw8NsDVArWN7BJDKFhLihTSNvnSxW09cKXivlb+UFCuI1fIK8j7EcowSxWmQp8cVfY65Ufgv2G
6QEh0RNiE9SPXnwT0kGh18fMwqST0ZupzBMTf90rLbxJiZ4yDTfG7IZrSlavg5AplFhlj31nwsyg
uGZ9HdKcWadz3hx+Zua63cjcSxwLG2+86CP8QlsMYErZlm3J3aDVfSryioFFyQi8fiC41iyhHmPl
ZG6Djyym3oRwWqSUaxwVIesWKbX3be6jiAHNX+oS4BTjy00ze32TWONl2LKN6PfxPdkCvNB3fk/Y
8qBtXrYi8L1Vv2kBYAtZj08SFkqcs24JUHqfPSb809gw06exh5MwiHodWj1JpSEaapKxIkoAYVc3
A4OaLNGGdlIwR9kqlpBIgy4OPZzBatS3lbDXDP3E1U9IJIVCC4xXZLOsTZ/EgvFvZTw+VUuGH7T6
o4PurLBIV27Rp0Nvo++xlhM7dDnk3sV4GSZYg+CM4eAq0iEhUypInCxBHvuvJQcOUbQPVm1Mouew
0NRPg0PiAr7KRHETyt2iCLisolMQk3bQUBglDFAPVDL8qG7JUfNkTe9vARk+6NyY5KIFsYnTcNJh
A5wFY6MZgGfyBJ8Lx4SXjMmI5LOdyWfJXQ6mgtExsZ2O6/GEJNHsiHoDqT3hDpQ2QT3hA3KKSnZv
I3+gf1969pZUGrQpEzF2w9cmKpFT2Oz3c5qz+Z0NzRpUvUeDK1v1I9wItDzV4GppwlxykMSYyZNY
pYRCYUTxAT7eWuaLXIFOsiW7qaScrghShPGbDczYqL5296aYty7fo5jk3L+bmjtXe9FadiJ/Lf19
MLsOPw9Ml1JAawpSbNeE7rgx8JEwZkHVXd85+c2qZHfI2cy832Q0RgxS3qIzDYmKlcqfB5N5nz9A
PAkuEYZ9IUoNTkokiumdjN6w/UTw7hISMQXo2z8KWQhx2ywWre4EbTXgo4qLJIB+ftSYds3u2xB1
+99bOezmIoBAXhKDh0smb8btpxjflr0x42dxY+U1LinjZ6j4/NPYKUZ1QZTKVYTsqDcgDm/4s31x
R4suKX/G8SNadLHK6obzHOuysQA0QkVhm+3s7vEPTrcOxuMyAG/YUYeu/2t0NoAXqTApGL3MBVBP
qzYUuQqrP2AHqLkDX5NvP4DKRno74mirgH+v/BlyrD3ujlREMVB5Ej1TzSKarGkpQr93+XxQwHbV
nKf83j7DMU9pp70SXVlpxSVNe1o3NWTIVN/PqVojtNiJcFw0HSA6OVhTmPy4sBEf3xCrDkkMFgGk
suh2yToUKqpG9vLvuFO73D+Gl7zCSCUUeZmUN/Uf/TX6yiJsDM1zwsnpUty7QStMMgmx8aBEDbQn
37Z6MZOMqe8IDkvxQPBHEZualQ1S5cJJctFaYx+yJw5ksXtssdLW0LJ0zr0uW9zSgXNkDrJBZCwJ
7lVddcKAejdzwTLWOt8yoD+HqVFbvRhsLZ9IhxVXkRXqd8LO4DGI/V1SYXnMnkkyb3voDWsDHQzc
bFySWpelWO3fpObgXpVdX2qnYX5f6YE4OZ/EJqoHEQNBIai1SO5BtKVytyscQKSCXzp7Vp0ZGKke
+9j8HWSL4mEcXZd1RYmV2KdHcz1FbGQouGVepGFpI+Lr9UPuSl8H/P1Op87s0jW3p4C5EIx2SFnF
iYswbtK9jFXmb/a19aUR4dpUVgkTn+r+8mzu4rPRpfZ2avyjeMVK5PV4wvN+ajBsGtvfHkdAnn6h
hbf8iIU985R88kKqArGNds9d6OwXiDyGeOT/lrB2rDvQKlZLIpSLPP6SWAzD/dAfqaPY7y7aj+ZF
26L9anAR1YY6yt5zuMQoLSvzl/ZlCarcYpDq+cyVxFpWU9IDLBDbkxtiMR3eZL1jKr3/NvKT0UqQ
8f1i/2ySrVIr5Q==
`protect end_protected
