//------------------------------------------------------------
// Project: HYBRID_CONTROL
// Author: Nicola Zaupa
// Date: (2023/11/08) (16:19:35)
// File: tb_hybrid_control_theta_phi.v
//------------------------------------------------------------
// Description:
// test-bench for the simulation of the hybrid control block.
// The idea is to test the proper operations of the state 
// machine.
//------------------------------------------------------------


`timescale 1 ns / 1 ps

module tb_hybrid_control_theta_phi();

reg clk_100M;
reg signed [13:0] vC, iC;
wire signed [13:0]vC_ADC, iC_ADC;
// reg [1:0] sigma; // from table
wire [1:0] sigma; // from modules
wire signed [31:0] vC_sim, iC_sim;


simulator_LLC #() simulator_LLC_inst (
   .vC_p(vC_sim), 
   .iS_p(iC_sim), 
   .Vo_p(),    
   .CLK(clk_100M),    
   .RESET(1'b1),   
   .sigma(sigma)
);

simulator_ADC_14bit #( .mu_I(65), .mu_V(140)
) simulator_ADC_14bit_inst ( 
   .v_in(vC_sim), 
   .i_in(iC_sim),
   .v_ADC(vC_ADC), 
   .i_ADC(iC_ADC)  
);

// CONTROLLER
hybrid_control_theta_phi #(.mu_z1(32'd86), .mu_z2(32'd90), .mu_Vg(32'd312000)
) hybrid_control_theta_phi_inst (
   .i_clock( clk_100M ), 
   .i_RESET( 1),    
   .i_vC( vC_ADC ),      
   .i_iC( iC_ADC ),       
   .i_theta( 32'd150 ),   
   .i_phi( 32'd15 ),
   .o_sigma(sigma)
);

// call the block to be simulated
hybrid_control_phi #(.mu_z1(32'd86), .mu_z2(32'd90), .mu_Vg(32'd312000)
) hybrid_control_phi_inst (
   .i_clock( clk_100M ), 
   .i_RESET(1'b1),    
   .i_vC( vC_ADC ),      
   .i_iC( iC_ADC ),       
   .i_phi( 32'd5 ),
   .o_sigma()
);

// create the clock signal
always begin //100MHz
   clk_100M = 1'b1;
   #5
   clk_100M = 1'b0;
   #5;
end


// initial begin // generate the input voltage and current
// // // samplings of current and voltage

// #10;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001001; // iC=  -55 
// vC = 14'b0000000000000000; // vC=    0 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010100; // iC= -108 
// vC = 14'b0000000001001001; // vC=   73 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111010; // iC=   -6 
// vC = 14'b1111111111010001; // vC=  -47 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011011; // iC=  155 
// vC = 14'b1111111111110100; // vC=  -12 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001001; // iC=   73 
// vC = 14'b1111111110001011; // vC= -117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000001; // iC=  -63 
// vC = 14'b0000000001101011; // vC=  107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100011; // iC=  163 
// vC = 14'b1111111111111101; // vC=   -3 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110011; // iC=  179 
// vC = 14'b0000000010010000; // vC=  144 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000000; // iC=  128 
// vC = 14'b1111111111101011; // vC=  -21 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111110110; // iC=  -10 
// vC = 14'b0000000000100010; // vC=   34 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100011; // iC=  163 
// vC = 14'b1111111110001110; // vC= -114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100001; // iC=  -31 
// vC = 14'b1111111111011001; // vC=  -39 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010001; // iC=   17 
// vC = 14'b0000000001000111; // vC=   71 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111001; // iC=  121 
// vC = 14'b0000000010000010; // vC=  130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100111; // iC=   39 
// vC = 14'b0000000001001011; // vC=   75 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011000; // iC=  152 
// vC = 14'b0000000000001101; // vC=   13 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111111; // iC=  191 
// vC = 14'b0000000010001000; // vC=  136 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000100; // iC=  132 
// vC = 14'b1111111110111111; // vC=  -65 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111100; // iC=  -68 
// vC = 14'b0000000010000011; // vC=  131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011111; // iC=  159 
// vC = 14'b0000000001101000; // vC=  104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101010; // iC=   42 
// vC = 14'b1111111111001100; // vC=  -52 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100101; // iC=  165 
// vC = 14'b0000000000111001; // vC=   57 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111110; // iC=   -2 
// vC = 14'b0000000001001000; // vC=   72 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101011; // iC=   43 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010100; // iC=  148 
// vC = 14'b0000000000110100; // vC=   52 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000010; // iC=  194 
// vC = 14'b0000000001011001; // vC=   89 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111101; // iC=   -3 
// vC = 14'b0000000001111011; // vC=  123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100111; // iC=  231 
// vC = 14'b0000000001010101; // vC=   85 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101111; // iC=  175 
// vC = 14'b0000000001100010; // vC=   98 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110010; // iC=  114 
// vC = 14'b1111111101101111; // vC= -145 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010010; // iC=   82 
// vC = 14'b0000000001111000; // vC=  120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111010; // iC=  122 
// vC = 14'b1111111110001000; // vC= -120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000110010; // iC=   50 
// vC = 14'b0000000010011011; // vC=  155 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000100; // iC=  132 
// vC = 14'b0000000000111011; // vC=   59 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001000; // iC=  200 
// vC = 14'b0000000001110000; // vC=  112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100010; // iC=  354 
// vC = 14'b0000000001011000; // vC=   88 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000001; // iC=  193 
// vC = 14'b1111111111011100; // vC=  -36 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010010; // iC=   82 
// vC = 14'b1111111110001100; // vC= -116 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011011010; // iC=  218 
// vC = 14'b0000000000011111; // vC=   31 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110000; // iC=  304 
// vC = 14'b0000000000111001; // vC=   57 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000110; // iC=  134 
// vC = 14'b0000000010100110; // vC=  166 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101011; // iC=  363 
// vC = 14'b0000000010000010; // vC=  130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111000; // iC=  440 
// vC = 14'b1111111111101011; // vC=  -21 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110110; // iC=  438 
// vC = 14'b1111111111010110; // vC=  -42 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000010; // iC=  450 
// vC = 14'b0000000000000011; // vC=    3 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100011; // iC=  355 
// vC = 14'b1111111111011110; // vC=  -34 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001110; // iC=  334 
// vC = 14'b0000000000100110; // vC=   38 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001110; // iC=  206 
// vC = 14'b1111111110010010; // vC= -110 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100000; // iC=  480 
// vC = 14'b0000000000101001; // vC=   41 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001001; // iC=  457 
// vC = 14'b1111111110011111; // vC=  -97 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010010; // iC=  402 
// vC = 14'b0000000001010011; // vC=   83 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110000; // iC=  432 
// vC = 14'b0000000010101101; // vC=  173 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010001; // iC=  529 
// vC = 14'b1111111111100010; // vC=  -30 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110110; // iC=  438 
// vC = 14'b1111111111111110; // vC=   -2 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101001; // iC=  233 
// vC = 14'b0000000001110110; // vC=  118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011001; // iC=  537 
// vC = 14'b1111111110011011; // vC= -101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001011; // iC=  331 
// vC = 14'b0000000010010100; // vC=  148 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111001; // iC=  505 
// vC = 14'b0000000001000010; // vC=   66 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100010; // iC=  290 
// vC = 14'b0000000000110000; // vC=   48 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001110; // iC=  590 
// vC = 14'b1111111111101001; // vC=  -23 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000111; // iC=  327 
// vC = 14'b0000000001011100; // vC=   92 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001111; // iC=  399 
// vC = 14'b0000000010001001; // vC=  137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111001; // iC=  505 
// vC = 14'b0000000001001100; // vC=   76 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110100; // iC=  308 
// vC = 14'b1111111110100011; // vC=  -93 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100101; // iC=  421 
// vC = 14'b1111111111000101; // vC=  -59 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101110; // iC=  622 
// vC = 14'b0000000010000011; // vC=  131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111110; // iC=  638 
// vC = 14'b0000000000100101; // vC=   37 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101100; // iC=  364 
// vC = 14'b1111111111011000; // vC=  -40 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010011; // iC=  339 
// vC = 14'b0000000000001010; // vC=   10 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101110; // iC=  494 
// vC = 14'b1111111111111100; // vC=   -4 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010110; // iC=  598 
// vC = 14'b0000000000011110; // vC=   30 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011100; // iC=  668 
// vC = 14'b0000000011001100; // vC=  204 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110010; // iC=  434 
// vC = 14'b0000000010011101; // vC=  157 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111110; // iC=  446 
// vC = 14'b0000000001101000; // vC=  104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000111; // iC=  519 
// vC = 14'b0000000011011111; // vC=  223 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101001; // iC=  553 
// vC = 14'b1111111110110101; // vC=  -75 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010010; // iC=  530 
// vC = 14'b1111111111100101; // vC=  -27 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111000; // iC=  696 
// vC = 14'b0000000001110010; // vC=  114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010010; // iC=  658 
// vC = 14'b0000000010001001; // vC=  137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100101; // iC=  549 
// vC = 14'b0000000000101011; // vC=   43 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110010; // iC=  626 
// vC = 14'b0000000001101000; // vC=  104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100000; // iC=  608 
// vC = 14'b0000000001011000; // vC=   88 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110110; // iC=  630 
// vC = 14'b1111111111001010; // vC=  -54 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111110; // iC=  638 
// vC = 14'b0000000000110010; // vC=   50 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011111; // iC=  543 
// vC = 14'b0000000011010100; // vC=  212 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000000; // iC=  576 
// vC = 14'b1111111111001011; // vC=  -53 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001111; // iC=  655 
// vC = 14'b1111111111001110; // vC=  -50 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000100; // iC=  580 
// vC = 14'b0000000000001011; // vC=   11 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110011; // iC=  691 
// vC = 14'b0000000001101011; // vC=  107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111010; // iC=  570 
// vC = 14'b0000000011000000; // vC=  192 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110110; // iC=  502 
// vC = 14'b0000000100011001; // vC=  281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110011; // iC=  627 
// vC = 14'b0000000100001000; // vC=  264 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010111; // iC=  791 
// vC = 14'b0000000011011010; // vC=  218 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011111; // iC=  543 
// vC = 14'b0000000001110011; // vC=  115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101010; // iC=  746 
// vC = 14'b0000000100000010; // vC=  258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010101; // iC=  725 
// vC = 14'b0000000001111110; // vC=  126 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001111; // iC=  783 
// vC = 14'b0000000001101101; // vC=  109 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110001; // iC=  625 
// vC = 14'b0000000010110000; // vC=  176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011011; // iC=  795 
// vC = 14'b0000000010010001; // vC=  145 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111011; // iC=  635 
// vC = 14'b0000000010110110; // vC=  182 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001101; // iC=  845 
// vC = 14'b0000000010000010; // vC=  130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100100; // iC=  740 
// vC = 14'b0000000001000011; // vC=   67 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001111; // iC=  719 
// vC = 14'b0000000010101011; // vC=  171 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101111; // iC=  815 
// vC = 14'b0000000001011011; // vC=   91 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111000; // iC=  632 
// vC = 14'b1111111111111101; // vC=   -3 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001000; // iC=  840 
// vC = 14'b0000000011000101; // vC=  197 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111100; // iC=  892 
// vC = 14'b0000000011100111; // vC=  231 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111100; // iC=  636 
// vC = 14'b0000000010100011; // vC=  163 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011111; // iC=  607 
// vC = 14'b0000000001111000; // vC=  120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110000; // iC=  752 
// vC = 14'b0000000011001011; // vC=  203 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110000; // iC=  688 
// vC = 14'b0000000010110010; // vC=  178 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100000; // iC=  736 
// vC = 14'b0000000001010010; // vC=   82 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100111; // iC=  743 
// vC = 14'b0000000011011110; // vC=  222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010011; // iC=  787 
// vC = 14'b0000000100011100; // vC=  284 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b0000000001110110; // vC=  118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011101; // iC=  797 
// vC = 14'b0000000100100011; // vC=  291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100011; // iC=  611 
// vC = 14'b0000000001010100; // vC=   84 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111110; // iC=  766 
// vC = 14'b0000000011110000; // vC=  240 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010111; // iC=  791 
// vC = 14'b0000000010000111; // vC=  135 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110111; // iC=  631 
// vC = 14'b0000000001100101; // vC=  101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101100; // iC=  684 
// vC = 14'b0000000100000101; // vC=  261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101011; // iC=  939 
// vC = 14'b0000000001110000; // vC=  112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111111; // iC=  895 
// vC = 14'b0000000101011000; // vC=  344 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101010; // iC=  682 
// vC = 14'b0000000011100000; // vC=  224 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111100; // iC=  700 
// vC = 14'b0000000100001011; // vC=  267 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010110; // iC=  726 
// vC = 14'b0000000001010001; // vC=   81 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101011; // iC=  747 
// vC = 14'b0000000100010110; // vC=  278 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111001; // iC=  761 
// vC = 14'b0000000101101000; // vC=  360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100011; // iC=  931 
// vC = 14'b0000000011010111; // vC=  215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100100; // iC=  932 
// vC = 14'b0000000001111011; // vC=  123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011110; // iC=  926 
// vC = 14'b0000000011011000; // vC=  216 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101100; // iC=  940 
// vC = 14'b0000000110011011; // vC=  411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110111; // iC=  759 
// vC = 14'b0000000100101100; // vC=  300 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010111; // iC=  663 
// vC = 14'b0000000101000000; // vC=  320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001000; // iC=  840 
// vC = 14'b0000000011111010; // vC=  250 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111000; // iC=  952 
// vC = 14'b0000000011100001; // vC=  225 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101110; // iC=  686 
// vC = 14'b0000000101001110; // vC=  334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011100; // iC=  860 
// vC = 14'b0000000100010000; // vC=  272 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011010; // iC=  666 
// vC = 14'b0000000110001001; // vC=  393 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110100; // iC=  948 
// vC = 14'b0000000101010001; // vC=  337 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011111; // iC=  799 
// vC = 14'b0000000101110110; // vC=  374 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110000; // iC=  752 
// vC = 14'b0000000100000001; // vC=  257 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011111; // iC=  671 
// vC = 14'b0000000100111010; // vC=  314 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011011; // iC=  731 
// vC = 14'b0000000011011011; // vC=  219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111101; // iC=  701 
// vC = 14'b0000000100001101; // vC=  269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101011; // iC=  875 
// vC = 14'b0000000101111101; // vC=  381 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110010; // iC=  946 
// vC = 14'b0000000110111010; // vC=  442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011010; // iC=  730 
// vC = 14'b0000000010111110; // vC=  190 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001111; // iC=  911 
// vC = 14'b0000000011001101; // vC=  205 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100100; // iC=  996 
// vC = 14'b0000000011111111; // vC=  255 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011101; // iC=  797 
// vC = 14'b0000000101111001; // vC=  377 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110000; // iC=  816 
// vC = 14'b0000000101010000; // vC=  336 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110011; // iC=  819 
// vC = 14'b0000000101010010; // vC=  338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110110; // iC=  822 
// vC = 14'b0000000101001001; // vC=  329 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010101; // iC=  725 
// vC = 14'b0000000010111000; // vC=  184 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010000; // iC=  912 
// vC = 14'b0000000110011111; // vC=  415 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010011; // iC=  723 
// vC = 14'b0000000100110110; // vC=  310 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000000; // iC=  768 
// vC = 14'b0000000111110110; // vC=  502 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000110; // iC=  902 
// vC = 14'b0000000101100000; // vC=  352 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011000; // iC=  856 
// vC = 14'b0000000101000110; // vC=  326 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111111; // iC=  959 
// vC = 14'b0000000111110001; // vC=  497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100010; // iC=  738 
// vC = 14'b0000000011111110; // vC=  254 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000100; // iC=  772 
// vC = 14'b0000000101001010; // vC=  330 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111111; // iC=  767 
// vC = 14'b0000000011100111; // vC=  231 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000001; // iC=  833 
// vC = 14'b0000000100100101; // vC=  293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110101; // iC=  821 
// vC = 14'b0000000110111100; // vC=  444 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000100; // iC=  708 
// vC = 14'b0000000110110101; // vC=  437 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000101; // iC=  773 
// vC = 14'b0000000110101111; // vC=  431 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011110; // iC=  926 
// vC = 14'b0000000100101101; // vC=  301 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000010; // iC=  770 
// vC = 14'b0000000101001110; // vC=  334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010111; // iC=  727 
// vC = 14'b0000000011101111; // vC=  239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000100; // iC=  964 
// vC = 14'b0000000111101010; // vC=  490 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101000; // iC=  936 
// vC = 14'b0000001000011010; // vC=  538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111100; // iC=  764 
// vC = 14'b0000000111100000; // vC=  480 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111101; // iC=  765 
// vC = 14'b0000000110100010; // vC=  418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100110; // iC=  870 
// vC = 14'b0000001000110001; // vC=  561 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101110; // iC=  814 
// vC = 14'b0000000100100010; // vC=  290 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001111; // iC=  719 
// vC = 14'b0000000100111111; // vC=  319 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110111; // iC=  695 
// vC = 14'b0000000100101110; // vC=  302 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111001; // iC=  825 
// vC = 14'b0000000110010000; // vC=  400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000001; // iC=  705 
// vC = 14'b0000000110011001; // vC=  409 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010100; // iC=  660 
// vC = 14'b0000000111011011; // vC=  475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100011; // iC=  739 
// vC = 14'b0000000110010111; // vC=  407 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010100; // iC=  724 
// vC = 14'b0000000100010010; // vC=  274 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110001; // iC=  689 
// vC = 14'b0000000110110101; // vC=  437 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110000; // iC=  880 
// vC = 14'b0000000111100110; // vC=  486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110110; // iC=  694 
// vC = 14'b0000000101111011; // vC=  379 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010010; // iC=  786 
// vC = 14'b0000000100011111; // vC=  287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101011; // iC=  683 
// vC = 14'b0000000100100001; // vC=  289 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110011; // iC=  883 
// vC = 14'b0000001001000111; // vC=  583 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101000; // iC=  936 
// vC = 14'b0000000110100010; // vC=  418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101101; // iC=  685 
// vC = 14'b0000000111110010; // vC=  498 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000100; // iC=  772 
// vC = 14'b0000000110110000; // vC=  432 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001100; // iC=  716 
// vC = 14'b0000001000111010; // vC=  570 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001111; // iC=  719 
// vC = 14'b0000001001001101; // vC=  589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011001; // iC=  729 
// vC = 14'b0000000101100110; // vC=  358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101101; // iC=  877 
// vC = 14'b0000000101001100; // vC=  332 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111000; // iC=  760 
// vC = 14'b0000000110011010; // vC=  410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111111; // iC=  767 
// vC = 14'b0000000101110110; // vC=  374 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001111; // iC=  847 
// vC = 14'b0000000110010111; // vC=  407 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001001; // iC=  841 
// vC = 14'b0000001000011101; // vC=  541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001010; // iC=  650 
// vC = 14'b0000001010001000; // vC=  648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101010; // iC=  618 
// vC = 14'b0000000111100110; // vC=  486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001011; // iC=  651 
// vC = 14'b0000001000011001; // vC=  537 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001000; // iC=  840 
// vC = 14'b0000000101101111; // vC=  367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101011; // iC=  747 
// vC = 14'b0000001000011111; // vC=  543 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101101; // iC=  749 
// vC = 14'b0000001010000100; // vC=  644 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111111; // iC=  575 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001000; // iC=  584 
// vC = 14'b0000000110010110; // vC=  406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110001; // iC=  561 
// vC = 14'b0000000111101100; // vC=  492 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010010; // iC=  722 
// vC = 14'b0000001000100011; // vC=  547 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010111; // iC=  791 
// vC = 14'b0000000101101110; // vC=  366 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000111; // iC=  711 
// vC = 14'b0000000110010110; // vC=  406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101011; // iC=  619 
// vC = 14'b0000000111001000; // vC=  456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110100; // iC=  564 
// vC = 14'b0000001010010100; // vC=  660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011001; // iC=  601 
// vC = 14'b0000000111100110; // vC=  486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011111; // iC=  671 
// vC = 14'b0000001010110010; // vC=  690 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101101; // iC=  621 
// vC = 14'b0000000110101110; // vC=  430 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011110; // iC=  606 
// vC = 14'b0000001010001010; // vC=  650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110110; // iC=  758 
// vC = 14'b0000001001110101; // vC=  629 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110000; // iC=  816 
// vC = 14'b0000001001011001; // vC=  601 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100100; // iC=  612 
// vC = 14'b0000001000110110; // vC=  566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110001; // iC=  561 
// vC = 14'b0000001001101000; // vC=  616 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100011; // iC=  739 
// vC = 14'b0000001001010011; // vC=  595 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000010; // iC=  514 
// vC = 14'b0000000110110011; // vC=  435 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110101; // iC=  693 
// vC = 14'b0000001001110000; // vC=  624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001100; // iC=  716 
// vC = 14'b0000000111110010; // vC=  498 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101010; // iC=  618 
// vC = 14'b0000001000101011; // vC=  555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001011; // iC=  715 
// vC = 14'b0000001001010111; // vC=  599 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000001; // iC=  769 
// vC = 14'b0000001000110110; // vC=  566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101100; // iC=  492 
// vC = 14'b0000001000110010; // vC=  562 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001001; // iC=  521 
// vC = 14'b0000000111001111; // vC=  463 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100101; // iC=  741 
// vC = 14'b0000000110111100; // vC=  444 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101111; // iC=  495 
// vC = 14'b0000001011010010; // vC=  722 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011011; // iC=  475 
// vC = 14'b0000001010011101; // vC=  669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001100; // iC=  524 
// vC = 14'b0000001000001111; // vC=  527 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001101; // iC=  653 
// vC = 14'b0000000111110101; // vC=  501 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011011; // iC=  475 
// vC = 14'b0000001010100101; // vC=  677 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111111; // iC=  511 
// vC = 14'b0000000111010011; // vC=  467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100110; // iC=  742 
// vC = 14'b0000000111001110; // vC=  462 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111011; // iC=  635 
// vC = 14'b0000001001010100; // vC=  596 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111011; // iC=  635 
// vC = 14'b0000001001010010; // vC=  594 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000111; // iC=  647 
// vC = 14'b0000001010000111; // vC=  647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000101; // iC=  645 
// vC = 14'b0000001011101100; // vC=  748 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111101; // iC=  573 
// vC = 14'b0000001001101001; // vC=  617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010111; // iC=  727 
// vC = 14'b0000001011111100; // vC=  764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010100; // iC=  468 
// vC = 14'b0000001010000111; // vC=  647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011001; // iC=  665 
// vC = 14'b0000001000011011; // vC=  539 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100100; // iC=  484 
// vC = 14'b0000001001110100; // vC=  628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110111; // iC=  503 
// vC = 14'b0000001000100000; // vC=  544 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011111; // iC=  479 
// vC = 14'b0000000111110011; // vC=  499 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100011; // iC=  419 
// vC = 14'b0000001000111010; // vC=  570 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011001; // iC=  409 
// vC = 14'b0000001011001110; // vC=  718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011000; // iC=  536 
// vC = 14'b0000001010000111; // vC=  647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000000; // iC=  448 
// vC = 14'b0000001010000001; // vC=  641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001101; // iC=  653 
// vC = 14'b0000001100000111; // vC=  775 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000100; // iC=  452 
// vC = 14'b0000001011010101; // vC=  725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110110; // iC=  694 
// vC = 14'b0000001011110100; // vC=  756 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011000; // iC=  600 
// vC = 14'b0000001011101111; // vC=  751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100010; // iC=  674 
// vC = 14'b0000001011001011; // vC=  715 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110001; // iC=  689 
// vC = 14'b0000001010100001; // vC=  673 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101011; // iC=  491 
// vC = 14'b0000000111101000; // vC=  488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001100; // iC=  524 
// vC = 14'b0000001000101010; // vC=  554 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111111; // iC=  383 
// vC = 14'b0000001001111010; // vC=  634 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001011; // iC=  459 
// vC = 14'b0000001011100110; // vC=  742 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011001; // iC=  473 
// vC = 14'b0000001001011001; // vC=  601 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111101; // iC=  509 
// vC = 14'b0000001000010100; // vC=  532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000010; // iC=  386 
// vC = 14'b0000001100010110; // vC=  790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011111; // iC=  607 
// vC = 14'b0000001100001100; // vC=  780 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101100; // iC=  492 
// vC = 14'b0000001010000011; // vC=  643 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010111; // iC=  663 
// vC = 14'b0000001001110111; // vC=  631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010010; // iC=  466 
// vC = 14'b0000001010101100; // vC=  684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101110; // iC=  366 
// vC = 14'b0000001011100100; // vC=  740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011000; // iC=  600 
// vC = 14'b0000001001110100; // vC=  628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011010; // iC=  346 
// vC = 14'b0000001001110100; // vC=  628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001100; // iC=  588 
// vC = 14'b0000001010100010; // vC=  674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110001; // iC=  497 
// vC = 14'b0000001001001100; // vC=  588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000100; // iC=  516 
// vC = 14'b0000001001111100; // vC=  636 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011111; // iC=  479 
// vC = 14'b0000001001111110; // vC=  638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011110; // iC=  414 
// vC = 14'b0000001001100100; // vC=  612 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001000; // iC=  584 
// vC = 14'b0000001010000011; // vC=  643 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001101; // iC=  589 
// vC = 14'b0000001000010110; // vC=  534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101110; // iC=  494 
// vC = 14'b0000001000110101; // vC=  565 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001011; // iC=  523 
// vC = 14'b0000001011110110; // vC=  758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011100; // iC=  476 
// vC = 14'b0000001000100010; // vC=  546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100011; // iC=  419 
// vC = 14'b0000001001000000; // vC=  576 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011111; // iC=  351 
// vC = 14'b0000001011010001; // vC=  721 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001000; // iC=  456 
// vC = 14'b0000001101001011; // vC=  843 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101110; // iC=  366 
// vC = 14'b0000001100110011; // vC=  819 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011010; // iC=  282 
// vC = 14'b0000001101011000; // vC=  856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000100; // iC=  452 
// vC = 14'b0000001100001111; // vC=  783 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011000; // iC=  472 
// vC = 14'b0000001101011111; // vC=  863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010011; // iC=  403 
// vC = 14'b0000001010011011; // vC=  667 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101000; // iC=  424 
// vC = 14'b0000001101011111; // vC=  863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111101; // iC=  445 
// vC = 14'b0000001011000100; // vC=  708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011100; // iC=  540 
// vC = 14'b0000001011110111; // vC=  759 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000100; // iC=  260 
// vC = 14'b0000001100111110; // vC=  830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000111; // iC=  455 
// vC = 14'b0000001101011101; // vC=  861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110000; // iC=  304 
// vC = 14'b0000001001011010; // vC=  602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011010; // iC=  474 
// vC = 14'b0000001011010101; // vC=  725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010010; // iC=  466 
// vC = 14'b0000001001101000; // vC=  616 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110001; // iC=  369 
// vC = 14'b0000001100111111; // vC=  831 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100000; // iC=  288 
// vC = 14'b0000001101001111; // vC=  847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100000; // iC=  416 
// vC = 14'b0000001101100101; // vC=  869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010011; // iC=  275 
// vC = 14'b0000001100110101; // vC=  821 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100010; // iC=  482 
// vC = 14'b0000001010111001; // vC=  697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100011; // iC=  291 
// vC = 14'b0000001100011101; // vC=  797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000011; // iC=  259 
// vC = 14'b0000001100101010; // vC=  810 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010001; // iC=  401 
// vC = 14'b0000001011101010; // vC=  746 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110011; // iC=  371 
// vC = 14'b0000001110000001; // vC=  897 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110011; // iC=  243 
// vC = 14'b0000001100100100; // vC=  804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110000; // iC=  496 
// vC = 14'b0000001011110010; // vC=  754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010010; // iC=  466 
// vC = 14'b0000001010100010; // vC=  674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110101; // iC=  309 
// vC = 14'b0000001100010011; // vC=  787 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000010; // iC=  450 
// vC = 14'b0000001101011011; // vC=  859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010101; // iC=  213 
// vC = 14'b0000001011011011; // vC=  731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101011; // iC=  363 
// vC = 14'b0000001101100101; // vC=  869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101010; // iC=  298 
// vC = 14'b0000001100100101; // vC=  805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010001; // iC=  401 
// vC = 14'b0000001011011001; // vC=  729 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111000; // iC=  248 
// vC = 14'b0000001100100110; // vC=  806 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100001; // iC=  161 
// vC = 14'b0000001010110001; // vC=  689 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101111; // iC=  431 
// vC = 14'b0000001001100011; // vC=  611 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011001; // iC=  409 
// vC = 14'b0000001100010100; // vC=  788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001110; // iC=  142 
// vC = 14'b0000001101111111; // vC=  895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101010; // iC=  170 
// vC = 14'b0000001100110011; // vC=  819 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111001; // iC=  185 
// vC = 14'b0000001101100000; // vC=  864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001011; // iC=  139 
// vC = 14'b0000001011110001; // vC=  753 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011011; // iC=  347 
// vC = 14'b0000001001110000; // vC=  624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011010; // iC=  282 
// vC = 14'b0000001100010100; // vC=  788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111000; // iC=  440 
// vC = 14'b0000001010000100; // vC=  644 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100100; // iC=  228 
// vC = 14'b0000001010111100; // vC=  700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000010; // iC=  322 
// vC = 14'b0000001101001001; // vC=  841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111000; // iC=  120 
// vC = 14'b0000001010101100; // vC=  684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010100; // iC=  212 
// vC = 14'b0000001101010001; // vC=  849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100010; // iC=  162 
// vC = 14'b0000001100100000; // vC=  800 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110110; // iC=  182 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000001; // iC=  257 
// vC = 14'b0000001101101011; // vC=  875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010111; // iC=  343 
// vC = 14'b0000001100100100; // vC=  804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110101; // iC=  181 
// vC = 14'b0000001110100100; // vC=  932 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000110; // iC=  262 
// vC = 14'b0000001100010101; // vC=  789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000111; // iC=  263 
// vC = 14'b0000001100101101; // vC=  813 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100101; // iC=  229 
// vC = 14'b0000001100010001; // vC=  785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110011; // iC=  115 
// vC = 14'b0000001010110000; // vC=  688 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010000; // iC=  336 
// vC = 14'b0000001010011011; // vC=  667 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000111; // iC=  263 
// vC = 14'b0000001001111100; // vC=  636 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000110; // iC=  134 
// vC = 14'b0000001101000011; // vC=  835 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000010; // iC=  130 
// vC = 14'b0000001110101010; // vC=  938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000111; // iC=  327 
// vC = 14'b0000001100101010; // vC=  810 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110111; // iC=  183 
// vC = 14'b0000001101011111; // vC=  863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001111; // iC=  271 
// vC = 14'b0000001011110011; // vC=  755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000111001; // iC=   57 
// vC = 14'b0000001010000011; // vC=  643 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001000110; // iC=   70 
// vC = 14'b0000001101101010; // vC=  874 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001110; // iC=  206 
// vC = 14'b0000001110100111; // vC=  935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000110; // iC=  134 
// vC = 14'b0000001101111111; // vC=  895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101011; // iC=  235 
// vC = 14'b0000001100001111; // vC=  783 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101011; // iC=  107 
// vC = 14'b0000001101000101; // vC=  837 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000111; // iC=  263 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100000; // iC=   32 
// vC = 14'b0000001010100101; // vC=  677 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111011; // iC=  187 
// vC = 14'b0000001010111100; // vC=  700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001110; // iC=   78 
// vC = 14'b0000001100100000; // vC=  800 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100000; // iC=  224 
// vC = 14'b0000001110011010; // vC=  922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010101; // iC=  213 
// vC = 14'b0000001101010110; // vC=  854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011101; // iC=  285 
// vC = 14'b0000001010111100; // vC=  700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000100; // iC=  260 
// vC = 14'b0000001010110100; // vC=  692 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001011; // iC=  331 
// vC = 14'b0000001100100010; // vC=  802 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101101; // iC=  109 
// vC = 14'b0000001011111100; // vC=  764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100111; // iC=   39 
// vC = 14'b0000001011000011; // vC=  707 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000100; // iC=  196 
// vC = 14'b0000001101000111; // vC=  839 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000001; // iC=  321 
// vC = 14'b0000001110001111; // vC=  911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101100; // iC=  300 
// vC = 14'b0000001010001101; // vC=  653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110001; // iC=  177 
// vC = 14'b0000001101011110; // vC=  862 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101111; // iC=  175 
// vC = 14'b0000001101010011; // vC=  851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110110; // iC=  246 
// vC = 14'b0000001011001100; // vC=  716 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100010; // iC=  162 
// vC = 14'b0000001110111001; // vC=  953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010101; // iC=   85 
// vC = 14'b0000001110101100; // vC=  940 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010000; // iC=  272 
// vC = 14'b0000001100101000; // vC=  808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001000011; // iC=   67 
// vC = 14'b0000001100011110; // vC=  798 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011001; // iC=   89 
// vC = 14'b0000001110010101; // vC=  917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110100; // iC=  180 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011001; // iC=   25 
// vC = 14'b0000001100010100; // vC=  788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011110; // iC=   30 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100101; // iC=  165 
// vC = 14'b0000001101110100; // vC=  884 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010000; // iC=  272 
// vC = 14'b0000001010011101; // vC=  669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110010; // iC=  114 
// vC = 14'b0000001100101000; // vC=  808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101010; // iC=  170 
// vC = 14'b0000001110111001; // vC=  953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101001; // iC=  -23 
// vC = 14'b0000001100110101; // vC=  821 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101100; // iC=  -20 
// vC = 14'b0000001100101110; // vC=  814 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010011; // iC=   83 
// vC = 14'b0000001010011010; // vC=  666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010101; // iC=  277 
// vC = 14'b0000001101001110; // vC=  846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100101; // iC=  101 
// vC = 14'b0000001100010101; // vC=  789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101110; // iC=  -18 
// vC = 14'b0000001101011101; // vC=  861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011110; // iC=  158 
// vC = 14'b0000001011101111; // vC=  751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100011; // iC=  163 
// vC = 14'b0000001010010011; // vC=  659 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100011; // iC=   35 
// vC = 14'b0000001101111000; // vC=  888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010011; // iC=  275 
// vC = 14'b0000001110100011; // vC=  931 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001001; // iC=    9 
// vC = 14'b0000001101100010; // vC=  866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001111; // iC=  271 
// vC = 14'b0000001110010101; // vC=  917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100100; // iC=  100 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001100; // iC=  204 
// vC = 14'b0000001010010111; // vC=  663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000110; // iC=  134 
// vC = 14'b0000001110000010; // vC=  898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100001; // iC=  -31 
// vC = 14'b0000001011001100; // vC=  716 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010001; // iC=   17 
// vC = 14'b0000001010001111; // vC=  655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101100; // iC=  236 
// vC = 14'b0000001101010001; // vC=  849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011101; // iC=   29 
// vC = 14'b0000001101111000; // vC=  888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000010; // iC=  258 
// vC = 14'b0000001011111001; // vC=  761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100111; // iC=   39 
// vC = 14'b0000001101111111; // vC=  895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001000; // iC=  264 
// vC = 14'b0000001110111101; // vC=  957 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000111011; // iC=   59 
// vC = 14'b0000001101110010; // vC=  882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011001; // iC=   89 
// vC = 14'b0000001010001101; // vC=  653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001000111; // iC=   71 
// vC = 14'b0000001010000110; // vC=  646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000110; // iC=  134 
// vC = 14'b0000001100101000; // vC=  808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010010; // iC=  146 
// vC = 14'b0000001100101111; // vC=  815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001110; // iC=  270 
// vC = 14'b0000001011110110; // vC=  758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101011; // iC=  -21 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000001; // iC=    1 
// vC = 14'b0000001011000111; // vC=  711 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001010; // iC=  266 
// vC = 14'b0000001010011111; // vC=  671 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011111; // iC=   95 
// vC = 14'b0000001101001110; // vC=  846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001100; // iC=   12 
// vC = 14'b0000001100010101; // vC=  789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011000; // iC=   88 
// vC = 14'b0000001101101111; // vC=  879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100010; // iC=  162 
// vC = 14'b0000001110010011; // vC=  915 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010000; // iC=   80 
// vC = 14'b0000001010101000; // vC=  680 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001111; // iC=  143 
// vC = 14'b0000001010010101; // vC=  661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000111; // iC=  199 
// vC = 14'b0000001010111000; // vC=  696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100010; // iC=  226 
// vC = 14'b0000001111010000; // vC=  976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101011; // iC=   43 
// vC = 14'b0000001101100000; // vC=  864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001011; // iC=  267 
// vC = 14'b0000001110011110; // vC=  926 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110111; // iC=  119 
// vC = 14'b0000001100000000; // vC=  768 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111011111; // iC=  -33 
// vC = 14'b0000001010110111; // vC=  695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100110; // iC=   38 
// vC = 14'b0000001110100000; // vC=  928 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101001; // iC=  169 
// vC = 14'b0000001010010000; // vC=  656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101110; // iC=  174 
// vC = 14'b0000001011001010; // vC=  714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000000; // iC=  192 
// vC = 14'b0000001101100010; // vC=  866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111000; // iC=  184 
// vC = 14'b0000001101011101; // vC=  861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000101; // iC=  261 
// vC = 14'b0000001100000010; // vC=  770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101010; // iC=  106 
// vC = 14'b0000001100100011; // vC=  803 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100110; // iC=  -26 
// vC = 14'b0000001011100101; // vC=  741 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000110001; // iC=   49 
// vC = 14'b0000001100100100; // vC=  804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001010; // iC=   74 
// vC = 14'b0000001101100000; // vC=  864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001011; // iC=   75 
// vC = 14'b0000001011100100; // vC=  740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011010; // iC=   26 
// vC = 14'b0000001010111001; // vC=  697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010011; // iC=   83 
// vC = 14'b0000001011010111; // vC=  727 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010001; // iC=   17 
// vC = 14'b0000001010011011; // vC=  667 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000110000; // iC=   48 
// vC = 14'b0000001010101100; // vC=  684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011001; // iC=   89 
// vC = 14'b0000001110101100; // vC=  940 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000011; // iC=    3 
// vC = 14'b0000001011000110; // vC=  710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101011; // iC=  107 
// vC = 14'b0000001011101010; // vC=  746 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011110; // iC=  286 
// vC = 14'b0000001101110010; // vC=  882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001011; // iC=  203 
// vC = 14'b0000001110111110; // vC=  958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100010; // iC=  290 
// vC = 14'b0000001101001101; // vC=  845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011101; // iC=  157 
// vC = 14'b0000001111001100; // vC=  972 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011011; // iC=   91 
// vC = 14'b0000001101101100; // vC=  876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011011110; // iC=  222 
// vC = 14'b0000001011011111; // vC=  735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000111; // iC=  135 
// vC = 14'b0000001111000110; // vC=  966 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010110; // iC=  278 
// vC = 14'b0000001100010001; // vC=  785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101000; // iC=  296 
// vC = 14'b0000001011101101; // vC=  749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001110; // iC=   14 
// vC = 14'b0000001101100100; // vC=  868 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001100; // iC=  332 
// vC = 14'b0000001010011010; // vC=  666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000110; // iC=  326 
// vC = 14'b0000001110011010; // vC=  922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111000; // iC=  184 
// vC = 14'b0000001100011011; // vC=  795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110110; // iC=  246 
// vC = 14'b0000001100000010; // vC=  770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111101; // iC=  253 
// vC = 14'b0000001101011101; // vC=  861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001000; // iC=  264 
// vC = 14'b0000001111010000; // vC=  976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101010; // iC=   42 
// vC = 14'b0000001100100100; // vC=  804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111000; // iC=  184 
// vC = 14'b0000001011101011; // vC=  747 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001010; // iC=  202 
// vC = 14'b0000001111011001; // vC=  985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100001; // iC=  353 
// vC = 14'b0000001101000001; // vC=  833 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010011; // iC=  211 
// vC = 14'b0000001011111000; // vC=  760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100000; // iC=  352 
// vC = 14'b0000001110111101; // vC=  957 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001000011; // iC=   67 
// vC = 14'b0000001110000111; // vC=  903 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110001; // iC=  369 
// vC = 14'b0000001011111001; // vC=  761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011101; // iC=   93 
// vC = 14'b0000001011101001; // vC=  745 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110000; // iC=  240 
// vC = 14'b0000001110101111; // vC=  943 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101001; // iC=  169 
// vC = 14'b0000001010110001; // vC=  689 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000110; // iC=  134 
// vC = 14'b0000001100000100; // vC=  772 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011111; // iC=   95 
// vC = 14'b0000001111011111; // vC=  991 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100100; // iC=  100 
// vC = 14'b0000001110010000; // vC=  912 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101010; // iC=  234 
// vC = 14'b0000001110100101; // vC=  933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001011; // iC=  203 
// vC = 14'b0000001110110100; // vC=  948 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001010; // iC=  394 
// vC = 14'b0000001101011011; // vC=  859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111100; // iC=  124 
// vC = 14'b0000001110001001; // vC=  905 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111110; // iC=  126 
// vC = 14'b0000001111010010; // vC=  978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110110; // iC=  118 
// vC = 14'b0000001110101111; // vC=  943 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100010; // iC=  418 
// vC = 14'b0000001011011001; // vC=  729 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011111; // iC=  415 
// vC = 14'b0000001110010000; // vC=  912 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001110; // iC=  142 
// vC = 14'b0000001010110010; // vC=  690 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100010; // iC=  418 
// vC = 14'b0000001110110011; // vC=  947 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011110; // iC=  350 
// vC = 14'b0000001100101000; // vC=  808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111111; // iC=  127 
// vC = 14'b0000001011101111; // vC=  751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111000; // iC=  376 
// vC = 14'b0000001011110101; // vC=  757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010101; // iC=  149 
// vC = 14'b0000001111010110; // vC=  982 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000001; // iC=  449 
// vC = 14'b0000001011001101; // vC=  717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110011; // iC=  243 
// vC = 14'b0000001111010011; // vC=  979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111100; // iC=  188 
// vC = 14'b0000001100011000; // vC=  792 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000110; // iC=  198 
// vC = 14'b0000001111000111; // vC=  967 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110000; // iC=  368 
// vC = 14'b0000001110001000; // vC=  904 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101100; // iC=  364 
// vC = 14'b0000001101111111; // vC=  895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000001; // iC=  257 
// vC = 14'b0000001110011111; // vC=  927 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000001; // iC=  385 
// vC = 14'b0000001011011000; // vC=  728 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001011; // iC=  203 
// vC = 14'b0000001100010000; // vC=  784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000100; // iC=  388 
// vC = 14'b0000001101101101; // vC=  877 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001100; // iC=  396 
// vC = 14'b0000001111011100; // vC=  988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111100; // iC=  316 
// vC = 14'b0000001101000111; // vC=  839 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000110; // iC=  454 
// vC = 14'b0000001111001111; // vC=  975 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100101; // iC=  357 
// vC = 14'b0000001110110011; // vC=  947 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011011; // iC=  411 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100100; // iC=  420 
// vC = 14'b0000010000000100; // vC= 1028 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111001; // iC=  313 
// vC = 14'b0000001110101010; // vC=  938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010101; // iC=  213 
// vC = 14'b0000001110100100; // vC=  932 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000000; // iC=  448 
// vC = 14'b0000001011100001; // vC=  737 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111101; // iC=  317 
// vC = 14'b0000001101010101; // vC=  853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000101; // iC=  517 
// vC = 14'b0000001111101101; // vC= 1005 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001011; // iC=  267 
// vC = 14'b0000010000000101; // vC= 1029 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011011; // iC=  475 
// vC = 14'b0000001111001100; // vC=  972 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110111; // iC=  375 
// vC = 14'b0000001110000001; // vC=  897 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111001; // iC=  505 
// vC = 14'b0000001100101101; // vC=  813 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011110; // iC=  350 
// vC = 14'b0000001110011100; // vC=  924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100100; // iC=  548 
// vC = 14'b0000001100111101; // vC=  829 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011110; // iC=  414 
// vC = 14'b0000001011011110; // vC=  734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110010; // iC=  306 
// vC = 14'b0000001110101010; // vC=  938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110000; // iC=  304 
// vC = 14'b0000001111100110; // vC=  998 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101011; // iC=  299 
// vC = 14'b0000001110010101; // vC=  917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110100; // iC=  372 
// vC = 14'b0000001101000000; // vC=  832 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100000; // iC=  608 
// vC = 14'b0000001100010100; // vC=  788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110001; // iC=  305 
// vC = 14'b0000001101010101; // vC=  853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001100; // iC=  524 
// vC = 14'b0000001100110111; // vC=  823 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001010; // iC=  458 
// vC = 14'b0000001111010001; // vC=  977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011010; // iC=  346 
// vC = 14'b0000001100001111; // vC=  783 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000100; // iC=  452 
// vC = 14'b0000010000100101; // vC= 1061 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100110; // iC=  550 
// vC = 14'b0000001111010100; // vC=  980 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000101; // iC=  645 
// vC = 14'b0000001100000000; // vC=  768 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011100; // iC=  412 
// vC = 14'b0000001110001110; // vC=  910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010111; // iC=  407 
// vC = 14'b0000001101111101; // vC=  893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111011; // iC=  635 
// vC = 14'b0000010000010000; // vC= 1040 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101100; // iC=  556 
// vC = 14'b0000001110011010; // vC=  922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111001; // iC=  505 
// vC = 14'b0000001100111001; // vC=  825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110110; // iC=  502 
// vC = 14'b0000001111001010; // vC=  970 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011000; // iC=  408 
// vC = 14'b0000001100000100; // vC=  772 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011010; // iC=  410 
// vC = 14'b0000001101111111; // vC=  895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111011; // iC=  379 
// vC = 14'b0000010000110000; // vC= 1072 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001001; // iC=  585 
// vC = 14'b0000001110011001; // vC=  921 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111111; // iC=  575 
// vC = 14'b0000010000001101; // vC= 1037 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100000; // iC=  416 
// vC = 14'b0000010000010111; // vC= 1047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100101; // iC=  485 
// vC = 14'b0000001111001110; // vC=  974 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100110; // iC=  486 
// vC = 14'b0000010000010001; // vC= 1041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000011; // iC=  515 
// vC = 14'b0000001110100001; // vC=  929 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110111; // iC=  695 
// vC = 14'b0000001111000001; // vC=  961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000010; // iC=  514 
// vC = 14'b0000001111001111; // vC=  975 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011010; // iC=  666 
// vC = 14'b0000001111001110; // vC=  974 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010100; // iC=  532 
// vC = 14'b0000001110011001; // vC=  921 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110101; // iC=  565 
// vC = 14'b0000010000111111; // vC= 1087 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000000; // iC=  704 
// vC = 14'b0000010000110010; // vC= 1074 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000010; // iC=  706 
// vC = 14'b0000001101101001; // vC=  873 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001111; // iC=  591 
// vC = 14'b0000010001001111; // vC= 1103 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011001; // iC=  665 
// vC = 14'b0000001101101110; // vC=  878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110010; // iC=  626 
// vC = 14'b0000010001011001; // vC= 1113 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000100; // iC=  644 
// vC = 14'b0000001101011000; // vC=  856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000111; // iC=  519 
// vC = 14'b0000010000000001; // vC= 1025 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110101; // iC=  693 
// vC = 14'b0000010000110000; // vC= 1072 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010100; // iC=  596 
// vC = 14'b0000010000100110; // vC= 1062 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100101; // iC=  613 
// vC = 14'b0000001101100010; // vC=  866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010010; // iC=  722 
// vC = 14'b0000010001101010; // vC= 1130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101011; // iC=  555 
// vC = 14'b0000001111110001; // vC= 1009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000100; // iC=  708 
// vC = 14'b0000010000010011; // vC= 1043 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010001; // iC=  529 
// vC = 14'b0000001111100101; // vC=  997 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101001; // iC=  681 
// vC = 14'b0000001111011011; // vC=  987 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001101; // iC=  717 
// vC = 14'b0000001111101111; // vC= 1007 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010110; // iC=  598 
// vC = 14'b0000001111111111; // vC= 1023 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110111; // iC=  823 
// vC = 14'b0000001111011111; // vC=  991 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001011; // iC=  715 
// vC = 14'b0000010010000101; // vC= 1157 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001110; // iC=  590 
// vC = 14'b0000001111111001; // vC= 1017 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010011; // iC=  723 
// vC = 14'b0000001111101001; // vC= 1001 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010001; // iC=  657 
// vC = 14'b0000010010000001; // vC= 1153 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011101; // iC=  669 
// vC = 14'b0000001111000010; // vC=  962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b0000010010000010; // vC= 1154 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100110; // iC=  806 
// vC = 14'b0000001111001001; // vC=  969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101000; // iC=  680 
// vC = 14'b0000001110111001; // vC=  953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000000; // iC=  704 
// vC = 14'b0000010000110001; // vC= 1073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101111; // iC=  815 
// vC = 14'b0000001110011010; // vC=  922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001100; // iC=  780 
// vC = 14'b0000010010011110; // vC= 1182 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111011; // iC=  635 
// vC = 14'b0000010000010000; // vC= 1040 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000011; // iC=  707 
// vC = 14'b0000001101101110; // vC=  878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001000; // iC=  712 
// vC = 14'b0000010000111100; // vC= 1084 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111000; // iC=  824 
// vC = 14'b0000010010110001; // vC= 1201 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101011; // iC=  811 
// vC = 14'b0000010000110001; // vC= 1073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000101; // iC=  709 
// vC = 14'b0000001110010101; // vC=  917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100000; // iC=  672 
// vC = 14'b0000001111110111; // vC= 1015 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001001; // iC=  841 
// vC = 14'b0000001110111111; // vC=  959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011000; // iC=  920 
// vC = 14'b0000010010010010; // vC= 1170 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111111; // iC=  767 
// vC = 14'b0000010001000010; // vC= 1090 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010100; // iC=  724 
// vC = 14'b0000010001011011; // vC= 1115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000001; // iC=  705 
// vC = 14'b0000010010011001; // vC= 1177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000010; // iC=  962 
// vC = 14'b0000010001011000; // vC= 1112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000110; // iC=  966 
// vC = 14'b0000001111110010; // vC= 1010 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100000; // iC=  800 
// vC = 14'b0000010001010000; // vC= 1104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100011; // iC=  931 
// vC = 14'b0000010001011010; // vC= 1114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100111; // iC=  743 
// vC = 14'b0000010000110001; // vC= 1073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101111; // iC=  879 
// vC = 14'b0000010001101000; // vC= 1128 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111111; // iC=  703 
// vC = 14'b0000001111011011; // vC=  987 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010100; // iC=  980 
// vC = 14'b0000001111000000; // vC=  960 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011011; // iC=  859 
// vC = 14'b0000010000001101; // vC= 1037 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011100; // iC=  924 
// vC = 14'b0000010001101010; // vC= 1130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111110; // iC=  894 
// vC = 14'b0000001111100111; // vC=  999 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111010; // iC=  762 
// vC = 14'b0000010011110011; // vC= 1267 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111100; // iC=  828 
// vC = 14'b0000001111000011; // vC=  963 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100011; // iC=  803 
// vC = 14'b0000010001001000; // vC= 1096 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110111; // iC=  887 
// vC = 14'b0000010001001011; // vC= 1099 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010010; // iC=  978 
// vC = 14'b0000010011000011; // vC= 1219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000011; // iC= 1027 
// vC = 14'b0000010001111100; // vC= 1148 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011001; // iC=  793 
// vC = 14'b0000010001001011; // vC= 1099 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000100; // iC=  900 
// vC = 14'b0000010011001001; // vC= 1225 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000100; // iC= 1028 
// vC = 14'b0000010001001010; // vC= 1098 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010010; // iC= 1042 
// vC = 14'b0000010000101010; // vC= 1066 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000101; // iC=  901 
// vC = 14'b0000010001110101; // vC= 1141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110001; // iC= 1073 
// vC = 14'b0000010011101011; // vC= 1259 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011111; // iC=  799 
// vC = 14'b0000010010010100; // vC= 1172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111000; // iC=  952 
// vC = 14'b0000010011101000; // vC= 1256 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000110; // iC=  966 
// vC = 14'b0000010000101001; // vC= 1065 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000110; // iC=  966 
// vC = 14'b0000010100100100; // vC= 1316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111000; // iC=  888 
// vC = 14'b0000010011100111; // vC= 1255 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101001; // iC=  937 
// vC = 14'b0000001111111000; // vC= 1016 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101100; // iC= 1004 
// vC = 14'b0000010010001000; // vC= 1160 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011111; // iC=  927 
// vC = 14'b0000010100100111; // vC= 1319 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010001; // iC= 1041 
// vC = 14'b0000010100111101; // vC= 1341 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100001; // iC=  929 
// vC = 14'b0000010010001100; // vC= 1164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001000; // iC= 1096 
// vC = 14'b0000010001010001; // vC= 1105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011011; // iC= 1051 
// vC = 14'b0000010010011010; // vC= 1178 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101001; // iC=  873 
// vC = 14'b0000010010101111; // vC= 1199 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010010; // iC=  914 
// vC = 14'b0000010101001101; // vC= 1357 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100011; // iC= 1123 
// vC = 14'b0000010100011111; // vC= 1311 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100111; // iC=  871 
// vC = 14'b0000010100000001; // vC= 1281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101101; // iC=  941 
// vC = 14'b0000010100000010; // vC= 1282 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111010; // iC= 1082 
// vC = 14'b0000010011010010; // vC= 1234 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110001; // iC= 1009 
// vC = 14'b0000010101100110; // vC= 1382 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010001; // iC=  977 
// vC = 14'b0000010000110010; // vC= 1074 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011110; // iC=  926 
// vC = 14'b0000010001111000; // vC= 1144 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110001; // iC=  945 
// vC = 14'b0000010010101111; // vC= 1199 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000111; // iC= 1031 
// vC = 14'b0000010101101110; // vC= 1390 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111000; // iC= 1080 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010100; // iC=  852 
// vC = 14'b0000010100111110; // vC= 1342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011001; // iC=  921 
// vC = 14'b0000010001101000; // vC= 1128 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010000; // iC=  912 
// vC = 14'b0000010101100000; // vC= 1376 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111000; // iC= 1016 
// vC = 14'b0000010101111011; // vC= 1403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000100; // iC=  964 
// vC = 14'b0000010011101111; // vC= 1263 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111011; // iC= 1083 
// vC = 14'b0000010110010010; // vC= 1426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110010; // iC= 1074 
// vC = 14'b0000010100000111; // vC= 1287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000000; // iC= 1088 
// vC = 14'b0000010100111000; // vC= 1336 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111011; // iC=  891 
// vC = 14'b0000010110100110; // vC= 1446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101000; // iC=  936 
// vC = 14'b0000010101100110; // vC= 1382 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111001; // iC= 1145 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111000; // iC= 1016 
// vC = 14'b0000010110001011; // vC= 1419 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010011; // iC= 1107 
// vC = 14'b0000010100111010; // vC= 1338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010111; // iC= 1111 
// vC = 14'b0000010001111111; // vC= 1151 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111001; // iC= 1017 
// vC = 14'b0000010100101101; // vC= 1325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011100; // iC= 1052 
// vC = 14'b0000010010111011; // vC= 1211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000110; // iC=  966 
// vC = 14'b0000010011010000; // vC= 1232 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001011; // iC= 1035 
// vC = 14'b0000010011101110; // vC= 1262 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100000; // iC= 1056 
// vC = 14'b0000010110100010; // vC= 1442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101000; // iC=  936 
// vC = 14'b0000010010110100; // vC= 1204 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010101; // iC= 1109 
// vC = 14'b0000010011000101; // vC= 1221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000001; // iC=  961 
// vC = 14'b0000010100101101; // vC= 1325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100000; // iC= 1184 
// vC = 14'b0000010101111100; // vC= 1404 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011110; // iC= 1054 
// vC = 14'b0000010011111000; // vC= 1272 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110000; // iC= 1136 
// vC = 14'b0000010110101001; // vC= 1449 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011000; // iC= 1112 
// vC = 14'b0000010101000100; // vC= 1348 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001001; // iC= 1225 
// vC = 14'b0000010110111110; // vC= 1470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110011; // iC= 1203 
// vC = 14'b0000010101000011; // vC= 1347 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000111; // iC=  967 
// vC = 14'b0000010111010110; // vC= 1494 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001011; // iC= 1163 
// vC = 14'b0000010110100001; // vC= 1441 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000111; // iC= 1031 
// vC = 14'b0000010100111100; // vC= 1340 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010010; // iC= 1106 
// vC = 14'b0000010111010001; // vC= 1489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100000; // iC=  992 
// vC = 14'b0000010011010000; // vC= 1232 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001110; // iC=  974 
// vC = 14'b0000010110001111; // vC= 1423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001100; // iC=  972 
// vC = 14'b0000010100111100; // vC= 1340 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100011; // iC=  931 
// vC = 14'b0000010100111011; // vC= 1339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010010; // iC=  978 
// vC = 14'b0000010011101101; // vC= 1261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000110; // iC= 1222 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110011; // iC= 1139 
// vC = 14'b0000010110001111; // vC= 1423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101110; // iC= 1134 
// vC = 14'b0000010100111011; // vC= 1339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011111; // iC=  991 
// vC = 14'b0000011000000101; // vC= 1541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011010; // iC= 1178 
// vC = 14'b0000010101001101; // vC= 1357 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001110; // iC= 1166 
// vC = 14'b0000010110111100; // vC= 1468 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110110; // iC= 1078 
// vC = 14'b0000010100100010; // vC= 1314 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101010; // iC= 1066 
// vC = 14'b0000011000010000; // vC= 1552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000111; // iC= 1159 
// vC = 14'b0000010110100110; // vC= 1446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111000; // iC= 1208 
// vC = 14'b0000011000100001; // vC= 1569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010000; // iC= 1232 
// vC = 14'b0000011000101011; // vC= 1579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110001; // iC= 1009 
// vC = 14'b0000011000000100; // vC= 1540 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100110; // iC= 1126 
// vC = 14'b0000010111010111; // vC= 1495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110011; // iC= 1075 
// vC = 14'b0000010111110000; // vC= 1520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110001; // iC=  945 
// vC = 14'b0000011000010011; // vC= 1555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100101; // iC= 1189 
// vC = 14'b0000010101111011; // vC= 1403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111100; // iC= 1084 
// vC = 14'b0000010110110011; // vC= 1459 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010100; // iC= 1044 
// vC = 14'b0000010101000001; // vC= 1345 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011100; // iC= 1116 
// vC = 14'b0000010110101100; // vC= 1452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101100; // iC= 1196 
// vC = 14'b0000010110101000; // vC= 1448 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000111; // iC= 1031 
// vC = 14'b0000010101000110; // vC= 1350 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001011; // iC= 1227 
// vC = 14'b0000010111011100; // vC= 1500 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101000; // iC= 1064 
// vC = 14'b0000011001010010; // vC= 1618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010100; // iC= 1172 
// vC = 14'b0000011000110100; // vC= 1588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100010; // iC= 1186 
// vC = 14'b0000011000001100; // vC= 1548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101010; // iC= 1194 
// vC = 14'b0000011001110000; // vC= 1648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011001; // iC= 1241 
// vC = 14'b0000010110111100; // vC= 1468 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001010; // iC= 1034 
// vC = 14'b0000010111001110; // vC= 1486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100101; // iC=  997 
// vC = 14'b0000011001011101; // vC= 1629 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011100; // iC= 1116 
// vC = 14'b0000010110110000; // vC= 1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100111; // iC= 1127 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000001; // iC= 1089 
// vC = 14'b0000010110101010; // vC= 1450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101000; // iC= 1000 
// vC = 14'b0000011000001101; // vC= 1549 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011111; // iC=  991 
// vC = 14'b0000011001000011; // vC= 1603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010011; // iC=  915 
// vC = 14'b0000011010000111; // vC= 1671 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001011; // iC=  971 
// vC = 14'b0000010110011000; // vC= 1432 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010110; // iC= 1174 
// vC = 14'b0000011001010000; // vC= 1616 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110110; // iC= 1078 
// vC = 14'b0000011010010111; // vC= 1687 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100100; // iC= 1060 
// vC = 14'b0000011001010100; // vC= 1620 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101011; // iC= 1195 
// vC = 14'b0000010111001010; // vC= 1482 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011101; // iC= 1181 
// vC = 14'b0000011011010001; // vC= 1745 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101000; // iC= 1128 
// vC = 14'b0000011010111110; // vC= 1726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000001; // iC= 1153 
// vC = 14'b0000011001010011; // vC= 1619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110001; // iC= 1201 
// vC = 14'b0000011001001100; // vC= 1612 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101101; // iC= 1005 
// vC = 14'b0000011000111110; // vC= 1598 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100011; // iC= 1187 
// vC = 14'b0000011001001110; // vC= 1614 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011000; // iC= 1048 
// vC = 14'b0000011001010111; // vC= 1623 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011001; // iC= 1049 
// vC = 14'b0000010111101010; // vC= 1514 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001000; // iC=  968 
// vC = 14'b0000010110110011; // vC= 1459 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101011; // iC= 1067 
// vC = 14'b0000011011000101; // vC= 1733 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000101; // iC= 1157 
// vC = 14'b0000011001011010; // vC= 1626 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110000; // iC= 1136 
// vC = 14'b0000011001101001; // vC= 1641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011110; // iC= 1054 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101101; // iC= 1133 
// vC = 14'b0000011001000100; // vC= 1604 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101100; // iC=  940 
// vC = 14'b0000011001111100; // vC= 1660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100010; // iC= 1058 
// vC = 14'b0000011100001101; // vC= 1805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100001; // iC= 1185 
// vC = 14'b0000011000101011; // vC= 1579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111000; // iC=  888 
// vC = 14'b0000011000010100; // vC= 1556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101000; // iC= 1064 
// vC = 14'b0000011001111100; // vC= 1660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101001; // iC= 1129 
// vC = 14'b0000011000110111; // vC= 1591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011010; // iC= 1114 
// vC = 14'b0000011010100000; // vC= 1696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010010; // iC= 1042 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011011; // iC=  987 
// vC = 14'b0000011010001001; // vC= 1673 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000011; // iC=  899 
// vC = 14'b0000011010000000; // vC= 1664 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111010; // iC= 1146 
// vC = 14'b0000011000001001; // vC= 1545 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000101; // iC=  965 
// vC = 14'b0000010111111000; // vC= 1528 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000010; // iC= 1154 
// vC = 14'b0000011000111101; // vC= 1597 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011110; // iC=  990 
// vC = 14'b0000011010100010; // vC= 1698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111000; // iC=  952 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111100; // iC=  892 
// vC = 14'b0000011000011101; // vC= 1565 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100101; // iC= 1061 
// vC = 14'b0000011011010001; // vC= 1745 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111011; // iC=  827 
// vC = 14'b0000011100000110; // vC= 1798 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000011; // iC=  835 
// vC = 14'b0000011100110100; // vC= 1844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100011; // iC=  867 
// vC = 14'b0000011011110101; // vC= 1781 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010101; // iC= 1045 
// vC = 14'b0000011101001010; // vC= 1866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111011; // iC=  955 
// vC = 14'b0000011100001111; // vC= 1807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011011; // iC= 1115 
// vC = 14'b0000011100101011; // vC= 1835 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111001; // iC= 1081 
// vC = 14'b0000011010100110; // vC= 1702 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110010; // iC=  946 
// vC = 14'b0000011011110001; // vC= 1777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000000; // iC= 1088 
// vC = 14'b0000011011110000; // vC= 1776 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000000; // iC=  832 
// vC = 14'b0000011100001110; // vC= 1806 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010001; // iC=  849 
// vC = 14'b0000011000111110; // vC= 1598 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001011; // iC=  907 
// vC = 14'b0000011011110110; // vC= 1782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010110; // iC=  854 
// vC = 14'b0000011011100100; // vC= 1764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000110; // iC=  774 
// vC = 14'b0000011100011010; // vC= 1818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001111; // iC=  847 
// vC = 14'b0000011101100011; // vC= 1891 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001101; // iC=  845 
// vC = 14'b0000011011110001; // vC= 1777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110000; // iC= 1008 
// vC = 14'b0000011001101100; // vC= 1644 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111111; // iC=  959 
// vC = 14'b0000011001101100; // vC= 1644 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010000; // iC=  848 
// vC = 14'b0000011101111101; // vC= 1917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001001; // iC=  969 
// vC = 14'b0000011010001111; // vC= 1679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100100; // iC=  932 
// vC = 14'b0000011001101011; // vC= 1643 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011111; // iC=  927 
// vC = 14'b0000011101010001; // vC= 1873 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100000; // iC=  736 
// vC = 14'b0000011101001110; // vC= 1870 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110100; // iC=  756 
// vC = 14'b0000011110101001; // vC= 1961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110011; // iC=  947 
// vC = 14'b0000011101000100; // vC= 1860 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000111; // iC=  967 
// vC = 14'b0000011110010000; // vC= 1936 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001100; // iC=  972 
// vC = 14'b0000011100100110; // vC= 1830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100101; // iC=  741 
// vC = 14'b0000011100111000; // vC= 1848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111011; // iC=  763 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101110; // iC= 1006 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110000; // iC=  752 
// vC = 14'b0000011010001101; // vC= 1677 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110011; // iC=  755 
// vC = 14'b0000011110111101; // vC= 1981 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011101; // iC=  989 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000000; // iC=  896 
// vC = 14'b0000011111001000; // vC= 1992 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010101; // iC=  725 
// vC = 14'b0000011100011010; // vC= 1818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b0000011100110101; // vC= 1845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101010; // iC=  874 
// vC = 14'b0000011110111011; // vC= 1979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110101; // iC=  949 
// vC = 14'b0000011110010101; // vC= 1941 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101100; // iC=  812 
// vC = 14'b0000011111000000; // vC= 1984 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111101; // iC=  701 
// vC = 14'b0000011101111011; // vC= 1915 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100110; // iC=  678 
// vC = 14'b0000011110100110; // vC= 1958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111010; // iC=  954 
// vC = 14'b0000011110110111; // vC= 1975 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010000; // iC=  848 
// vC = 14'b0000011010110011; // vC= 1715 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000110; // iC=  710 
// vC = 14'b0000011101011001; // vC= 1881 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010011; // iC=  787 
// vC = 14'b0000011011110010; // vC= 1778 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100100; // iC=  676 
// vC = 14'b0000011111100100; // vC= 2020 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100101; // iC=  677 
// vC = 14'b0000011100101111; // vC= 1839 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011111; // iC=  671 
// vC = 14'b0000011011010001; // vC= 1745 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110100; // iC=  628 
// vC = 14'b0000011011001001; // vC= 1737 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000010; // iC=  770 
// vC = 14'b0000011100001100; // vC= 1804 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010010; // iC=  786 
// vC = 14'b0000011011010011; // vC= 1747 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101111; // iC=  879 
// vC = 14'b0000011011101011; // vC= 1771 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010010; // iC=  786 
// vC = 14'b0000011111110110; // vC= 2038 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010111; // iC=  727 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111111; // iC=  895 
// vC = 14'b0000011101100110; // vC= 1894 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101111; // iC=  815 
// vC = 14'b0000011011111001; // vC= 1785 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100000; // iC=  672 
// vC = 14'b0000011111100110; // vC= 2022 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110010; // iC=  626 
// vC = 14'b0000011100101010; // vC= 1834 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100110; // iC=  550 
// vC = 14'b0000011101011110; // vC= 1886 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000001; // iC=  833 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111101; // iC=  701 
// vC = 14'b0000011111110111; // vC= 2039 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010010; // iC=  786 
// vC = 14'b0000011110101010; // vC= 1962 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001010; // iC=  586 
// vC = 14'b0000011100011000; // vC= 1816 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011011; // iC=  731 
// vC = 14'b0000011101111010; // vC= 1914 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010011; // iC=  595 
// vC = 14'b0000011110010000; // vC= 1936 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010001; // iC=  593 
// vC = 14'b0000011101110101; // vC= 1909 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010111; // iC=  535 
// vC = 14'b0000011110111001; // vC= 1977 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100001; // iC=  545 
// vC = 14'b0000011111100000; // vC= 2016 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111001; // iC=  505 
// vC = 14'b0000011101110100; // vC= 1908 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001001; // iC=  649 
// vC = 14'b0000011110001011; // vC= 1931 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110111; // iC=  567 
// vC = 14'b0000011011110111; // vC= 1783 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011110; // iC=  606 
// vC = 14'b0000100000001010; // vC= 2058 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011011; // iC=  475 
// vC = 14'b0000011111110001; // vC= 2033 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101101; // iC=  493 
// vC = 14'b0000011110011001; // vC= 1945 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001000; // iC=  648 
// vC = 14'b0000011110000011; // vC= 1923 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111011; // iC=  379 
// vC = 14'b0000011110001101; // vC= 1933 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010011; // iC=  403 
// vC = 14'b0000011100011101; // vC= 1821 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111011; // iC=  571 
// vC = 14'b0000100000001001; // vC= 2057 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011000; // iC=  408 
// vC = 14'b0000011101011010; // vC= 1882 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110000; // iC=  304 
// vC = 14'b0000011110010100; // vC= 1940 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010010; // iC=  594 
// vC = 14'b0000011100101010; // vC= 1834 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110110; // iC=  374 
// vC = 14'b0000011100101111; // vC= 1839 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111011; // iC=  379 
// vC = 14'b0000100000000010; // vC= 2050 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001011; // iC=  523 
// vC = 14'b0000100001001100; // vC= 2124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111011; // iC=  251 
// vC = 14'b0000011101011010; // vC= 1882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000011; // iC=  515 
// vC = 14'b0000011111011000; // vC= 2008 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011010; // iC=  410 
// vC = 14'b0000100000101100; // vC= 2092 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101011; // iC=  235 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011111; // iC=  415 
// vC = 14'b0000011111101011; // vC= 2027 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001100; // iC=  460 
// vC = 14'b0000011111101011; // vC= 2027 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100001; // iC=  289 
// vC = 14'b0000100000010100; // vC= 2068 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111011; // iC=  443 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001010; // iC=  394 
// vC = 14'b0000011110000111; // vC= 1927 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001110; // iC=  334 
// vC = 14'b0000011111001100; // vC= 1996 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001100; // iC=  268 
// vC = 14'b0000011101100001; // vC= 1889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100000; // iC=  224 
// vC = 14'b0000011101101100; // vC= 1900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101001; // iC=  233 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100000; // iC=   96 
// vC = 14'b0000011101110001; // vC= 1905 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111001; // iC=  249 
// vC = 14'b0000011100111000; // vC= 1848 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010101; // iC=  213 
// vC = 14'b0000011110101100; // vC= 1964 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101000; // iC=   40 
// vC = 14'b0000011111000010; // vC= 1986 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011111; // iC=  287 
// vC = 14'b0000011100111001; // vC= 1849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100110; // iC=  102 
// vC = 14'b0000011110010010; // vC= 1938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001000; // iC=    8 
// vC = 14'b0000100000111001; // vC= 2105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000000; // iC=  128 
// vC = 14'b0000100000011101; // vC= 2077 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001010; // iC=   10 
// vC = 14'b0000011100011111; // vC= 1823 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000000; // iC=  192 
// vC = 14'b0000011101111110; // vC= 1918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011110; // iC=  -98 
// vC = 14'b0000011110100010; // vC= 1954 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101011; // iC=   43 
// vC = 14'b0000011101110100; // vC= 1908 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000010; // iC= -126 
// vC = 14'b0000011111010001; // vC= 2001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100001; // iC=   97 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001110; // iC= -178 
// vC = 14'b0000011101001001; // vC= 1865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000010; // iC= -126 
// vC = 14'b0000011111110110; // vC= 2038 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011110010; // iC= -270 
// vC = 14'b0000011111110101; // vC= 2037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000100; // iC= -124 
// vC = 14'b0000100000010011; // vC= 2067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011100101; // iC= -283 
// vC = 14'b0000100001010010; // vC= 2130 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101010; // iC=  -22 
// vC = 14'b0000100001001111; // vC= 2127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100010; // iC= -158 
// vC = 14'b0000011100010010; // vC= 1810 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010000; // iC= -176 
// vC = 14'b0000011111101100; // vC= 2028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100101; // iC= -347 
// vC = 14'b0000100000110100; // vC= 2100 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001001; // iC= -119 
// vC = 14'b0000011100101001; // vC= 1833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101010; // iC= -406 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110000; // iC= -400 
// vC = 14'b0000100000001000; // vC= 2056 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111001; // iC= -327 
// vC = 14'b0000011101000110; // vC= 1862 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001110; // iC= -370 
// vC = 14'b0000011111101100; // vC= 2028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001001; // iC= -439 
// vC = 14'b0000100000001100; // vC= 2060 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100011; // iC= -413 
// vC = 14'b0000011100011011; // vC= 1819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101111; // iC= -465 
// vC = 14'b0000011110111011; // vC= 1979 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011111; // iC= -481 
// vC = 14'b0000011101010011; // vC= 1875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011101; // iC= -483 
// vC = 14'b0000011110001010; // vC= 1930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000110; // iC= -570 
// vC = 14'b0000011110011101; // vC= 1949 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101011; // iC= -533 
// vC = 14'b0000100000000011; // vC= 2051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111001; // iC= -647 
// vC = 14'b0000011101111111; // vC= 1919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111111; // iC= -641 
// vC = 14'b0000011101001000; // vC= 1864 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010001; // iC= -623 
// vC = 14'b0000011111010000; // vC= 2000 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001000; // iC= -440 
// vC = 14'b0000011101011000; // vC= 1880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111000; // iC= -648 
// vC = 14'b0000011110101101; // vC= 1965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011100; // iC= -548 
// vC = 14'b0000011101101001; // vC= 1897 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100111; // iC= -537 
// vC = 14'b0000011011101001; // vC= 1769 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011111; // iC= -673 
// vC = 14'b0000011011011110; // vC= 1758 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110111; // iC= -649 
// vC = 14'b0000011110001011; // vC= 1931 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111110; // iC= -834 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010100; // iC= -748 
// vC = 14'b0000011100110011; // vC= 1843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100001; // iC= -671 
// vC = 14'b0000011100001101; // vC= 1805 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011001; // iC= -871 
// vC = 14'b0000011110001101; // vC= 1933 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101011; // iC= -597 
// vC = 14'b0000011111000100; // vC= 1988 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111000; // iC= -776 
// vC = 14'b0000011100001110; // vC= 1806 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101000; // iC= -792 
// vC = 14'b0000011101100001; // vC= 1889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000101; // iC= -827 
// vC = 14'b0000011110011001; // vC= 1945 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011000; // iC= -744 
// vC = 14'b0000011011011101; // vC= 1757 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101011; // iC= -981 
// vC = 14'b0000011011010111; // vC= 1751 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101010; // iC= -854 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101001; // iC= -727 
// vC = 14'b0000011110101111; // vC= 1967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111010; // iC= -774 
// vC = 14'b0000011011001110; // vC= 1742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100011; // iC= -861 
// vC = 14'b0000011100010111; // vC= 1815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111110; // iC= -898 
// vC = 14'b0000011010111101; // vC= 1725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000101; // iC=-1083 
// vC = 14'b0000011110111011; // vC= 1979 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100010; // iC= -990 
// vC = 14'b0000011110000100; // vC= 1924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001000; // iC= -824 
// vC = 14'b0000011011101000; // vC= 1768 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000010; // iC=-1086 
// vC = 14'b0000011010101011; // vC= 1707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101000; // iC= -920 
// vC = 14'b0000011010011001; // vC= 1689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001011; // iC=-1013 
// vC = 14'b0000011110111001; // vC= 1977 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001101; // iC= -947 
// vC = 14'b0000011101011100; // vC= 1884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010100; // iC=-1132 
// vC = 14'b0000011101010100; // vC= 1876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b0000011010011000; // vC= 1688 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011001; // iC=-1127 
// vC = 14'b0000011110010011; // vC= 1939 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111111; // iC=-1025 
// vC = 14'b0000011110000001; // vC= 1921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100100; // iC=-1052 
// vC = 14'b0000011110101010; // vC= 1962 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001101; // iC=-1139 
// vC = 14'b0000011101010011; // vC= 1875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000001; // iC=-1279 
// vC = 14'b0000011101101001; // vC= 1897 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010100; // iC=-1132 
// vC = 14'b0000011010001110; // vC= 1678 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010101; // iC=-1131 
// vC = 14'b0000011101100110; // vC= 1894 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101011; // iC=-1045 
// vC = 14'b0000011011100000; // vC= 1760 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110001; // iC=-1231 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001011; // iC=-1077 
// vC = 14'b0000011110000000; // vC= 1920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110111; // iC=-1353 
// vC = 14'b0000011101010010; // vC= 1874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010110; // iC=-1130 
// vC = 14'b0000011001111100; // vC= 1660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101100; // iC=-1236 
// vC = 14'b0000011001001111; // vC= 1615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101001; // iC=-1303 
// vC = 14'b0000011001001000; // vC= 1608 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000001; // iC=-1407 
// vC = 14'b0000011011001011; // vC= 1739 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010110; // iC=-1194 
// vC = 14'b0000011011010110; // vC= 1750 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110100; // iC=-1292 
// vC = 14'b0000011100011011; // vC= 1819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101101; // iC=-1427 
// vC = 14'b0000011100111000; // vC= 1848 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110001; // iC=-1359 
// vC = 14'b0000011000101001; // vC= 1577 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111100; // iC=-1348 
// vC = 14'b0000011011110011; // vC= 1779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101000; // iC=-1176 
// vC = 14'b0000011011100000; // vC= 1760 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010011; // iC=-1453 
// vC = 14'b0000011011000000; // vC= 1728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111001; // iC=-1351 
// vC = 14'b0000011000110001; // vC= 1585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111010; // iC=-1414 
// vC = 14'b0000011001110101; // vC= 1653 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010011; // iC=-1453 
// vC = 14'b0000010111110000; // vC= 1520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000100; // iC=-1532 
// vC = 14'b0000011000010100; // vC= 1556 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001101; // iC=-1395 
// vC = 14'b0000011011011011; // vC= 1755 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111101; // iC=-1539 
// vC = 14'b0000011011001110; // vC= 1742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101110; // iC=-1554 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000111; // iC=-1401 
// vC = 14'b0000011000011111; // vC= 1567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011101; // iC=-1571 
// vC = 14'b0000011001000000; // vC= 1600 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111010; // iC=-1350 
// vC = 14'b0000011010101011; // vC= 1707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011100; // iC=-1380 
// vC = 14'b0000011000011010; // vC= 1562 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101110; // iC=-1490 
// vC = 14'b0000011010101101; // vC= 1709 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110000; // iC=-1552 
// vC = 14'b0000011011010011; // vC= 1747 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010100; // iC=-1516 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101010; // iC=-1302 
// vC = 14'b0000010111100010; // vC= 1506 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000101; // iC=-1595 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110100; // iC=-1420 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101010; // iC=-1430 
// vC = 14'b0000011010000100; // vC= 1668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011000; // iC=-1640 
// vC = 14'b0000010110010000; // vC= 1424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001010; // iC=-1334 
// vC = 14'b0000010110001101; // vC= 1421 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010011; // iC=-1581 
// vC = 14'b0000010110010100; // vC= 1428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000011; // iC=-1533 
// vC = 14'b0000011001111101; // vC= 1661 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011110; // iC=-1442 
// vC = 14'b0000010110111011; // vC= 1467 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000000; // iC=-1664 
// vC = 14'b0000010110110000; // vC= 1456 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111011; // iC=-1477 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011011; // iC=-1445 
// vC = 14'b0000010111110001; // vC= 1521 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011010; // iC=-1702 
// vC = 14'b0000010101011111; // vC= 1375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010101; // iC=-1515 
// vC = 14'b0000010111101001; // vC= 1513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110110; // iC=-1610 
// vC = 14'b0000010110011101; // vC= 1437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101111; // iC=-1617 
// vC = 14'b0000010111101100; // vC= 1516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011110; // iC=-1506 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111001; // iC=-1543 
// vC = 14'b0000011000010110; // vC= 1558 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001011; // iC=-1653 
// vC = 14'b0000011001011100; // vC= 1628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110101; // iC=-1675 
// vC = 14'b0000010110111001; // vC= 1465 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100010; // iC=-1694 
// vC = 14'b0000010111011001; // vC= 1497 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011001; // iC=-1447 
// vC = 14'b0000011001010001; // vC= 1617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011010; // iC=-1510 
// vC = 14'b0000010100001100; // vC= 1292 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101010; // iC=-1686 
// vC = 14'b0000010100101111; // vC= 1327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101110; // iC=-1618 
// vC = 14'b0000010100111011; // vC= 1339 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010011; // iC=-1773 
// vC = 14'b0000010100010001; // vC= 1297 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110101; // iC=-1483 
// vC = 14'b0000010111101100; // vC= 1516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000010; // iC=-1470 
// vC = 14'b0000010111101000; // vC= 1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110010; // iC=-1486 
// vC = 14'b0000011000011010; // vC= 1562 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110001; // iC=-1807 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110100; // iC=-1548 
// vC = 14'b0000010110001001; // vC= 1417 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000001; // iC=-1599 
// vC = 14'b0000010011110100; // vC= 1268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111011; // iC=-1605 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100001; // iC=-1503 
// vC = 14'b0000010101101100; // vC= 1388 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011000; // iC=-1640 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100001; // iC=-1567 
// vC = 14'b0000010110111111; // vC= 1471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000011; // iC=-1725 
// vC = 14'b0000010101011100; // vC= 1372 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b0000010011110010; // vC= 1266 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000100; // iC=-1596 
// vC = 14'b0000010110000001; // vC= 1409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011001; // iC=-1703 
// vC = 14'b0000010101010010; // vC= 1362 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111000; // iC=-1672 
// vC = 14'b0000010011001111; // vC= 1231 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101110; // iC=-1810 
// vC = 14'b0000010101100000; // vC= 1376 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100100; // iC=-1628 
// vC = 14'b0000010011101101; // vC= 1261 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000101; // iC=-1787 
// vC = 14'b0000010011100101; // vC= 1253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001001; // iC=-1655 
// vC = 14'b0000010100100000; // vC= 1312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100001; // iC=-1759 
// vC = 14'b0000010011110001; // vC= 1265 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011010; // iC=-1702 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000000; // iC=-1664 
// vC = 14'b0000010001010111; // vC= 1111 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010010; // iC=-1646 
// vC = 14'b0000010001111001; // vC= 1145 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000111; // iC=-1913 
// vC = 14'b0000010001010010; // vC= 1106 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111110; // iC=-1794 
// vC = 14'b0000010100101010; // vC= 1322 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b0000010101010001; // vC= 1361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111010; // iC=-1734 
// vC = 14'b0000010011111111; // vC= 1279 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111011; // iC=-1669 
// vC = 14'b0000010100001000; // vC= 1288 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b0000010010000111; // vC= 1159 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b0000010001110000; // vC= 1136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b0000010000111011; // vC= 1083 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011111; // iC=-1761 
// vC = 14'b0000010011001101; // vC= 1229 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b0000010000010011; // vC= 1043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111100; // iC=-1732 
// vC = 14'b0000010100110010; // vC= 1330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b0000010011011001; // vC= 1241 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001110; // iC=-1906 
// vC = 14'b0000010010100100; // vC= 1188 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b0000010011101110; // vC= 1262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111110; // iC=-1666 
// vC = 14'b0000010001100011; // vC= 1123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111110; // iC=-1730 
// vC = 14'b0000010010010011; // vC= 1171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100111; // iC=-1753 
// vC = 14'b0000010001100001; // vC= 1121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b0000010011110100; // vC= 1268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b0000010010010101; // vC= 1173 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100111; // iC=-1945 
// vC = 14'b0000010001110111; // vC= 1143 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100111; // iC=-1945 
// vC = 14'b0000010011001010; // vC= 1226 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001011; // iC=-1781 
// vC = 14'b0000010000110011; // vC= 1075 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000010; // iC=-1726 
// vC = 14'b0000010000001010; // vC= 1034 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110000; // iC=-1936 
// vC = 14'b0000010010100000; // vC= 1184 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111100; // iC=-1796 
// vC = 14'b0000010000110111; // vC= 1079 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b0000010000111110; // vC= 1086 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b0000001110000111; // vC=  903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b0000001110001110; // vC=  910 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b0000001111101100; // vC= 1004 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b0000010001010101; // vC= 1109 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001011; // iC=-1973 
// vC = 14'b0000001110101010; // vC=  938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000110; // iC=-1850 
// vC = 14'b0000010001010111; // vC= 1111 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b0000001101100011; // vC=  867 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b0000001100111110; // vC=  830 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000101; // iC=-2043 
// vC = 14'b0000001111101001; // vC= 1001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b0000001101000001; // vC=  833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b0000010000100000; // vC= 1056 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000010000111010; // vC= 1082 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b0000001110011000; // vC=  920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000001111000000; // vC=  960 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100011; // iC=-1821 
// vC = 14'b0000010000100010; // vC= 1058 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b0000001100001001; // vC=  777 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100111; // iC=-1881 
// vC = 14'b0000001111101011; // vC= 1003 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b0000001011101101; // vC=  749 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b0000001101000011; // vC=  835 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000010000001101; // vC= 1037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000001110000111; // vC=  903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100101; // iC=-2075 
// vC = 14'b0000001110111111; // vC=  959 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000011; // iC=-1981 
// vC = 14'b0000001100000011; // vC=  771 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000011; // iC=-1853 
// vC = 14'b0000001010111101; // vC=  701 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000001110000010; // vC=  898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b0000001010011100; // vC=  668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b0000001100101110; // vC=  814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110011; // iC=-1933 
// vC = 14'b0000001010110110; // vC=  694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b0000001111000111; // vC=  967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100010; // iC=-2142 
// vC = 14'b0000001101001001; // vC=  841 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000001100111010; // vC=  826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000101; // iC=-1851 
// vC = 14'b0000001101110100; // vC=  884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000001101101111; // vC=  879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000111; // iC=-1913 
// vC = 14'b0000001100010010; // vC=  786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000001110001100; // vC=  908 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b0000001001001010; // vC=  586 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100010; // iC=-1886 
// vC = 14'b0000001101001011; // vC=  843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111001; // iC=-2119 
// vC = 14'b0000001010100011; // vC=  675 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b0000001100001111; // vC=  783 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000001001001101; // vC=  589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b0000001010000111; // vC=  647 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111111; // iC=-1921 
// vC = 14'b0000001011011110; // vC=  734 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011111; // iC=-2081 
// vC = 14'b0000001010000111; // vC=  647 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011111; // iC=-1953 
// vC = 14'b0000001011011101; // vC=  733 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000110; // iC=-2170 
// vC = 14'b0000001100100100; // vC=  804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110110; // iC=-2186 
// vC = 14'b0000001001101111; // vC=  623 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000001001011101; // vC=  605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011100; // iC=-2148 
// vC = 14'b0000001000010101; // vC=  533 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b0000001011101100; // vC=  748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b0000001010110010; // vC=  690 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111100; // iC=-2180 
// vC = 14'b0000001001110101; // vC=  629 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000000110111111; // vC=  447 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000001010110100; // vC=  692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000011; // iC=-2173 
// vC = 14'b0000001000111010; // vC=  570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111011; // iC=-2117 
// vC = 14'b0000001010110100; // vC=  692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101010; // iC=-2198 
// vC = 14'b0000001001000000; // vC=  576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111110; // iC=-2242 
// vC = 14'b0000001000111001; // vC=  569 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b0000001001000110; // vC=  582 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000100; // iC=-2236 
// vC = 14'b0000000101111011; // vC=  379 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101010; // iC=-2198 
// vC = 14'b0000000110101101; // vC=  429 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101101; // iC=-2259 
// vC = 14'b0000000101110010; // vC=  370 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010101; // iC=-2091 
// vC = 14'b0000001000101000; // vC=  552 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101101; // iC=-2131 
// vC = 14'b0000001010001011; // vC=  651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101010; // iC=-2134 
// vC = 14'b0000000111001010; // vC=  458 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b0000001001110111; // vC=  631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b0000001001110010; // vC=  626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000000111011000; // vC=  472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101011; // iC=-2133 
// vC = 14'b0000000100101111; // vC=  303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b0000001000011110; // vC=  542 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000011; // iC=-2173 
// vC = 14'b0000001000111010; // vC=  570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010100; // iC=-2156 
// vC = 14'b0000000101101101; // vC=  365 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010111; // iC=-2217 
// vC = 14'b0000000111111110; // vC=  510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111001; // iC=-2183 
// vC = 14'b0000000100011110; // vC=  286 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000000110111011; // vC=  443 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110001; // iC=-2127 
// vC = 14'b0000000101000010; // vC=  322 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000000011110000; // vC=  240 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110001; // iC=-2127 
// vC = 14'b0000000100100001; // vC=  289 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011100; // iC=-2212 
// vC = 14'b0000000111101000; // vC=  488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001101; // iC=-2163 
// vC = 14'b0000000011011100; // vC=  220 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011111; // iC=-2081 
// vC = 14'b0000000011111101; // vC=  253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010100; // iC=-2092 
// vC = 14'b0000000100000000; // vC=  256 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101101; // iC=-2131 
// vC = 14'b0000000111100010; // vC=  482 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010001; // iC=-2223 
// vC = 14'b0000000101100111; // vC=  359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110101; // iC=-2251 
// vC = 14'b0000000010011011; // vC=  155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010001; // iC=-2223 
// vC = 14'b0000000101011001; // vC=  345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111001; // iC=-2183 
// vC = 14'b0000000011011011; // vC=  219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111001; // iC=-2119 
// vC = 14'b0000000110110011; // vC=  435 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011011000; // iC=-2344 
// vC = 14'b0000000100100000; // vC=  288 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011111; // iC=-2209 
// vC = 14'b0000000110000001; // vC=  385 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011111111; // iC=-2305 
// vC = 14'b0000000001010101; // vC=   85 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000111; // iC=-2233 
// vC = 14'b0000000100111100; // vC=  316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100001110; // iC=-2290 
// vC = 14'b0000000100100101; // vC=  293 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100001010; // iC=-2294 
// vC = 14'b0000000001110001; // vC=  113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011011000; // iC=-2344 
// vC = 14'b0000000010100010; // vC=  162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b0000000100111001; // vC=  313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100000; // iC=-2208 
// vC = 14'b0000000010001011; // vC=  139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000001; // iC=-2239 
// vC = 14'b0000000100111100; // vC=  316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111110; // iC=-2050 
// vC = 14'b0000000011110000; // vC=  240 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011010101; // iC=-2347 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011010111; // iC=-2345 
// vC = 14'b0000000010011001; // vC=  153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010100; // iC=-2220 
// vC = 14'b0000000011010001; // vC=  209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011011100; // iC=-2340 
// vC = 14'b1111111111110111; // vC=   -9 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011101100; // iC=-2324 
// vC = 14'b0000000010000101; // vC=  133 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101100; // iC=-2196 
// vC = 14'b1111111111100110; // vC=  -26 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011100111; // iC=-2329 
// vC = 14'b0000000010110011; // vC=  179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100000100; // iC=-2300 
// vC = 14'b0000000011001111; // vC=  207 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011000011; // iC=-2365 
// vC = 14'b1111111111011000; // vC=  -40 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011000110; // iC=-2362 
// vC = 14'b0000000000011111; // vC=   31 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100100; // iC=-2204 
// vC = 14'b0000000010011011; // vC=  155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001000; // iC=-2232 
// vC = 14'b0000000010000100; // vC=  132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100001; // iC=-2143 
// vC = 14'b0000000000110010; // vC=   50 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000111; // iC=-2105 
// vC = 14'b0000000000000100; // vC=    4 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001100; // iC=-2228 
// vC = 14'b1111111110011010; // vC= -102 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100011011; // iC=-2277 
// vC = 14'b0000000001001101; // vC=   77 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010111000; // iC=-2376 
// vC = 14'b1111111101110011; // vC= -141 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010000; // iC=-2224 
// vC = 14'b1111111101111000; // vC= -136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011100; // iC=-2212 
// vC = 14'b0000000001100011; // vC=   99 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111001; // iC=-2119 
// vC = 14'b1111111101001111; // vC= -177 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011101111; // iC=-2321 
// vC = 14'b0000000001101001; // vC=  105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000001; // iC=-2239 
// vC = 14'b0000000000001010; // vC=   10 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011100; // iC=-2212 
// vC = 14'b1111111111000111; // vC=  -57 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100111; // iC=-2201 
// vC = 14'b0000000001000000; // vC=   64 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011010110; // iC=-2346 
// vC = 14'b1111111101100000; // vC= -160 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100100; // iC=-2204 
// vC = 14'b1111111110000000; // vC= -128 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011111; // iC=-2145 
// vC = 14'b1111111100111111; // vC= -193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101000; // iC=-2200 
// vC = 14'b0000000000010100; // vC=   20 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111001; // iC=-2119 
// vC = 14'b1111111111001010; // vC=  -54 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b1111111100111101; // vC= -195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100011111; // iC=-2273 
// vC = 14'b1111111111011010; // vC=  -38 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010011011; // iC=-2405 
// vC = 14'b1111111100101110; // vC= -210 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100111; // iC=-2137 
// vC = 14'b1111111110101011; // vC=  -85 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110101; // iC=-2123 
// vC = 14'b1111111111101110; // vC=  -18 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111100; // iC=-2180 
// vC = 14'b1111111111011100; // vC=  -36 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110101; // iC=-2187 
// vC = 14'b1111111100000101; // vC= -251 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000101; // iC=-2171 
// vC = 14'b1111111010111001; // vC= -327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100001110; // iC=-2290 
// vC = 14'b1111111111001100; // vC=  -52 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011001; // iC=-2215 
// vC = 14'b1111111010101011; // vC= -341 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010001110; // iC=-2418 
// vC = 14'b1111111010110010; // vC= -334 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010010110; // iC=-2410 
// vC = 14'b1111111101001100; // vC= -180 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001101; // iC=-2227 
// vC = 14'b1111111010100110; // vC= -346 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011010; // iC=-2214 
// vC = 14'b1111111010100011; // vC= -349 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100110; // iC=-2138 
// vC = 14'b1111111011100110; // vC= -282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011101011; // iC=-2325 
// vC = 14'b1111111011100011; // vC= -285 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101001; // iC=-2199 
// vC = 14'b1111111011101110; // vC= -274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010001; // iC=-2223 
// vC = 14'b1111111001111110; // vC= -386 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010100000; // iC=-2400 
// vC = 14'b1111111010000111; // vC= -377 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100011110; // iC=-2274 
// vC = 14'b1111111100000011; // vC= -253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011011; // iC=-2149 
// vC = 14'b1111111011110110; // vC= -266 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010010011; // iC=-2413 
// vC = 14'b1111111101000010; // vC= -190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010101; // iC=-2219 
// vC = 14'b1111111001101101; // vC= -403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b1111111100001010; // vC= -246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011001001; // iC=-2359 
// vC = 14'b1111111010010111; // vC= -361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011100101; // iC=-2331 
// vC = 14'b1111111011001111; // vC= -305 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011101010; // iC=-2326 
// vC = 14'b1111111100110011; // vC= -205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010110111; // iC=-2377 
// vC = 14'b1111111001101110; // vC= -402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101001; // iC=-2135 
// vC = 14'b1111111011000100; // vC= -316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010111; // iC=-2217 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111110; // iC=-2242 
// vC = 14'b1111111011100111; // vC= -281 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011101; // iC=-2211 
// vC = 14'b1111111010010100; // vC= -364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011010101; // iC=-2347 
// vC = 14'b1111111000110001; // vC= -463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011010; // iC=-2214 
// vC = 14'b1111111010100100; // vC= -348 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001001; // iC=-2231 
// vC = 14'b1111111010110011; // vC= -333 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011001001; // iC=-2359 
// vC = 14'b1111111000111001; // vC= -455 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011100001; // iC=-2335 
// vC = 14'b1111110111011110; // vC= -546 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010011000; // iC=-2408 
// vC = 14'b1111111000001100; // vC= -500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010111110; // iC=-2370 
// vC = 14'b1111111000110111; // vC= -457 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000111; // iC=-2169 
// vC = 14'b1111110111001000; // vC= -568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011100011; // iC=-2333 
// vC = 14'b1111111010101101; // vC= -339 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101010; // iC=-2262 
// vC = 14'b1111111010011101; // vC= -355 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010110010; // iC=-2382 
// vC = 14'b1111111000111000; // vC= -456 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110011; // iC=-2253 
// vC = 14'b1111110111100000; // vC= -544 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010101100; // iC=-2388 
// vC = 14'b1111110110000010; // vC= -638 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110111; // iC=-2249 
// vC = 14'b1111111001000101; // vC= -443 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100011101; // iC=-2275 
// vC = 14'b1111110111111000; // vC= -520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100001001; // iC=-2295 
// vC = 14'b1111111000011011; // vC= -485 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010100111; // iC=-2393 
// vC = 14'b1111111001001011; // vC= -437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100100101; // iC=-2267 
// vC = 14'b1111110111011000; // vC= -552 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000010; // iC=-2238 
// vC = 14'b1111110110100111; // vC= -601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001100; // iC=-2228 
// vC = 14'b1111110100110000; // vC= -720 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111101; // iC=-2179 
// vC = 14'b1111110110100010; // vC= -606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100101; // iC=-2203 
// vC = 14'b1111110110011001; // vC= -615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100100110; // iC=-2266 
// vC = 14'b1111110110010101; // vC= -619 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110111; // iC=-2121 
// vC = 14'b1111110101001111; // vC= -689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000100; // iC=-2172 
// vC = 14'b1111110111000010; // vC= -574 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000100; // iC=-2172 
// vC = 14'b1111110101010000; // vC= -688 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011100000; // iC=-2336 
// vC = 14'b1111110011001110; // vC= -818 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111011; // iC=-2181 
// vC = 14'b1111110100110010; // vC= -718 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010011001; // iC=-2407 
// vC = 14'b1111110110011110; // vC= -610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100010000; // iC=-2288 
// vC = 14'b1111110101001111; // vC= -689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011101001; // iC=-2327 
// vC = 14'b1111110110010110; // vC= -618 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011010000; // iC=-2352 
// vC = 14'b1111110110111011; // vC= -581 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010111110; // iC=-2370 
// vC = 14'b1111110010100001; // vC= -863 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110100; // iC=-2188 
// vC = 14'b1111110010111011; // vC= -837 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110110; // iC=-2186 
// vC = 14'b1111110101000111; // vC= -697 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100001; // iC=-2207 
// vC = 14'b1111110100000110; // vC= -762 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011001; // iC=-2087 
// vC = 14'b1111110010101010; // vC= -854 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110110; // iC=-2122 
// vC = 14'b1111110100100100; // vC= -732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011001000; // iC=-2360 
// vC = 14'b1111110101110111; // vC= -649 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b1111110101011011; // vC= -677 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011101; // iC=-2211 
// vC = 14'b1111110011000110; // vC= -826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101001; // iC=-2263 
// vC = 14'b1111110011101110; // vC= -786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011000100; // iC=-2364 
// vC = 14'b1111110010110001; // vC= -847 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001100; // iC=-2164 
// vC = 14'b1111110001001001; // vC= -951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111000; // iC=-2120 
// vC = 14'b1111110010011011; // vC= -869 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100011101; // iC=-2275 
// vC = 14'b1111110101000001; // vC= -703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101100; // iC=-2132 
// vC = 14'b1111110001111011; // vC= -901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001000; // iC=-2168 
// vC = 14'b1111110100001101; // vC= -755 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011011; // iC=-2085 
// vC = 14'b1111110001001100; // vC= -948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011101101; // iC=-2323 
// vC = 14'b1111110010111110; // vC= -834 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101001; // iC=-2135 
// vC = 14'b1111110010101111; // vC= -849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011010110111; // iC=-2377 
// vC = 14'b1111110001100101; // vC= -923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011001; // iC=-2087 
// vC = 14'b1111110011001011; // vC= -821 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110101; // iC=-2123 
// vC = 14'b1111101111010110; // vC=-1066 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110111; // iC=-2249 
// vC = 14'b1111110010100010; // vC= -862 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b1111110001101010; // vC= -918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001010; // iC=-2230 
// vC = 14'b1111101111011100; // vC=-1060 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010110; // iC=-2218 
// vC = 14'b1111101111000111; // vC=-1081 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b1111110010100011; // vC= -861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111100; // iC=-2116 
// vC = 14'b1111110010100011; // vC= -861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001000; // iC=-2232 
// vC = 14'b1111101110000100; // vC=-1148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b1111101111100101; // vC=-1051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111000; // iC=-2056 
// vC = 14'b1111101101101101; // vC=-1171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011010111; // iC=-2345 
// vC = 14'b1111110000000000; // vC=-1024 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011010010; // iC=-2350 
// vC = 14'b1111101111011001; // vC=-1063 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010001; // iC=-2095 
// vC = 14'b1111110000000011; // vC=-1021 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011101; // iC=-2147 
// vC = 14'b1111101111000000; // vC=-1088 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010100; // iC=-2156 
// vC = 14'b1111110001111001; // vC= -903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011001; // iC=-2151 
// vC = 14'b1111101101010000; // vC=-1200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100000011; // iC=-2301 
// vC = 14'b1111101100111110; // vC=-1218 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011100011; // iC=-2333 
// vC = 14'b1111101110011010; // vC=-1126 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100011011; // iC=-2277 
// vC = 14'b1111101111110001; // vC=-1039 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b1111101110000100; // vC=-1148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011011110111; // iC=-2313 
// vC = 14'b1111101110100011; // vC=-1117 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101010; // iC=-2262 
// vC = 14'b1111110000001111; // vC=-1009 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011100; // iC=-2212 
// vC = 14'b1111101110100101; // vC=-1115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110001; // iC=-2063 
// vC = 14'b1111101111110011; // vC=-1037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111000; // iC=-2056 
// vC = 14'b1111101101100110; // vC=-1178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101100; // iC=-2132 
// vC = 14'b1111101111110100; // vC=-1036 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110111; // iC=-2185 
// vC = 14'b1111101111101001; // vC=-1047 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b1111101100010101; // vC=-1259 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110100; // iC=-2252 
// vC = 14'b1111101011000100; // vC=-1340 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100000; // iC=-2080 
// vC = 14'b1111101110111001; // vC=-1095 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b1111101101001101; // vC=-1203 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010101; // iC=-2027 
// vC = 14'b1111101110010111; // vC=-1129 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100010100; // iC=-2284 
// vC = 14'b1111101011100011; // vC=-1309 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b1111101011110110; // vC=-1290 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011010; // iC=-2214 
// vC = 14'b1111101001111111; // vC=-1409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100001; // iC=-2079 
// vC = 14'b1111101011011011; // vC=-1317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110001; // iC=-1999 
// vC = 14'b1111101100101110; // vC=-1234 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101001; // iC=-2199 
// vC = 14'b1111101001111011; // vC=-1413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100010001; // iC=-2287 
// vC = 14'b1111101110001101; // vC=-1139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101001; // iC=-2263 
// vC = 14'b1111101010101110; // vC=-1362 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b1111101100110100; // vC=-1228 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111011; // iC=-2117 
// vC = 14'b1111101100101001; // vC=-1239 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100001110; // iC=-2290 
// vC = 14'b1111101101111101; // vC=-1155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b1111101001100011; // vC=-1437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110010; // iC=-2062 
// vC = 14'b1111101100000111; // vC=-1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b1111101000101011; // vC=-1493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b1111101000110100; // vC=-1484 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011011; // iC=-2213 
// vC = 14'b1111101000110000; // vC=-1488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100101; // iC=-2011 
// vC = 14'b1111101100011010; // vC=-1254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b1111101011001011; // vC=-1333 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011001; // iC=-2151 
// vC = 14'b1111101000110000; // vC=-1488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b1111101001000000; // vC=-1472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b1111101011111000; // vC=-1288 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111000; // iC=-2248 
// vC = 14'b1111101011010010; // vC=-1326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b1111101000011010; // vC=-1510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b1111101001110101; // vC=-1419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110001; // iC=-2063 
// vC = 14'b1111100111111101; // vC=-1539 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000111; // iC=-2169 
// vC = 14'b1111100111011011; // vC=-1573 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011100; // iC=-2212 
// vC = 14'b1111101000101100; // vC=-1492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001100; // iC=-2228 
// vC = 14'b1111101000011101; // vC=-1507 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101101; // iC=-2195 
// vC = 14'b1111101010001001; // vC=-1399 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010110; // iC=-2090 
// vC = 14'b1111101011000011; // vC=-1341 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101010; // iC=-2198 
// vC = 14'b1111101001110011; // vC=-1421 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b1111101001010111; // vC=-1449 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b1111101000110001; // vC=-1487 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110011; // iC=-1997 
// vC = 14'b1111101010101110; // vC=-1362 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101111; // iC=-2001 
// vC = 14'b1111101010011111; // vC=-1377 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100111; // iC=-1945 
// vC = 14'b1111100101011100; // vC=-1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100011; // iC=-2077 
// vC = 14'b1111100101110010; // vC=-1678 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b1111100101001111; // vC=-1713 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000100; // iC=-2172 
// vC = 14'b1111100111101000; // vC=-1560 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b1111100110010110; // vC=-1642 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b1111100110000101; // vC=-1659 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b1111100100111011; // vC=-1733 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b1111100111111010; // vC=-1542 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000110; // iC=-1978 
// vC = 14'b1111100100111110; // vC=-1730 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000101; // iC=-1915 
// vC = 14'b1111100100011100; // vC=-1764 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010100; // iC=-1900 
// vC = 14'b1111100101011101; // vC=-1699 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111111; // iC=-1985 
// vC = 14'b1111101000101010; // vC=-1494 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001111; // iC=-2161 
// vC = 14'b1111101000100110; // vC=-1498 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001110; // iC=-1906 
// vC = 14'b1111100111010111; // vC=-1577 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b1111100110010100; // vC=-1644 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111100; // iC=-1860 
// vC = 14'b1111100111010101; // vC=-1579 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b1111100101101000; // vC=-1688 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101000; // iC=-2136 
// vC = 14'b1111100100011011; // vC=-1765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b1111100101010110; // vC=-1706 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b1111100111000001; // vC=-1599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011111; // iC=-2081 
// vC = 14'b1111100100011101; // vC=-1763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b1111100011010110; // vC=-1834 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b1111100010101111; // vC=-1873 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011001; // iC=-2087 
// vC = 14'b1111100110110101; // vC=-1611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110011; // iC=-1933 
// vC = 14'b1111100010101110; // vC=-1874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b1111100110101010; // vC=-1622 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011011; // iC=-1829 
// vC = 14'b1111100010011110; // vC=-1890 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b1111100010000010; // vC=-1918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110100; // iC=-2060 
// vC = 14'b1111100010010100; // vC=-1900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b1111100101100100; // vC=-1692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b1111100011100111; // vC=-1817 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b1111100101011010; // vC=-1702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b1111100101010100; // vC=-1708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011011; // iC=-1829 
// vC = 14'b1111100101101101; // vC=-1683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011001; // iC=-1895 
// vC = 14'b1111100001011101; // vC=-1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000011; // iC=-1853 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b1111100101111001; // vC=-1671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b1111100000101111; // vC=-2001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101010; // iC=-1878 
// vC = 14'b1111100010101101; // vC=-1875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100111; // iC=-1881 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b1111100011101101; // vC=-1811 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b1111100100111010; // vC=-1734 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b1111100000011001; // vC=-2023 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b1111100000011100; // vC=-2020 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b1111100010110111; // vC=-1865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001010; // iC=-1782 
// vC = 14'b1111100001010011; // vC=-1965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b1111100100100110; // vC=-1754 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b1111100010010010; // vC=-1902 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010100; // iC=-1772 
// vC = 14'b1111100010100011; // vC=-1885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b1111100011010111; // vC=-1833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010110; // iC=-1770 
// vC = 14'b1111100000010011; // vC=-2029 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110001; // iC=-1999 
// vC = 14'b1111011111000011; // vC=-2109 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b1111100001101011; // vC=-1941 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100110; // iC=-1690 
// vC = 14'b1111100000111110; // vC=-1986 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b1111100000001000; // vC=-2040 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b1111100011001101; // vC=-1843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b1111100000110110; // vC=-1994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001011; // iC=-1717 
// vC = 14'b1111100001110000; // vC=-1936 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111000; // iC=-1736 
// vC = 14'b1111100000101111; // vC=-2001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100101; // iC=-1755 
// vC = 14'b1111100010000001; // vC=-1919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b1111011110100000; // vC=-2144 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100010; // iC=-1694 
// vC = 14'b1111011110111111; // vC=-2113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000111; // iC=-1913 
// vC = 14'b1111100000101110; // vC=-2002 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111100000011001; // vC=-2023 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011010; // iC=-1894 
// vC = 14'b1111011101111001; // vC=-2183 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b1111100000001111; // vC=-2033 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011000; // iC=-1640 
// vC = 14'b1111011111001110; // vC=-2098 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000010; // iC=-1726 
// vC = 14'b1111100000111000; // vC=-1992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110100; // iC=-1932 
// vC = 14'b1111011110111110; // vC=-2114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110000; // iC=-1616 
// vC = 14'b1111011110000010; // vC=-2174 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101100; // iC=-1684 
// vC = 14'b1111011110100010; // vC=-2142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101000; // iC=-1880 
// vC = 14'b1111011111001000; // vC=-2104 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000111; // iC=-1913 
// vC = 14'b1111011111011010; // vC=-2086 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000010; // iC=-1598 
// vC = 14'b1111011100110100; // vC=-2252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101111; // iC=-1745 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100101; // iC=-1755 
// vC = 14'b1111100000001000; // vC=-2040 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b1111011110000101; // vC=-2171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110111; // iC=-1609 
// vC = 14'b1111011100001011; // vC=-2293 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000011; // iC=-1853 
// vC = 14'b1111011110001011; // vC=-2165 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b1111011111000111; // vC=-2105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100001; // iC=-1695 
// vC = 14'b1111011101011100; // vC=-2212 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001011; // iC=-1781 
// vC = 14'b1111011110110001; // vC=-2127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010100; // iC=-1772 
// vC = 14'b1111011110000001; // vC=-2175 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101101; // iC=-1683 
// vC = 14'b1111011111000111; // vC=-2105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011110; // iC=-1698 
// vC = 14'b1111011101101011; // vC=-2197 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111000; // iC=-1608 
// vC = 14'b1111011011100011; // vC=-2333 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110011; // iC=-1549 
// vC = 14'b1111011101001101; // vC=-2227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001101; // iC=-1523 
// vC = 14'b1111011100110011; // vC=-2253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010101; // iC=-1643 
// vC = 14'b1111011101010101; // vC=-2219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111010; // iC=-1670 
// vC = 14'b1111011100101010; // vC=-2262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000111; // iC=-1657 
// vC = 14'b1111011101000011; // vC=-2237 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111011; // iC=-1669 
// vC = 14'b1111011100010101; // vC=-2283 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000110; // iC=-1722 
// vC = 14'b1111011100010111; // vC=-2281 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111101; // iC=-1603 
// vC = 14'b1111011010010110; // vC=-2410 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110001; // iC=-1679 
// vC = 14'b1111011100011110; // vC=-2274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111001; // iC=-1735 
// vC = 14'b1111011101010011; // vC=-2221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111101; // iC=-1475 
// vC = 14'b1111011100011111; // vC=-2273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111000; // iC=-1608 
// vC = 14'b1111011010111011; // vC=-2373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110010; // iC=-1614 
// vC = 14'b1111011101100100; // vC=-2204 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111010; // iC=-1478 
// vC = 14'b1111011101011010; // vC=-2214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101100; // iC=-1556 
// vC = 14'b1111011011110110; // vC=-2314 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010101; // iC=-1515 
// vC = 14'b1111011100110000; // vC=-2256 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010100; // iC=-1580 
// vC = 14'b1111011010101100; // vC=-2388 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100011; // iC=-1693 
// vC = 14'b1111011011111110; // vC=-2306 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011011; // iC=-1509 
// vC = 14'b1111011001100001; // vC=-2463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001111; // iC=-1649 
// vC = 14'b1111011010111011; // vC=-2373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100001; // iC=-1503 
// vC = 14'b1111011100000100; // vC=-2300 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010100; // iC=-1708 
// vC = 14'b1111011010011000; // vC=-2408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011011; // iC=-1701 
// vC = 14'b1111011010011110; // vC=-2402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010001; // iC=-1583 
// vC = 14'b1111011010111000; // vC=-2376 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001010; // iC=-1654 
// vC = 14'b1111011010110110; // vC=-2378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101111; // iC=-1425 
// vC = 14'b1111011100010000; // vC=-2288 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010001; // iC=-1391 
// vC = 14'b1111011011100000; // vC=-2336 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011011; // iC=-1445 
// vC = 14'b1111011001100010; // vC=-2462 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101110; // iC=-1426 
// vC = 14'b1111011000100101; // vC=-2523 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011100; // iC=-1572 
// vC = 14'b1111011001101000; // vC=-2456 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001101; // iC=-1651 
// vC = 14'b1111010111111011; // vC=-2565 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011011; // iC=-1509 
// vC = 14'b1111011000111001; // vC=-2503 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110100; // iC=-1420 
// vC = 14'b1111011100000001; // vC=-2303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010000; // iC=-1648 
// vC = 14'b1111011001111110; // vC=-2434 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101001; // iC=-1559 
// vC = 14'b1111011100010111; // vC=-2281 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011110; // iC=-1378 
// vC = 14'b1111011010101001; // vC=-2391 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001011; // iC=-1397 
// vC = 14'b1111010111100011; // vC=-2589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100010; // iC=-1502 
// vC = 14'b1111011000110110; // vC=-2506 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111010; // iC=-1414 
// vC = 14'b1111010111110000; // vC=-2576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100000; // iC=-1504 
// vC = 14'b1111011010001111; // vC=-2417 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110001; // iC=-1551 
// vC = 14'b1111011011000001; // vC=-2367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111011; // iC=-1285 
// vC = 14'b1111010111101011; // vC=-2581 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100001; // iC=-1311 
// vC = 14'b1111011010010110; // vC=-2410 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100101; // iC=-1371 
// vC = 14'b1111011010101011; // vC=-2389 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010010; // iC=-1582 
// vC = 14'b1111010111101101; // vC=-2579 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111001; // iC=-1543 
// vC = 14'b1111011001010110; // vC=-2474 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111011; // iC=-1413 
// vC = 14'b1111011000011000; // vC=-2536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011010; // iC=-1254 
// vC = 14'b1111011010110110; // vC=-2378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101110; // iC=-1298 
// vC = 14'b1111011000000111; // vC=-2553 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110000; // iC=-1424 
// vC = 14'b1111010111100101; // vC=-2587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000110; // iC=-1402 
// vC = 14'b1111010110110101; // vC=-2635 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110110; // iC=-1354 
// vC = 14'b1111011000111001; // vC=-2503 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101010; // iC=-1366 
// vC = 14'b1111011010110001; // vC=-2383 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101110; // iC=-1234 
// vC = 14'b1111010111011011; // vC=-2597 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000101; // iC=-1467 
// vC = 14'b1111010111111101; // vC=-2563 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000001; // iC=-1471 
// vC = 14'b1111011000000011; // vC=-2557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110111; // iC=-1481 
// vC = 14'b1111010111010111; // vC=-2601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111000; // iC=-1224 
// vC = 14'b1111011010100010; // vC=-2398 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010100; // iC=-1388 
// vC = 14'b1111011000100011; // vC=-2525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010010; // iC=-1390 
// vC = 14'b1111011000011000; // vC=-2536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001010; // iC=-1206 
// vC = 14'b1111010101111001; // vC=-2695 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010111; // iC=-1321 
// vC = 14'b1111011010010000; // vC=-2416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011101; // iC=-1315 
// vC = 14'b1111010110110011; // vC=-2637 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110000; // iC=-1296 
// vC = 14'b1111010110111010; // vC=-2630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110011; // iC=-1357 
// vC = 14'b1111010110111111; // vC=-2625 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010101; // iC=-1387 
// vC = 14'b1111010101011110; // vC=-2722 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001001; // iC=-1335 
// vC = 14'b1111011001011110; // vC=-2466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101010; // iC=-1238 
// vC = 14'b1111010110111110; // vC=-2626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100001; // iC=-1119 
// vC = 14'b1111011001000100; // vC=-2492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111110; // iC=-1410 
// vC = 14'b1111010110111000; // vC=-2632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100110; // iC=-1114 
// vC = 14'b1111011001011101; // vC=-2467 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000100; // iC=-1084 
// vC = 14'b1111010110111111; // vC=-2625 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000100; // iC=-1212 
// vC = 14'b1111011000100000; // vC=-2528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110001; // iC=-1103 
// vC = 14'b1111010110001000; // vC=-2680 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010101; // iC=-1259 
// vC = 14'b1111010110001111; // vC=-2673 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101001; // iC=-1303 
// vC = 14'b1111010100111010; // vC=-2758 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000011; // iC=-1149 
// vC = 14'b1111010110111100; // vC=-2628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010001; // iC=-1263 
// vC = 14'b1111011000011001; // vC=-2535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010011; // iC=-1133 
// vC = 14'b1111010100110001; // vC=-2767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010101; // iC=-1195 
// vC = 14'b1111010101000100; // vC=-2748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111010; // iC=-1094 
// vC = 14'b1111010100111101; // vC=-2755 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100011; // iC=-1117 
// vC = 14'b1111010011111010; // vC=-2822 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110011; // iC=-1293 
// vC = 14'b1111010110101000; // vC=-2648 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111010; // iC=-1222 
// vC = 14'b1111010110111001; // vC=-2631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100000; // iC=-1184 
// vC = 14'b1111010011101111; // vC=-2833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011010; // iC=-1254 
// vC = 14'b1111010110010111; // vC=-2665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011100; // iC=-1060 
// vC = 14'b1111010110000010; // vC=-2686 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001101; // iC=-1075 
// vC = 14'b1111010100111001; // vC=-2759 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111010; // iC=-1030 
// vC = 14'b1111010101000111; // vC=-2745 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000101; // iC= -955 
// vC = 14'b1111010110001000; // vC=-2680 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001011; // iC=-1077 
// vC = 14'b1111010101100011; // vC=-2717 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011011; // iC=-1061 
// vC = 14'b1111010110110011; // vC=-2637 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010010; // iC=-1134 
// vC = 14'b1111010110000011; // vC=-2685 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000110; // iC=-1018 
// vC = 14'b1111010111100100; // vC=-2588 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110110; // iC=-1162 
// vC = 14'b1111010111100010; // vC=-2590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110000; // iC=-1040 
// vC = 14'b1111010011010101; // vC=-2859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001101; // iC=-1075 
// vC = 14'b1111010110010101; // vC=-2667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011001; // iC=-1127 
// vC = 14'b1111010100101000; // vC=-2776 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010101; // iC= -939 
// vC = 14'b1111010100111000; // vC=-2760 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010101; // iC= -939 
// vC = 14'b1111010101100000; // vC=-2720 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010100; // iC= -940 
// vC = 14'b1111010110110000; // vC=-2640 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101011; // iC= -917 
// vC = 14'b1111010011101111; // vC=-2833 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001111; // iC=-1137 
// vC = 14'b1111010011110011; // vC=-2829 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110011; // iC=-1165 
// vC = 14'b1111010011111100; // vC=-2820 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011001; // iC=-1127 
// vC = 14'b1111010011010110; // vC=-2858 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001010; // iC=-1014 
// vC = 14'b1111010100010011; // vC=-2797 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101110; // iC= -978 
// vC = 14'b1111010011010010; // vC=-2862 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001000; // iC=-1016 
// vC = 14'b1111010101100001; // vC=-2719 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111110; // iC=-1026 
// vC = 14'b1111010010000110; // vC=-2938 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101110; // iC= -914 
// vC = 14'b1111010011010000; // vC=-2864 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000000; // iC=-1024 
// vC = 14'b1111010011001010; // vC=-2870 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110101; // iC= -843 
// vC = 14'b1111010010110101; // vC=-2891 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100101; // iC= -795 
// vC = 14'b1111010010100010; // vC=-2910 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010001; // iC= -943 
// vC = 14'b1111010110001001; // vC=-2679 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110100; // iC= -780 
// vC = 14'b1111010110001100; // vC=-2676 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011111; // iC= -801 
// vC = 14'b1111010100010011; // vC=-2797 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100000; // iC= -928 
// vC = 14'b1111010101100000; // vC=-2720 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000010; // iC= -894 
// vC = 14'b1111010101100000; // vC=-2720 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110011; // iC= -973 
// vC = 14'b1111010100101000; // vC=-2776 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001110; // iC= -882 
// vC = 14'b1111010100001100; // vC=-2804 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011011; // iC= -933 
// vC = 14'b1111010001111110; // vC=-2946 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010001; // iC=-1007 
// vC = 14'b1111010001111011; // vC=-2949 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100001; // iC= -927 
// vC = 14'b1111010100001110; // vC=-2802 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101110; // iC= -722 
// vC = 14'b1111010100101011; // vC=-2773 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000000; // iC= -832 
// vC = 14'b1111010101111101; // vC=-2691 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b1111010001100001; // vC=-2975 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110110; // iC= -650 
// vC = 14'b1111010001111000; // vC=-2952 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111001; // iC= -775 
// vC = 14'b1111010001011100; // vC=-2980 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010100; // iC= -748 
// vC = 14'b1111010100011101; // vC=-2787 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111010; // iC= -646 
// vC = 14'b1111010011011000; // vC=-2856 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011101; // iC= -803 
// vC = 14'b1111010010000010; // vC=-2942 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111010; // iC= -710 
// vC = 14'b1111010011111011; // vC=-2821 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111101; // iC= -771 
// vC = 14'b1111010100011000; // vC=-2792 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101011; // iC= -725 
// vC = 14'b1111010011111010; // vC=-2822 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000100; // iC= -572 
// vC = 14'b1111010100101100; // vC=-2772 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111111; // iC= -577 
// vC = 14'b1111010100111011; // vC=-2757 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010110; // iC= -746 
// vC = 14'b1111010011100000; // vC=-2848 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010010; // iC= -750 
// vC = 14'b1111010010100100; // vC=-2908 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011010; // iC= -678 
// vC = 14'b1111010101011100; // vC=-2724 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010001; // iC= -687 
// vC = 14'b1111010011001100; // vC=-2868 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100011; // iC= -477 
// vC = 14'b1111010001011101; // vC=-2979 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010010; // iC= -494 
// vC = 14'b1111010100000101; // vC=-2811 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111111; // iC= -705 
// vC = 14'b1111010101000101; // vC=-2747 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101111; // iC= -465 
// vC = 14'b1111010011110001; // vC=-2831 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011111; // iC= -609 
// vC = 14'b1111010101011100; // vC=-2724 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100111; // iC= -409 
// vC = 14'b1111010010010001; // vC=-2927 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110100; // iC= -332 
// vC = 14'b1111010100111101; // vC=-2755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011110; // iC= -610 
// vC = 14'b1111010100001101; // vC=-2803 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101100; // iC= -404 
// vC = 14'b1111010010110111; // vC=-2889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101001; // iC= -279 
// vC = 14'b1111010001011011; // vC=-2981 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101010; // iC= -534 
// vC = 14'b1111010011011101; // vC=-2851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100000; // iC= -480 
// vC = 14'b1111010100100110; // vC=-2778 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001100; // iC= -500 
// vC = 14'b1111010011001000; // vC=-2872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011111111; // iC= -257 
// vC = 14'b1111010001111001; // vC=-2951 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110010; // iC= -462 
// vC = 14'b1111010000101010; // vC=-3030 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011000; // iC= -360 
// vC = 14'b1111010010111111; // vC=-2881 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000011; // iC= -317 
// vC = 14'b1111010000111001; // vC=-3015 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101101; // iC= -147 
// vC = 14'b1111010010010011; // vC=-2925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101011110; // iC= -162 
// vC = 14'b1111010001100110; // vC=-2970 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010001; // iC= -239 
// vC = 14'b1111010011010001; // vC=-2863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100100; // iC=  -92 
// vC = 14'b1111010100110100; // vC=-2764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010101; // iC= -363 
// vC = 14'b1111010001001001; // vC=-2999 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011100110; // iC= -282 
// vC = 14'b1111010011111011; // vC=-2821 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010111; // iC=  -41 
// vC = 14'b1111010001010110; // vC=-2986 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101101; // iC= -211 
// vC = 14'b1111010001101100; // vC=-2964 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100101; // iC=  -27 
// vC = 14'b1111010010110000; // vC=-2896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001100; // iC= -116 
// vC = 14'b1111010000000011; // vC=-3069 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000111; // iC=  -57 
// vC = 14'b1111010011011111; // vC=-2849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000010; // iC= -126 
// vC = 14'b1111010010011000; // vC=-2920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111100; // iC=  -68 
// vC = 14'b1111010011010011; // vC=-2861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101010; // iC=   42 
// vC = 14'b1111010100110110; // vC=-2762 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111110; // iC= -130 
// vC = 14'b1111010101001000; // vC=-2744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011010; // iC=  154 
// vC = 14'b1111010001010111; // vC=-2985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010010; // iC=   82 
// vC = 14'b1111010100000001; // vC=-2815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111111; // iC=  191 
// vC = 14'b1111010001101101; // vC=-2963 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101001; // iC=   41 
// vC = 14'b1111010000011001; // vC=-3047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011011011; // iC=  219 
// vC = 14'b1111010101001101; // vC=-2739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011101; // iC=  157 
// vC = 14'b1111010011000001; // vC=-2879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101111; // iC=  111 
// vC = 14'b1111010011000010; // vC=-2878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101110; // iC=  110 
// vC = 14'b1111010010100001; // vC=-2911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001011; // iC=  139 
// vC = 14'b1111010001110001; // vC=-2959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001001; // iC=  201 
// vC = 14'b1111010000110001; // vC=-3023 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101111; // iC=  239 
// vC = 14'b1111010000100000; // vC=-3040 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001000; // iC=  264 
// vC = 14'b1111010000101100; // vC=-3028 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110110; // iC=  182 
// vC = 14'b1111010000100110; // vC=-3034 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010110; // iC=  214 
// vC = 14'b1111010000101101; // vC=-3027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011001; // iC=  473 
// vC = 14'b1111010100100000; // vC=-2784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001100; // iC=  460 
// vC = 14'b1111010100110000; // vC=-2768 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101001; // iC=  425 
// vC = 14'b1111010010011011; // vC=-2917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010110; // iC=  534 
// vC = 14'b1111010101001110; // vC=-2738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100011; // iC=  547 
// vC = 14'b1111010010011010; // vC=-2918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110010; // iC=  562 
// vC = 14'b1111010010010010; // vC=-2926 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011010; // iC=  410 
// vC = 14'b1111010101000001; // vC=-2751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011111; // iC=  607 
// vC = 14'b1111010101101101; // vC=-2707 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101001; // iC=  617 
// vC = 14'b1111010100001001; // vC=-2807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100110; // iC=  678 
// vC = 14'b1111010011101111; // vC=-2833 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110010; // iC=  754 
// vC = 14'b1111010010111001; // vC=-2887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011110; // iC=  542 
// vC = 14'b1111010010011000; // vC=-2920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111110; // iC=  766 
// vC = 14'b1111010101011010; // vC=-2726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111100; // iC=  700 
// vC = 14'b1111010010101001; // vC=-2903 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110100; // iC=  628 
// vC = 14'b1111010101111010; // vC=-2694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011100; // iC=  732 
// vC = 14'b1111010010000111; // vC=-2937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011001; // iC=  793 
// vC = 14'b1111010101110100; // vC=-2700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010001; // iC=  785 
// vC = 14'b1111010110010100; // vC=-2668 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111100; // iC=  892 
// vC = 14'b1111010101010011; // vC=-2733 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111100; // iC=  764 
// vC = 14'b1111010100011111; // vC=-2785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100001; // iC=  993 
// vC = 14'b1111010010101111; // vC=-2897 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010000; // iC=  976 
// vC = 14'b1111010110011100; // vC=-2660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001000; // iC=  776 
// vC = 14'b1111010101100000; // vC=-2720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000010; // iC= 1026 
// vC = 14'b1111010010111011; // vC=-2885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110111; // iC= 1079 
// vC = 14'b1111010101001101; // vC=-2739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100011; // iC=  995 
// vC = 14'b1111010010100001; // vC=-2911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110000; // iC= 1136 
// vC = 14'b1111010110001000; // vC=-2680 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010001; // iC=  977 
// vC = 14'b1111010110100011; // vC=-2653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000111; // iC= 1223 
// vC = 14'b1111010111000111; // vC=-2617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110000; // iC= 1136 
// vC = 14'b1111010110101000; // vC=-2648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101001; // iC= 1065 
// vC = 14'b1111010011100111; // vC=-2841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010111; // iC=  983 
// vC = 14'b1111010011100100; // vC=-2844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001101; // iC= 1293 
// vC = 14'b1111010110110100; // vC=-2636 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111010; // iC= 1338 
// vC = 14'b1111010111000011; // vC=-2621 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110010; // iC= 1138 
// vC = 14'b1111010101110001; // vC=-2703 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111101; // iC= 1341 
// vC = 14'b1111010101000001; // vC=-2751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100110; // iC= 1254 
// vC = 14'b1111010011011001; // vC=-2855 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111110; // iC= 1214 
// vC = 14'b1111010110101110; // vC=-2642 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101111; // iC= 1199 
// vC = 14'b1111010111111111; // vC=-2561 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110000; // iC= 1200 
// vC = 14'b1111010110000100; // vC=-2684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000001; // iC= 1473 
// vC = 14'b1111010011001000; // vC=-2872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000000; // iC= 1472 
// vC = 14'b1111010011010110; // vC=-2858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011100; // iC= 1372 
// vC = 14'b1111010110010100; // vC=-2668 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110110; // iC= 1398 
// vC = 14'b1111010100001100; // vC=-2804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101001; // iC= 1321 
// vC = 14'b1111010100110011; // vC=-2765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011111; // iC= 1567 
// vC = 14'b1111011000001110; // vC=-2546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000010; // iC= 1346 
// vC = 14'b1111010101111101; // vC=-2691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010100; // iC= 1364 
// vC = 14'b1111010100111101; // vC=-2755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010101; // iC= 1557 
// vC = 14'b1111010110011000; // vC=-2664 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000110; // iC= 1414 
// vC = 14'b1111010100011110; // vC=-2786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011101; // iC= 1501 
// vC = 14'b1111010101010000; // vC=-2736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000000; // iC= 1408 
// vC = 14'b1111010111001101; // vC=-2611 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001111; // iC= 1679 
// vC = 14'b1111010111100011; // vC=-2589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000111; // iC= 1415 
// vC = 14'b1111010101001100; // vC=-2740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110111; // iC= 1655 
// vC = 14'b1111010111100101; // vC=-2587 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011001; // iC= 1625 
// vC = 14'b1111010101111001; // vC=-2695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010000; // iC= 1744 
// vC = 14'b1111011000101011; // vC=-2517 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001000; // iC= 1672 
// vC = 14'b1111011001110011; // vC=-2445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111001; // iC= 1721 
// vC = 14'b1111010111000110; // vC=-2618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111010; // iC= 1530 
// vC = 14'b1111010110101100; // vC=-2644 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000110; // iC= 1798 
// vC = 14'b1111010110011011; // vC=-2661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111011; // iC= 1595 
// vC = 14'b1111011000011100; // vC=-2532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100001; // iC= 1569 
// vC = 14'b1111011000101010; // vC=-2518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b1111010101101011; // vC=-2709 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110100; // iC= 1716 
// vC = 14'b1111011001000011; // vC=-2493 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111000; // iC= 1720 
// vC = 14'b1111011001011101; // vC=-2467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000100; // iC= 1732 
// vC = 14'b1111010111100111; // vC=-2585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101111; // iC= 1647 
// vC = 14'b1111010111101111; // vC=-2577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000001; // iC= 1857 
// vC = 14'b1111011000100111; // vC=-2521 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000110; // iC= 1798 
// vC = 14'b1111011000001001; // vC=-2551 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101111; // iC= 1711 
// vC = 14'b1111010111000001; // vC=-2623 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b1111010110111001; // vC=-2631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b1111011011011101; // vC=-2339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010110; // iC= 1814 
// vC = 14'b1111011001010001; // vC=-2479 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b1111011011011010; // vC=-2342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110001; // iC= 2033 
// vC = 14'b1111011100010001; // vC=-2287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b1111011001000001; // vC=-2495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b1111011001110011; // vC=-2445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011110; // iC= 2078 
// vC = 14'b1111011010000010; // vC=-2430 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b1111011000111111; // vC=-2497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100010; // iC= 2018 
// vC = 14'b1111011011001101; // vC=-2355 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111011001001000; // vC=-2488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110100; // iC= 2100 
// vC = 14'b1111011100111011; // vC=-2245 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010100; // iC= 2068 
// vC = 14'b1111011010011000; // vC=-2408 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111101; // iC= 2045 
// vC = 14'b1111011101100010; // vC=-2206 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b1111011001100011; // vC=-2461 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100000; // iC= 2080 
// vC = 14'b1111011001001001; // vC=-2487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b1111011001100010; // vC=-2462 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010000; // iC= 2064 
// vC = 14'b1111011101011100; // vC=-2212 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101010; // iC= 1898 
// vC = 14'b1111011101110100; // vC=-2188 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111111; // iC= 2111 
// vC = 14'b1111011100110111; // vC=-2249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b1111011010000100; // vC=-2428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101111; // iC= 2159 
// vC = 14'b1111011011101011; // vC=-2325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000001; // iC= 2241 
// vC = 14'b1111011110010101; // vC=-2155 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100101; // iC= 2149 
// vC = 14'b1111011001111110; // vC=-2434 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001010; // iC= 2250 
// vC = 14'b1111011010001101; // vC=-2419 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011100010; // iC= 2274 
// vC = 14'b1111011110000010; // vC=-2174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111111; // iC= 2239 
// vC = 14'b1111011110111011; // vC=-2117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000000; // iC= 2112 
// vC = 14'b1111011101110111; // vC=-2185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000001; // iC= 2177 
// vC = 14'b1111011100011110; // vC=-2274 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111011101100111; // vC=-2201 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b1111011111001100; // vC=-2100 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111011111101111; // vC=-2065 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b1111011110001100; // vC=-2164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011110010; // iC= 2290 
// vC = 14'b1111011101011111; // vC=-2209 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111011011110111; // vC=-2313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001000; // iC= 2248 
// vC = 14'b1111011101000101; // vC=-2235 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010011; // iC= 2259 
// vC = 14'b1111011011111110; // vC=-2306 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100100110; // iC= 2342 
// vC = 14'b1111011100111000; // vC=-2248 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010000; // iC= 2256 
// vC = 14'b1111100000100001; // vC=-2015 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000111; // iC= 2055 
// vC = 14'b1111011101010010; // vC=-2222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110110; // iC= 2166 
// vC = 14'b1111100001001010; // vC=-1974 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100001100; // iC= 2316 
// vC = 14'b1111011110001011; // vC=-2165 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000100; // iC= 2180 
// vC = 14'b1111100001011001; // vC=-1959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111000; // iC= 2104 
// vC = 14'b1111011110101000; // vC=-2136 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100101101; // iC= 2349 
// vC = 14'b1111011101101001; // vC=-2199 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011110111; // iC= 2295 
// vC = 14'b1111100001001100; // vC=-1972 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010000; // iC= 2256 
// vC = 14'b1111011110111011; // vC=-2117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b1111100001010000; // vC=-1968 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010011; // iC= 2131 
// vC = 14'b1111100010011011; // vC=-1893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010011; // iC= 2259 
// vC = 14'b1111011111000000; // vC=-2112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000111; // iC= 2247 
// vC = 14'b1111011110111011; // vC=-2117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101001101; // iC= 2381 
// vC = 14'b1111100000100010; // vC=-2014 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111101; // iC= 2109 
// vC = 14'b1111011110011011; // vC=-2149 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011110010; // iC= 2290 
// vC = 14'b1111100001000101; // vC=-1979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011011; // iC= 2075 
// vC = 14'b1111100011000001; // vC=-1855 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000011; // iC= 2243 
// vC = 14'b1111100010111111; // vC=-1857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001100; // iC= 2188 
// vC = 14'b1111100010010011; // vC=-1901 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011110; // iC= 2142 
// vC = 14'b1111100000100111; // vC=-2009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101000101; // iC= 2373 
// vC = 14'b1111100010110010; // vC=-1870 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101000111; // iC= 2375 
// vC = 14'b1111100010011011; // vC=-1893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101111; // iC= 2159 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110110; // iC= 2166 
// vC = 14'b1111100001000001; // vC=-1983 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b1111100001111100; // vC=-1924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101100; // iC= 2220 
// vC = 14'b1111100000111011; // vC=-1989 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111100000111111; // vC=-1985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101101001; // iC= 2409 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111110; // iC= 2174 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101001011; // iC= 2379 
// vC = 14'b1111100101001100; // vC=-1716 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101101; // iC= 2093 
// vC = 14'b1111100001011000; // vC=-1960 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001000; // iC= 2248 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001101; // iC= 2253 
// vC = 14'b1111100101010100; // vC=-1708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001100; // iC= 2188 
// vC = 14'b1111100101111001; // vC=-1671 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100110011; // iC= 2355 
// vC = 14'b1111100110100011; // vC=-1629 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111100110001100; // vC=-1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010001; // iC= 2257 
// vC = 14'b1111100010001011; // vC=-1909 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011100101; // iC= 2277 
// vC = 14'b1111100101111010; // vC=-1670 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011001; // iC= 2201 
// vC = 14'b1111100011000000; // vC=-1856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b1111100011011000; // vC=-1832 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101010000; // iC= 2384 
// vC = 14'b1111100110101100; // vC=-1620 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000011; // iC= 2179 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001001; // iC= 2185 
// vC = 14'b1111100101000111; // vC=-1721 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011011110; // iC= 2270 
// vC = 14'b1111100011101010; // vC=-1814 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010101; // iC= 2133 
// vC = 14'b1111100100010100; // vC=-1772 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000101; // iC= 2181 
// vC = 14'b1111100111111011; // vC=-1541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011101; // iC= 2141 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110100; // iC= 2228 
// vC = 14'b1111100101101100; // vC=-1684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010000; // iC= 2192 
// vC = 14'b1111100100011111; // vC=-1761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100010001; // iC= 2321 
// vC = 14'b1111101000111000; // vC=-1480 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001011; // iC= 2187 
// vC = 14'b1111100100101000; // vC=-1752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100101011; // iC= 2347 
// vC = 14'b1111101000110011; // vC=-1485 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100100110; // iC= 2342 
// vC = 14'b1111100101010010; // vC=-1710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110011; // iC= 2163 
// vC = 14'b1111100110001111; // vC=-1649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110011; // iC= 2227 
// vC = 14'b1111101001010111; // vC=-1449 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101000; // iC= 2152 
// vC = 14'b1111100111100111; // vC=-1561 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100010; // iC= 2146 
// vC = 14'b1111101001001111; // vC=-1457 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100000100; // iC= 2308 
// vC = 14'b1111100111001100; // vC=-1588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011101010; // iC= 2282 
// vC = 14'b1111101001011011; // vC=-1445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100011001; // iC= 2329 
// vC = 14'b1111101001111011; // vC=-1413 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101011001; // iC= 2393 
// vC = 14'b1111101001011001; // vC=-1447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100110111; // iC= 2359 
// vC = 14'b1111100111000000; // vC=-1600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100000010; // iC= 2306 
// vC = 14'b1111101010110000; // vC=-1360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100101101; // iC= 2349 
// vC = 14'b1111101000101100; // vC=-1492 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101000111; // iC= 2375 
// vC = 14'b1111100111011000; // vC=-1576 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100010011; // iC= 2323 
// vC = 14'b1111100111011011; // vC=-1573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111011; // iC= 2235 
// vC = 14'b1111101011001110; // vC=-1330 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010010; // iC= 2194 
// vC = 14'b1111101001100010; // vC=-1438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101001; // iC= 2153 
// vC = 14'b1111101000010100; // vC=-1516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011100001; // iC= 2273 
// vC = 14'b1111101010100101; // vC=-1371 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100110001001; // iC= 2441 
// vC = 14'b1111101001010001; // vC=-1455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011101001; // iC= 2281 
// vC = 14'b1111101011001101; // vC=-1331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011101001; // iC= 2281 
// vC = 14'b1111101011011101; // vC=-1315 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001111; // iC= 2255 
// vC = 14'b1111101000010100; // vC=-1516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b1111101001010100; // vC=-1452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100110000001; // iC= 2433 
// vC = 14'b1111101000100010; // vC=-1502 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110001; // iC= 2161 
// vC = 14'b1111101010110100; // vC=-1356 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100100110; // iC= 2342 
// vC = 14'b1111101100100011; // vC=-1245 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100100; // iC= 2212 
// vC = 14'b1111101011010000; // vC=-1328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100110001001; // iC= 2441 
// vC = 14'b1111101100000001; // vC=-1279 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b1111101100000101; // vC=-1275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101000000; // iC= 2368 
// vC = 14'b1111101010111100; // vC=-1348 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101000000; // iC= 2368 
// vC = 14'b1111101001000100; // vC=-1468 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011011000; // iC= 2264 
// vC = 14'b1111101100110001; // vC=-1231 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100001; // iC= 2145 
// vC = 14'b1111101110000100; // vC=-1148 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100110100; // iC= 2356 
// vC = 14'b1111101011001101; // vC=-1331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011110001; // iC= 2289 
// vC = 14'b1111101010010101; // vC=-1387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101011100; // iC= 2396 
// vC = 14'b1111101011010111; // vC=-1321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101111101; // iC= 2429 
// vC = 14'b1111101100110010; // vC=-1230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011011; // iC= 2139 
// vC = 14'b1111101110011001; // vC=-1127 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101110000; // iC= 2416 
// vC = 14'b1111101110001101; // vC=-1139 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100001001; // iC= 2313 
// vC = 14'b1111101010100101; // vC=-1371 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100001000; // iC= 2312 
// vC = 14'b1111101011001100; // vC=-1332 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101000111; // iC= 2375 
// vC = 14'b1111101110000000; // vC=-1152 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100110001001; // iC= 2441 
// vC = 14'b1111101111110011; // vC=-1037 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011111011; // iC= 2299 
// vC = 14'b1111101100100010; // vC=-1246 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011000; // iC= 2200 
// vC = 14'b1111101011111011; // vC=-1285 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011011; // iC= 2139 
// vC = 14'b1111101101100110; // vC=-1178 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100110010; // iC= 2354 
// vC = 14'b1111101111000011; // vC=-1085 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100100; // iC= 2148 
// vC = 14'b1111101011111110; // vC=-1282 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101000111; // iC= 2375 
// vC = 14'b1111101101000101; // vC=-1211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001010; // iC= 2250 
// vC = 14'b1111101111100011; // vC=-1053 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101111101; // iC= 2429 
// vC = 14'b1111110000001001; // vC=-1015 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100101101; // iC= 2349 
// vC = 14'b1111110001010000; // vC= -944 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001110; // iC= 2254 
// vC = 14'b1111110001010111; // vC= -937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011011100; // iC= 2268 
// vC = 14'b1111101100110000; // vC=-1232 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101011100; // iC= 2396 
// vC = 14'b1111101111011000; // vC=-1064 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110000; // iC= 2224 
// vC = 14'b1111101101111101; // vC=-1155 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100011111; // iC= 2335 
// vC = 14'b1111101101011001; // vC=-1191 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000010; // iC= 2114 
// vC = 14'b1111110001110110; // vC= -906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111111; // iC= 2239 
// vC = 14'b1111110000111010; // vC= -966 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101110; // iC= 2158 
// vC = 14'b1111101111100011; // vC=-1053 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101001; // iC= 2153 
// vC = 14'b1111110000010001; // vC=-1007 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011110100; // iC= 2292 
// vC = 14'b1111110000011001; // vC= -999 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010000; // iC= 2192 
// vC = 14'b1111101110000101; // vC=-1147 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100110011; // iC= 2355 
// vC = 14'b1111101111101110; // vC=-1042 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011011011; // iC= 2267 
// vC = 14'b1111101111100000; // vC=-1056 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111101; // iC= 2109 
// vC = 14'b1111110000001001; // vC=-1015 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101101110; // iC= 2414 
// vC = 14'b1111110010110011; // vC= -845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100110000000; // iC= 2432 
// vC = 14'b1111110010011111; // vC= -865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001101; // iC= 2253 
// vC = 14'b1111110000100101; // vC= -987 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000101; // iC= 2181 
// vC = 14'b1111110001101010; // vC= -918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011011010; // iC= 2266 
// vC = 14'b1111110011011000; // vC= -808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011111110; // iC= 2302 
// vC = 14'b1111110010100111; // vC= -857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100010100; // iC= 2324 
// vC = 14'b1111110100101011; // vC= -725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100110; // iC= 2214 
// vC = 14'b1111110000011101; // vC= -995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011111; // iC= 2143 
// vC = 14'b1111110000000111; // vC=-1017 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011110110; // iC= 2294 
// vC = 14'b1111110100100010; // vC= -734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100010000; // iC= 2320 
// vC = 14'b1111110100101001; // vC= -727 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101101100; // iC= 2412 
// vC = 14'b1111110100000011; // vC= -765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101101011; // iC= 2411 
// vC = 14'b1111110100001100; // vC= -756 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011111110; // iC= 2302 
// vC = 14'b1111110100011110; // vC= -738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111010; // iC= 2234 
// vC = 14'b1111110100011000; // vC= -744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001101; // iC= 2253 
// vC = 14'b1111110100100111; // vC= -729 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101000101; // iC= 2373 
// vC = 14'b1111110100001011; // vC= -757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111011; // iC= 2171 
// vC = 14'b1111110100111000; // vC= -712 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011111000; // iC= 2296 
// vC = 14'b1111110001111100; // vC= -900 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b1111110101110011; // vC= -653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100110000; // iC= 2352 
// vC = 14'b1111110110000101; // vC= -635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011111011; // iC= 2299 
// vC = 14'b1111110101000110; // vC= -698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101000111; // iC= 2375 
// vC = 14'b1111110101100100; // vC= -668 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100011101; // iC= 2333 
// vC = 14'b1111110010111100; // vC= -836 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010011; // iC= 2259 
// vC = 14'b1111110101001001; // vC= -695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100111100; // iC= 2364 
// vC = 14'b1111110100000010; // vC= -766 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011100111; // iC= 2279 
// vC = 14'b1111110110011110; // vC= -610 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b1111110100101010; // vC= -726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100000001; // iC= 2305 
// vC = 14'b1111111000000100; // vC= -508 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011100011; // iC= 2275 
// vC = 14'b1111110111001111; // vC= -561 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111010; // iC= 2234 
// vC = 14'b1111110111100010; // vC= -542 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b1111111000001010; // vC= -502 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101001; // iC= 2217 
// vC = 14'b1111110110000011; // vC= -637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111110100100110; // vC= -730 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110110; // iC= 2102 
// vC = 14'b1111110100001101; // vC= -755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001111; // iC= 2191 
// vC = 14'b1111111000010011; // vC= -493 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100000001; // iC= 2305 
// vC = 14'b1111110101111110; // vC= -642 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100110110; // iC= 2358 
// vC = 14'b1111110100011011; // vC= -741 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100111000; // iC= 2360 
// vC = 14'b1111110101100011; // vC= -669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101011; // iC= 2219 
// vC = 14'b1111110101111001; // vC= -647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111001; // iC= 2169 
// vC = 14'b1111110111111010; // vC= -518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100001; // iC= 2145 
// vC = 14'b1111111001100110; // vC= -410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100101000011; // iC= 2371 
// vC = 14'b1111110111011100; // vC= -548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011010; // iC= 2074 
// vC = 14'b1111111000010101; // vC= -491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011101010; // iC= 2282 
// vC = 14'b1111111010100011; // vC= -349 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100010010; // iC= 2322 
// vC = 14'b1111111001110101; // vC= -395 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100111; // iC= 2151 
// vC = 14'b1111110111100000; // vC= -544 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000011; // iC= 2179 
// vC = 14'b1111111001111110; // vC= -386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011100111; // iC= 2279 
// vC = 14'b1111110110001111; // vC= -625 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011000; // iC= 2200 
// vC = 14'b1111111010001000; // vC= -376 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000010; // iC= 2050 
// vC = 14'b1111111010011010; // vC= -358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111110111001111; // vC= -561 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110100; // iC= 2228 
// vC = 14'b1111111011011000; // vC= -296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100000010; // iC= 2306 
// vC = 14'b1111111001001011; // vC= -437 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110110; // iC= 2102 
// vC = 14'b1111110111111111; // vC= -513 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101010; // iC= 2090 
// vC = 14'b1111111001100111; // vC= -409 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000111; // iC= 2183 
// vC = 14'b1111111000001000; // vC= -504 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101101; // iC= 2029 
// vC = 14'b1111110111101100; // vC= -532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110011; // iC= 2227 
// vC = 14'b1111111010101100; // vC= -340 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100001; // iC= 2017 
// vC = 14'b1111111011011001; // vC= -295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000100; // iC= 2244 
// vC = 14'b1111111100011010; // vC= -230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100100000010; // iC= 2306 
// vC = 14'b1111111100010010; // vC= -238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000001; // iC= 2049 
// vC = 14'b1111111000100101; // vC= -475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011111; // iC= 2015 
// vC = 14'b1111111100111101; // vC= -195 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101111; // iC= 2095 
// vC = 14'b1111111011000110; // vC= -314 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101001; // iC= 2217 
// vC = 14'b1111111010010100; // vC= -364 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111110; // iC= 2238 
// vC = 14'b1111111000111001; // vC= -455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010010; // iC= 2130 
// vC = 14'b1111111101011011; // vC= -165 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011111110; // iC= 2302 
// vC = 14'b1111111101111110; // vC= -130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011011010; // iC= 2266 
// vC = 14'b1111111101001000; // vC= -184 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100000; // iC= 2080 
// vC = 14'b1111111010010100; // vC= -364 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000001; // iC= 2177 
// vC = 14'b1111111010111001; // vC= -327 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b1111111010001100; // vC= -372 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010110; // iC= 2198 
// vC = 14'b1111111001110000; // vC= -400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100111; // iC= 2215 
// vC = 14'b1111111001111010; // vC= -390 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100111; // iC= 2151 
// vC = 14'b1111111011001011; // vC= -309 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100011; // iC= 2147 
// vC = 14'b1111111111001011; // vC=  -53 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011011; // iC= 2203 
// vC = 14'b1111111100101101; // vC= -211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101100; // iC= 2092 
// vC = 14'b1111111110010001; // vC= -111 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010110; // iC= 2070 
// vC = 14'b1111111111011000; // vC=  -40 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b1111111110010100; // vC= -108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010001; // iC= 2129 
// vC = 14'b1111111100101111; // vC= -209 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b1111111011001110; // vC= -306 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110010; // iC= 2034 
// vC = 14'b1111111101110000; // vC= -144 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111011; // iC= 2107 
// vC = 14'b1111111111001111; // vC=  -49 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001000; // iC= 1992 
// vC = 14'b1111111110111000; // vC=  -72 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101100; // iC= 2220 
// vC = 14'b1111111110001100; // vC= -116 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110001; // iC= 1969 
// vC = 14'b1111111101000011; // vC= -189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b1111111101001111; // vC= -177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101000; // iC= 2216 
// vC = 14'b1111111111011111; // vC=  -33 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001101; // iC= 1997 
// vC = 14'b1111111111100111; // vC=  -25 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111100; // iC= 1980 
// vC = 14'b1111111101010010; // vC= -174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001010; // iC= 2250 
// vC = 14'b0000000000101101; // vC=   45 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011100; // iC= 2204 
// vC = 14'b0000000001101100; // vC=  108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101100; // iC= 2220 
// vC = 14'b1111111110001101; // vC= -115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111010; // iC= 2234 
// vC = 14'b0000000000011111; // vC=   31 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b1111111110010001; // vC= -111 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b1111111111001101; // vC=  -51 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000010; // iC= 1986 
// vC = 14'b1111111111011110; // vC=  -34 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b0000000010000100; // vC=  132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b1111111111010110; // vC=  -42 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101010; // iC= 2090 
// vC = 14'b1111111111001000; // vC=  -56 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100101; // iC= 2149 
// vC = 14'b0000000010000011; // vC=  131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000011; // iC= 2179 
// vC = 14'b1111111111100001; // vC=  -31 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101010; // iC= 2154 
// vC = 14'b0000000001100101; // vC=  101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b0000000000000101; // vC=    5 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010100; // iC= 2068 
// vC = 14'b1111111110100101; // vC=  -91 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111111111010001; // vC=  -47 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111111111100101; // vC=  -27 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010001; // iC= 1937 
// vC = 14'b0000000010000110; // vC=  134 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100101; // iC= 2149 
// vC = 14'b1111111111010000; // vC=  -48 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b0000000011111000; // vC=  248 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001110; // iC= 2126 
// vC = 14'b0000000000101100; // vC=   44 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b0000000100010111; // vC=  279 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001001; // iC= 2057 
// vC = 14'b0000000001101000; // vC=  104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b0000000001000100; // vC=   68 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b0000000100110000; // vC=  304 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010001; // iC= 2065 
// vC = 14'b0000000011000010; // vC=  194 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b0000000001111011; // vC=  123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b0000000001111001; // vC=  121 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b0000000011011110; // vC=  222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001010; // iC= 1994 
// vC = 14'b0000000000100110; // vC=   38 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001100; // iC= 1868 
// vC = 14'b0000000010011001; // vC=  153 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b0000000011000110; // vC=  198 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b0000000011011010; // vC=  218 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011100; // iC= 2076 
// vC = 14'b0000000001111111; // vC=  127 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b0000000010010100; // vC=  148 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011010; // iC= 1818 
// vC = 14'b0000000001100011; // vC=   99 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b0000000011110100; // vC=  244 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b0000000001100110; // vC=  102 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110010; // iC= 2034 
// vC = 14'b0000000101100100; // vC=  356 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100111; // iC= 1895 
// vC = 14'b0000000011101101; // vC=  237 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101010; // iC= 1834 
// vC = 14'b0000000110000011; // vC=  387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b0000000011101001; // vC=  233 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110110; // iC= 1974 
// vC = 14'b0000000100110001; // vC=  305 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000110; // iC= 1862 
// vC = 14'b0000000110101000; // vC=  424 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000110; // iC= 1862 
// vC = 14'b0000000011110110; // vC=  246 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100000; // iC= 1888 
// vC = 14'b0000000010101110; // vC=  174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101001; // iC= 1769 
// vC = 14'b0000000011100110; // vC=  230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b0000000101010110; // vC=  342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b0000000110101010; // vC=  426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101100; // iC= 1772 
// vC = 14'b0000000110101100; // vC=  428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b0000000110001110; // vC=  398 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111100; // iC= 1916 
// vC = 14'b0000000110000100; // vC=  388 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010101; // iC= 1877 
// vC = 14'b0000000101010110; // vC=  342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011010; // iC= 1754 
// vC = 14'b0000000110011100; // vC=  412 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b0000000100011000; // vC=  280 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100110; // iC= 1830 
// vC = 14'b0000001000110000; // vC=  560 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001110; // iC= 1742 
// vC = 14'b0000000111111101; // vC=  509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000010; // iC= 1794 
// vC = 14'b0000000101001100; // vC=  332 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000100; // iC= 1860 
// vC = 14'b0000000110011100; // vC=  412 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000100; // iC= 1924 
// vC = 14'b0000001000011011; // vC=  539 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b0000000110010100; // vC=  404 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111000; // iC= 1848 
// vC = 14'b0000001001000001; // vC=  577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111110; // iC= 1918 
// vC = 14'b0000001001101010; // vC=  618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011000; // iC= 1752 
// vC = 14'b0000000101100000; // vC=  352 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101010; // iC= 1898 
// vC = 14'b0000000110001010; // vC=  394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b0000000101001001; // vC=  329 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010111; // iC= 1687 
// vC = 14'b0000001010001010; // vC=  650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100000; // iC= 1760 
// vC = 14'b0000001001101000; // vC=  616 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000010; // iC= 1986 
// vC = 14'b0000001000000110; // vC=  518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b0000001000100001; // vC=  545 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101111; // iC= 1711 
// vC = 14'b0000000110111001; // vC=  441 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101001; // iC= 1769 
// vC = 14'b0000000111010011; // vC=  467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b0000000110000010; // vC=  386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110110; // iC= 1718 
// vC = 14'b0000000110000111; // vC=  391 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001110; // iC= 1742 
// vC = 14'b0000001001011011; // vC=  603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000010; // iC= 1794 
// vC = 14'b0000000111001111; // vC=  463 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000000; // iC= 1792 
// vC = 14'b0000000111101101; // vC=  493 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000110; // iC= 1862 
// vC = 14'b0000000111100111; // vC=  487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100001; // iC= 1633 
// vC = 14'b0000001011011101; // vC=  733 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100100; // iC= 1828 
// vC = 14'b0000000111000100; // vC=  452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111001; // iC= 1785 
// vC = 14'b0000000111101010; // vC=  490 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110011; // iC= 1779 
// vC = 14'b0000001010011001; // vC=  665 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100100; // iC= 1700 
// vC = 14'b0000000111010101; // vC=  469 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b0000001011010000; // vC=  720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010000; // iC= 1616 
// vC = 14'b0000001000000100; // vC=  516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111101; // iC= 1597 
// vC = 14'b0000001000001110; // vC=  526 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b0000001001001111; // vC=  591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100100; // iC= 1636 
// vC = 14'b0000001000101000; // vC=  552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000010; // iC= 1794 
// vC = 14'b0000001001100101; // vC=  613 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101110; // iC= 1710 
// vC = 14'b0000001001101011; // vC=  619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101100; // iC= 1580 
// vC = 14'b0000001100111111; // vC=  831 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001101; // iC= 1677 
// vC = 14'b0000001100001101; // vC=  781 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011110; // iC= 1822 
// vC = 14'b0000001001111010; // vC=  634 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000100; // iC= 1732 
// vC = 14'b0000001100110000; // vC=  816 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b0000001001100011; // vC=  611 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001010; // iC= 1802 
// vC = 14'b0000001100001001; // vC=  777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111011; // iC= 1723 
// vC = 14'b0000001010001100; // vC=  652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000111; // iC= 1799 
// vC = 14'b0000001101001011; // vC=  843 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110000; // iC= 1648 
// vC = 14'b0000001010100011; // vC=  675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000100; // iC= 1540 
// vC = 14'b0000001010111001; // vC=  697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101100; // iC= 1772 
// vC = 14'b0000001110001100; // vC=  908 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b0000001100000000; // vC=  768 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111010; // iC= 1530 
// vC = 14'b0000001001110011; // vC=  627 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101100; // iC= 1772 
// vC = 14'b0000001110010010; // vC=  914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011111; // iC= 1695 
// vC = 14'b0000001101101001; // vC=  873 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100100; // iC= 1700 
// vC = 14'b0000001010101001; // vC=  681 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101011; // iC= 1515 
// vC = 14'b0000001010011010; // vC=  666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001111; // iC= 1615 
// vC = 14'b0000001100000110; // vC=  774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101100; // iC= 1516 
// vC = 14'b0000001101001010; // vC=  842 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011001; // iC= 1625 
// vC = 14'b0000001111001011; // vC=  971 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001100; // iC= 1676 
// vC = 14'b0000001011001111; // vC=  719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001000; // iC= 1480 
// vC = 14'b0000001110001110; // vC=  910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111001; // iC= 1657 
// vC = 14'b0000001111000011; // vC=  963 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001101; // iC= 1549 
// vC = 14'b0000001101110101; // vC=  885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100011; // iC= 1507 
// vC = 14'b0000001100110101; // vC=  821 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011000; // iC= 1560 
// vC = 14'b0000001111010011; // vC=  979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111101; // iC= 1725 
// vC = 14'b0000001110011101; // vC=  925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101101; // iC= 1709 
// vC = 14'b0000001100111111; // vC=  831 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100110; // iC= 1638 
// vC = 14'b0000001100000100; // vC=  772 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100101; // iC= 1701 
// vC = 14'b0000001100001001; // vC=  777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011000; // iC= 1688 
// vC = 14'b0000001011111110; // vC=  766 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111110; // iC= 1662 
// vC = 14'b0000001110111001; // vC=  953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001011; // iC= 1611 
// vC = 14'b0000001110100101; // vC=  933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001111; // iC= 1487 
// vC = 14'b0000001100010111; // vC=  791 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010010; // iC= 1682 
// vC = 14'b0000001100100000; // vC=  800 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011010; // iC= 1498 
// vC = 14'b0000010000110000; // vC= 1072 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110111; // iC= 1655 
// vC = 14'b0000010000100100; // vC= 1060 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011101; // iC= 1565 
// vC = 14'b0000001110011110; // vC=  926 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101100; // iC= 1580 
// vC = 14'b0000001101001101; // vC=  845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101001; // iC= 1513 
// vC = 14'b0000001101100101; // vC=  869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010100; // iC= 1684 
// vC = 14'b0000001111000011; // vC=  963 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000110; // iC= 1670 
// vC = 14'b0000010000000000; // vC= 1024 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110111; // iC= 1527 
// vC = 14'b0000001101010101; // vC=  853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000111; // iC= 1543 
// vC = 14'b0000001101111100; // vC=  892 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110101; // iC= 1397 
// vC = 14'b0000001111000110; // vC=  966 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110101; // iC= 1589 
// vC = 14'b0000001111011100; // vC=  988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101100; // iC= 1644 
// vC = 14'b0000001101010000; // vC=  848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101101; // iC= 1453 
// vC = 14'b0000001101110111; // vC=  887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100001; // iC= 1633 
// vC = 14'b0000001111111000; // vC= 1016 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000111; // iC= 1415 
// vC = 14'b0000001101011011; // vC=  859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111000; // iC= 1464 
// vC = 14'b0000001110010011; // vC=  915 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011010; // iC= 1498 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111111; // iC= 1535 
// vC = 14'b0000001110100010; // vC=  930 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010011; // iC= 1363 
// vC = 14'b0000001110001001; // vC=  905 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101100; // iC= 1388 
// vC = 14'b0000010001010000; // vC= 1104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010101; // iC= 1557 
// vC = 14'b0000010000111011; // vC= 1083 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010100; // iC= 1300 
// vC = 14'b0000010000000000; // vC= 1024 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001100; // iC= 1484 
// vC = 14'b0000001110111000; // vC=  952 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100111; // iC= 1383 
// vC = 14'b0000010000010111; // vC= 1047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011010; // iC= 1562 
// vC = 14'b0000001110100100; // vC=  932 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101011; // iC= 1579 
// vC = 14'b0000001111111001; // vC= 1017 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100100; // iC= 1444 
// vC = 14'b0000010001011010; // vC= 1114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011100; // iC= 1308 
// vC = 14'b0000010001000011; // vC= 1091 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101100; // iC= 1452 
// vC = 14'b0000001110111001; // vC=  953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101000; // iC= 1448 
// vC = 14'b0000001111010000; // vC=  976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100100; // iC= 1508 
// vC = 14'b0000010011110100; // vC= 1268 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001100; // iC= 1548 
// vC = 14'b0000010011011010; // vC= 1242 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100110; // iC= 1254 
// vC = 14'b0000010000100010; // vC= 1058 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000101; // iC= 1221 
// vC = 14'b0000010100000001; // vC= 1281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011110; // iC= 1502 
// vC = 14'b0000010011110000; // vC= 1264 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100110; // iC= 1510 
// vC = 14'b0000010001101001; // vC= 1129 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011010; // iC= 1434 
// vC = 14'b0000010000010001; // vC= 1041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011011; // iC= 1371 
// vC = 14'b0000010000011001; // vC= 1049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110000; // iC= 1456 
// vC = 14'b0000010000010010; // vC= 1042 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110101; // iC= 1397 
// vC = 14'b0000010100000000; // vC= 1280 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110011; // iC= 1203 
// vC = 14'b0000010000101010; // vC= 1066 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011111; // iC= 1247 
// vC = 14'b0000010011010011; // vC= 1235 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011010; // iC= 1434 
// vC = 14'b0000010000001001; // vC= 1033 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000111; // iC= 1159 
// vC = 14'b0000010000011111; // vC= 1055 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111111; // iC= 1343 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010100; // iC= 1428 
// vC = 14'b0000010000101011; // vC= 1067 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011111; // iC= 1311 
// vC = 14'b0000010000110110; // vC= 1078 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000100; // iC= 1284 
// vC = 14'b0000010011110110; // vC= 1270 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010001; // iC= 1169 
// vC = 14'b0000010001001000; // vC= 1096 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001001; // iC= 1225 
// vC = 14'b0000010001111011; // vC= 1147 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011000; // iC= 1368 
// vC = 14'b0000010011000001; // vC= 1217 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110000; // iC= 1136 
// vC = 14'b0000010100000101; // vC= 1285 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001111; // iC= 1167 
// vC = 14'b0000010101011111; // vC= 1375 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010100; // iC= 1300 
// vC = 14'b0000010010011100; // vC= 1180 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100111; // iC= 1127 
// vC = 14'b0000010001010000; // vC= 1104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010100; // iC= 1300 
// vC = 14'b0000010100100111; // vC= 1319 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100110; // iC= 1254 
// vC = 14'b0000010100001010; // vC= 1290 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100010; // iC= 1378 
// vC = 14'b0000010101110001; // vC= 1393 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110110; // iC= 1142 
// vC = 14'b0000010101101101; // vC= 1389 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111001; // iC= 1145 
// vC = 14'b0000010011101010; // vC= 1258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110100; // iC= 1332 
// vC = 14'b0000010101000110; // vC= 1350 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101001; // iC= 1065 
// vC = 14'b0000010010001101; // vC= 1165 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110001; // iC= 1265 
// vC = 14'b0000010011100001; // vC= 1249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100001; // iC= 1057 
// vC = 14'b0000010010101001; // vC= 1193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011100; // iC= 1180 
// vC = 14'b0000010110100010; // vC= 1442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001101; // iC= 1101 
// vC = 14'b0000010100010000; // vC= 1296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100101; // iC= 1317 
// vC = 14'b0000010101000011; // vC= 1347 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110000; // iC= 1328 
// vC = 14'b0000010100000000; // vC= 1280 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100111; // iC= 1319 
// vC = 14'b0000010100001000; // vC= 1288 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101111; // iC= 1071 
// vC = 14'b0000010101000101; // vC= 1349 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110000; // iC= 1008 
// vC = 14'b0000010101001110; // vC= 1358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100111; // iC=  999 
// vC = 14'b0000010011001100; // vC= 1228 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001100; // iC= 1228 
// vC = 14'b0000010111001101; // vC= 1485 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010111; // iC= 1239 
// vC = 14'b0000010101101001; // vC= 1385 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111000; // iC= 1144 
// vC = 14'b0000010011110101; // vC= 1269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011110; // iC= 1118 
// vC = 14'b0000010111000110; // vC= 1478 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100000; // iC= 1184 
// vC = 14'b0000010111000001; // vC= 1473 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111111; // iC= 1087 
// vC = 14'b0000010111010101; // vC= 1493 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101100; // iC= 1068 
// vC = 14'b0000010011101101; // vC= 1261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000001; // iC= 1153 
// vC = 14'b0000010110101101; // vC= 1453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010111; // iC= 1111 
// vC = 14'b0000010111000001; // vC= 1473 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110011; // iC= 1139 
// vC = 14'b0000010101100100; // vC= 1380 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011100; // iC=  988 
// vC = 14'b0000010101010100; // vC= 1364 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011111; // iC= 1055 
// vC = 14'b0000010110100111; // vC= 1447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101111; // iC= 1007 
// vC = 14'b0000010110010100; // vC= 1428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110001; // iC=  945 
// vC = 14'b0000010011101101; // vC= 1261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000111; // iC=  967 
// vC = 14'b0000010101011111; // vC= 1375 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000110; // iC= 1158 
// vC = 14'b0000010101110011; // vC= 1395 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111110; // iC= 1086 
// vC = 14'b0000010100110111; // vC= 1335 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100010; // iC=  930 
// vC = 14'b0000010100000010; // vC= 1282 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110100; // iC=  948 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111010; // iC= 1082 
// vC = 14'b0000010110111100; // vC= 1468 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010101; // iC=  853 
// vC = 14'b0000010100111000; // vC= 1336 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101101; // iC=  941 
// vC = 14'b0000010100110110; // vC= 1334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011100; // iC=  988 
// vC = 14'b0000010101001110; // vC= 1358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010000; // iC= 1104 
// vC = 14'b0000010100101100; // vC= 1324 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010011; // iC=  979 
// vC = 14'b0000010110011010; // vC= 1434 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001110; // iC=  846 
// vC = 14'b0000010100110000; // vC= 1328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101100; // iC= 1068 
// vC = 14'b0000011000011100; // vC= 1564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110101; // iC= 1077 
// vC = 14'b0000010111111101; // vC= 1533 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101001; // iC=  873 
// vC = 14'b0000010100111101; // vC= 1341 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101010; // iC=  938 
// vC = 14'b0000010101110100; // vC= 1396 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100001; // iC=  865 
// vC = 14'b0000011000100001; // vC= 1569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100011; // iC= 1059 
// vC = 14'b0000010100010000; // vC= 1296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110111; // iC=  823 
// vC = 14'b0000011000011111; // vC= 1567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001001; // iC=  905 
// vC = 14'b0000010111110010; // vC= 1522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001111; // iC=  783 
// vC = 14'b0000010100011011; // vC= 1307 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101011; // iC= 1067 
// vC = 14'b0000010111000011; // vC= 1475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000110; // iC=  838 
// vC = 14'b0000010100101010; // vC= 1322 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111011; // iC=  827 
// vC = 14'b0000010101100100; // vC= 1380 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011110; // iC= 1054 
// vC = 14'b0000010101010100; // vC= 1364 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001101; // iC=  973 
// vC = 14'b0000011000000101; // vC= 1541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110111; // iC= 1015 
// vC = 14'b0000010110101010; // vC= 1450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001010; // iC=  714 
// vC = 14'b0000010100111001; // vC= 1337 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001110; // iC=  846 
// vC = 14'b0000011000100011; // vC= 1571 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110110; // iC=  822 
// vC = 14'b0000010110110000; // vC= 1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001101; // iC=  845 
// vC = 14'b0000010101010001; // vC= 1361 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101000; // iC=  936 
// vC = 14'b0000011000111110; // vC= 1598 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011111; // iC=  799 
// vC = 14'b0000011001000001; // vC= 1601 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000111; // iC=  839 
// vC = 14'b0000010110110100; // vC= 1460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010110; // iC=  982 
// vC = 14'b0000010101100010; // vC= 1378 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111000; // iC=  888 
// vC = 14'b0000011001111100; // vC= 1660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111001; // iC=  889 
// vC = 14'b0000011001101110; // vC= 1646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111110; // iC=  702 
// vC = 14'b0000010101110000; // vC= 1392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001111; // iC=  847 
// vC = 14'b0000010101101111; // vC= 1391 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101010; // iC=  874 
// vC = 14'b0000011000000001; // vC= 1537 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000010; // iC=  706 
// vC = 14'b0000011010011011; // vC= 1691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110111; // iC=  823 
// vC = 14'b0000011000111110; // vC= 1598 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001101; // iC=  909 
// vC = 14'b0000010110101101; // vC= 1453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011100; // iC=  860 
// vC = 14'b0000010101111000; // vC= 1400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101101; // iC=  685 
// vC = 14'b0000010110100111; // vC= 1447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101110; // iC=  750 
// vC = 14'b0000010111100111; // vC= 1511 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001000; // iC=  584 
// vC = 14'b0000011010101100; // vC= 1708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110001; // iC=  753 
// vC = 14'b0000010110010110; // vC= 1430 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111001; // iC=  633 
// vC = 14'b0000010111000010; // vC= 1474 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010110; // iC=  790 
// vC = 14'b0000011000101101; // vC= 1581 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011010; // iC=  730 
// vC = 14'b0000011000110011; // vC= 1587 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110111; // iC=  631 
// vC = 14'b0000010111110011; // vC= 1523 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001010; // iC=  842 
// vC = 14'b0000011001010011; // vC= 1619 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001011; // iC=  651 
// vC = 14'b0000010110011010; // vC= 1434 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110000; // iC=  624 
// vC = 14'b0000011000000010; // vC= 1538 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000010; // iC=  834 
// vC = 14'b0000011000101100; // vC= 1580 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000011; // iC=  707 
// vC = 14'b0000011010100011; // vC= 1699 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000101; // iC=  517 
// vC = 14'b0000011001100111; // vC= 1639 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100000; // iC=  544 
// vC = 14'b0000011000110000; // vC= 1584 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101011; // iC=  747 
// vC = 14'b0000011010010010; // vC= 1682 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100001; // iC=  609 
// vC = 14'b0000010111100101; // vC= 1509 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111000; // iC=  568 
// vC = 14'b0000011001111010; // vC= 1658 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110011; // iC=  499 
// vC = 14'b0000011011010011; // vC= 1747 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110110; // iC=  630 
// vC = 14'b0000011001001011; // vC= 1611 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100111; // iC=  615 
// vC = 14'b0000011001010101; // vC= 1621 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010000; // iC=  592 
// vC = 14'b0000010111011011; // vC= 1499 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111111; // iC=  575 
// vC = 14'b0000010111100001; // vC= 1505 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110010; // iC=  626 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110110; // iC=  438 
// vC = 14'b0000011001111110; // vC= 1662 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111000; // iC=  696 
// vC = 14'b0000011000010110; // vC= 1558 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111000; // iC=  504 
// vC = 14'b0000011010110011; // vC= 1715 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101000; // iC=  424 
// vC = 14'b0000010110101111; // vC= 1455 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011111; // iC=  607 
// vC = 14'b0000011000011011; // vC= 1563 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000011; // iC=  579 
// vC = 14'b0000011001011011; // vC= 1627 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011100; // iC=  540 
// vC = 14'b0000011000000010; // vC= 1538 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111011; // iC=  379 
// vC = 14'b0000010111001100; // vC= 1484 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011001; // iC=  409 
// vC = 14'b0000011011000111; // vC= 1735 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001101; // iC=  461 
// vC = 14'b0000011001000000; // vC= 1600 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000101; // iC=  325 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000101; // iC=  581 
// vC = 14'b0000011011001100; // vC= 1740 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011101; // iC=  349 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100011; // iC=  483 
// vC = 14'b0000011001010111; // vC= 1623 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111010; // iC=  442 
// vC = 14'b0000011011111011; // vC= 1787 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111100; // iC=  252 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100100; // iC=  420 
// vC = 14'b0000011001100111; // vC= 1639 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010111; // iC=  407 
// vC = 14'b0000011001001110; // vC= 1614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110011; // iC=  179 
// vC = 14'b0000011010100100; // vC= 1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100111; // iC=  359 
// vC = 14'b0000011011000000; // vC= 1728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110000; // iC=  304 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111110; // iC=  318 
// vC = 14'b0000011010000001; // vC= 1665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001000; // iC=  264 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010100; // iC=  404 
// vC = 14'b0000010111111111; // vC= 1535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110111; // iC=  119 
// vC = 14'b0000011000001001; // vC= 1545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000111; // iC=  263 
// vC = 14'b0000011011011111; // vC= 1759 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110010; // iC=  178 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101100; // iC=  108 
// vC = 14'b0000011001001111; // vC= 1615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001101; // iC=  141 
// vC = 14'b0000011000110001; // vC= 1585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011101; // iC=  157 
// vC = 14'b0000011001000100; // vC= 1604 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001100; // iC=   76 
// vC = 14'b0000010111100011; // vC= 1507 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100111; // iC=  103 
// vC = 14'b0000011000000100; // vC= 1540 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110000; // iC=  240 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101100; // iC=  108 
// vC = 14'b0000011001010100; // vC= 1620 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000110001; // iC=   49 
// vC = 14'b0000010111111101; // vC= 1533 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110101111; // iC=  -81 
// vC = 14'b0000011010001110; // vC= 1678 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010100; // iC=   20 
// vC = 14'b0000011000010001; // vC= 1553 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100011; // iC=  -29 
// vC = 14'b0000011001000100; // vC= 1604 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100010; // iC=   98 
// vC = 14'b0000011000101111; // vC= 1583 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010110; // iC=  -42 
// vC = 14'b0000011011011011; // vC= 1755 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101000; // iC= -152 
// vC = 14'b0000011011100001; // vC= 1761 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101001; // iC=   41 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011100; // iC= -228 
// vC = 14'b0000011011001100; // vC= 1740 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011101; // iC=  -99 
// vC = 14'b0000011001100000; // vC= 1632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000000; // iC= -192 
// vC = 14'b0000011001011000; // vC= 1624 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010011; // iC= -301 
// vC = 14'b0000011000011111; // vC= 1567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110110; // iC= -330 
// vC = 14'b0000010111100101; // vC= 1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101101; // iC= -211 
// vC = 14'b0000011010000111; // vC= 1671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010111; // iC= -169 
// vC = 14'b0000011001110111; // vC= 1655 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011110111; // iC= -265 
// vC = 14'b0000011010111000; // vC= 1720 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010011; // iC= -365 
// vC = 14'b0000011010000001; // vC= 1665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100010; // iC= -158 
// vC = 14'b0000011000110011; // vC= 1587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110011; // iC= -205 
// vC = 14'b0000011011000110; // vC= 1734 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010101; // iC= -235 
// vC = 14'b0000011010011100; // vC= 1692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101000; // iC= -536 
// vC = 14'b0000011000001110; // vC= 1550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110010; // iC= -462 
// vC = 14'b0000011001000110; // vC= 1606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111101; // iC= -579 
// vC = 14'b0000010111010110; // vC= 1494 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110110; // iC= -458 
// vC = 14'b0000011011010000; // vC= 1744 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011011; // iC= -485 
// vC = 14'b0000011010100000; // vC= 1696 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101100; // iC= -468 
// vC = 14'b0000010111000111; // vC= 1479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011001; // iC= -551 
// vC = 14'b0000011011000000; // vC= 1728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011011; // iC= -613 
// vC = 14'b0000011000010001; // vC= 1553 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110010; // iC= -718 
// vC = 14'b0000011001001110; // vC= 1614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010011; // iC= -557 
// vC = 14'b0000011010010001; // vC= 1681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111011; // iC= -453 
// vC = 14'b0000010110110100; // vC= 1460 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000101; // iC= -763 
// vC = 14'b0000010111010111; // vC= 1495 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011100; // iC= -804 
// vC = 14'b0000010111010111; // vC= 1495 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010001; // iC= -623 
// vC = 14'b0000010111111001; // vC= 1529 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010000; // iC= -624 
// vC = 14'b0000011011010111; // vC= 1751 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011001; // iC= -807 
// vC = 14'b0000011000110110; // vC= 1590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000011; // iC= -829 
// vC = 14'b0000010111110000; // vC= 1520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100011; // iC= -733 
// vC = 14'b0000011000101000; // vC= 1576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010001; // iC= -815 
// vC = 14'b0000011000101101; // vC= 1581 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011100; // iC= -740 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101100; // iC= -724 
// vC = 14'b0000011000110110; // vC= 1590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000011; // iC= -829 
// vC = 14'b0000010110100011; // vC= 1443 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111111; // iC=-1025 
// vC = 14'b0000011001001111; // vC= 1615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001010; // iC= -822 
// vC = 14'b0000010111100001; // vC= 1505 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101010; // iC=-1046 
// vC = 14'b0000010110101011; // vC= 1451 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010000; // iC= -944 
// vC = 14'b0000010111010100; // vC= 1492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011000; // iC=-1000 
// vC = 14'b0000010101111111; // vC= 1407 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010010; // iC= -814 
// vC = 14'b0000010110000001; // vC= 1409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111100; // iC= -836 
// vC = 14'b0000010111010101; // vC= 1493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111100; // iC=-1092 
// vC = 14'b0000011001000100; // vC= 1604 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000111; // iC= -953 
// vC = 14'b0000010111010101; // vC= 1493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001010; // iC=-1078 
// vC = 14'b0000010110100100; // vC= 1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100000; // iC=-1184 
// vC = 14'b0000010111100100; // vC= 1508 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011011; // iC= -997 
// vC = 14'b0000010110010010; // vC= 1426 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001111; // iC=-1073 
// vC = 14'b0000011001100010; // vC= 1634 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011101; // iC=-1059 
// vC = 14'b0000010101100110; // vC= 1382 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010101; // iC=-1003 
// vC = 14'b0000011000100011; // vC= 1571 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100110; // iC=-1306 
// vC = 14'b0000010101010000; // vC= 1360 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110101; // iC=-1099 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110000; // iC=-1104 
// vC = 14'b0000010101010001; // vC= 1361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100100; // iC=-1116 
// vC = 14'b0000010101010110; // vC= 1366 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101110; // iC=-1234 
// vC = 14'b0000010101100100; // vC= 1380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111110; // iC=-1410 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110111; // iC=-1289 
// vC = 14'b0000010101000001; // vC= 1345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000011; // iC=-1405 
// vC = 14'b0000010100110111; // vC= 1335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110101; // iC=-1355 
// vC = 14'b0000010111111011; // vC= 1531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110011; // iC=-1421 
// vC = 14'b0000010110011100; // vC= 1436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111110; // iC=-1410 
// vC = 14'b0000010110111010; // vC= 1466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111001; // iC=-1351 
// vC = 14'b0000011000110011; // vC= 1587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100001; // iC=-1311 
// vC = 14'b0000010100001011; // vC= 1291 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101100; // iC=-1492 
// vC = 14'b0000010101100001; // vC= 1377 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101000; // iC=-1432 
// vC = 14'b0000010101000011; // vC= 1347 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110101; // iC=-1355 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101011; // iC=-1429 
// vC = 14'b0000010110000101; // vC= 1413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111001; // iC=-1415 
// vC = 14'b0000010111011100; // vC= 1500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110011; // iC=-1421 
// vC = 14'b0000010100000100; // vC= 1284 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011100; // iC=-1508 
// vC = 14'b0000010111001111; // vC= 1487 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111101; // iC=-1603 
// vC = 14'b0000010110000110; // vC= 1414 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011111; // iC=-1377 
// vC = 14'b0000010101011011; // vC= 1371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110010; // iC=-1550 
// vC = 14'b0000010101111111; // vC= 1407 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101100; // iC=-1556 
// vC = 14'b0000010110000001; // vC= 1409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001100; // iC=-1588 
// vC = 14'b0000010101111100; // vC= 1404 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011100; // iC=-1444 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001011; // iC=-1461 
// vC = 14'b0000010010111110; // vC= 1214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010101; // iC=-1451 
// vC = 14'b0000010111001101; // vC= 1485 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100111; // iC=-1561 
// vC = 14'b0000010011100001; // vC= 1249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001111; // iC=-1649 
// vC = 14'b0000010010010100; // vC= 1172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110011; // iC=-1677 
// vC = 14'b0000010110100000; // vC= 1440 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001101; // iC=-1779 
// vC = 14'b0000010101000100; // vC= 1348 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000011; // iC=-1789 
// vC = 14'b0000010100101111; // vC= 1327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010000; // iC=-1648 
// vC = 14'b0000010010001001; // vC= 1161 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101010; // iC=-1686 
// vC = 14'b0000010110011001; // vC= 1433 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101101; // iC=-1555 
// vC = 14'b0000010001100000; // vC= 1120 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000111; // iC=-1721 
// vC = 14'b0000010001010001; // vC= 1105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111010; // iC=-1670 
// vC = 14'b0000010010000011; // vC= 1155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101111; // iC=-1617 
// vC = 14'b0000010011000001; // vC= 1217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000010; // iC=-1662 
// vC = 14'b0000010011100110; // vC= 1254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011000; // iC=-1640 
// vC = 14'b0000010100100001; // vC= 1313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011111; // iC=-1761 
// vC = 14'b0000010100110111; // vC= 1335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000011; // iC=-1725 
// vC = 14'b0000010010101011; // vC= 1195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010011; // iC=-1645 
// vC = 14'b0000010101011010; // vC= 1370 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000111; // iC=-1785 
// vC = 14'b0000010000110010; // vC= 1074 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100101; // iC=-1691 
// vC = 14'b0000010010001010; // vC= 1162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011010; // iC=-1638 
// vC = 14'b0000010011111111; // vC= 1279 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000101; // iC=-1659 
// vC = 14'b0000010000000111; // vC= 1031 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011001; // iC=-1895 
// vC = 14'b0000010000000100; // vC= 1028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011100; // iC=-1636 
// vC = 14'b0000010010001000; // vC= 1160 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011110; // iC=-1762 
// vC = 14'b0000010000100000; // vC= 1056 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001110; // iC=-1842 
// vC = 14'b0000001111011100; // vC=  988 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110010; // iC=-1742 
// vC = 14'b0000010000101011; // vC= 1067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000100; // iC=-1660 
// vC = 14'b0000010011110100; // vC= 1268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b0000010011111011; // vC= 1275 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b0000001110110110; // vC=  950 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000101; // iC=-1915 
// vC = 14'b0000010011011001; // vC= 1241 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001100; // iC=-1716 
// vC = 14'b0000001111010000; // vC=  976 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110100; // iC=-1740 
// vC = 14'b0000010010100010; // vC= 1186 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000010010111110; // vC= 1214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111111; // iC=-1921 
// vC = 14'b0000001111011101; // vC=  989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011110; // iC=-1698 
// vC = 14'b0000001111100100; // vC=  996 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b0000010010100010; // vC= 1186 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011011; // iC=-1829 
// vC = 14'b0000001111101011; // vC= 1003 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b0000010001011001; // vC= 1113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000000; // iC=-1792 
// vC = 14'b0000001111110001; // vC= 1009 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b0000001110100011; // vC=  931 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100010; // iC=-1886 
// vC = 14'b0000001101111101; // vC=  893 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000110; // iC=-1722 
// vC = 14'b0000001110111011; // vC=  955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011001; // iC=-1895 
// vC = 14'b0000001111100101; // vC=  997 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100111; // iC=-1945 
// vC = 14'b0000001111100010; // vC=  994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b0000001110111111; // vC=  959 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b0000001101100010; // vC=  866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b0000001101001110; // vC=  846 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010001; // iC=-1839 
// vC = 14'b0000010001010010; // vC= 1106 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100000; // iC=-1760 
// vC = 14'b0000001111001011; // vC=  971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010000; // iC=-1904 
// vC = 14'b0000001111011001; // vC=  985 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110101; // iC=-1867 
// vC = 14'b0000010000111100; // vC= 1084 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b0000001100110110; // vC=  822 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111001; // iC=-1799 
// vC = 14'b0000001110011100; // vC=  924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111111; // iC=-1793 
// vC = 14'b0000001100110000; // vC=  816 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010111; // iC=-1833 
// vC = 14'b0000001110001011; // vC=  907 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b0000001100001000; // vC=  776 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011110; // iC=-1826 
// vC = 14'b0000001110010111; // vC=  919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b0000001110110000; // vC=  944 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001101; // iC=-2035 
// vC = 14'b0000001101100111; // vC=  871 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b0000001111110100; // vC= 1012 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b0000001101100110; // vC=  870 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000100; // iC=-1852 
// vC = 14'b0000001101100010; // vC=  866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b0000001110110000; // vC=  944 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010010; // iC=-1966 
// vC = 14'b0000001110111101; // vC=  957 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011110; // iC=-2082 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110011; // iC=-1805 
// vC = 14'b0000001101000100; // vC=  836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b0000001110000011; // vC=  899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b0000001010010111; // vC=  663 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000101; // iC=-2043 
// vC = 14'b0000001100011111; // vC=  799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000001011000001; // vC=  705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101110; // iC=-1810 
// vC = 14'b0000001101010101; // vC=  853 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b0000001101101111; // vC=  879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000001100111100; // vC=  828 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000001001001111; // vC=  591 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110101; // iC=-1867 
// vC = 14'b0000001011011010; // vC=  730 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b0000001001000011; // vC=  579 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b0000001000101010; // vC=  554 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000001001110001; // vC=  625 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001010; // iC=-1910 
// vC = 14'b0000001101000100; // vC=  836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011100; // iC=-1892 
// vC = 14'b0000001000101111; // vC=  559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011000; // iC=-2024 
// vC = 14'b0000001010110111; // vC=  695 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100111; // iC=-1945 
// vC = 14'b0000001011101111; // vC=  751 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b0000001001111101; // vC=  637 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b0000001001110001; // vC=  625 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b0000001000000000; // vC=  512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000001010110011; // vC=  691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010100; // iC=-1900 
// vC = 14'b0000001000000001; // vC=  513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b0000000111010010; // vC=  466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b0000001001010000; // vC=  592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b0000001001101111; // vC=  623 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b0000000110100110; // vC=  422 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000001000001001; // vC=  521 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101001; // iC=-2071 
// vC = 14'b0000001001010011; // vC=  595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b0000001001011100; // vC=  604 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b0000000110010111; // vC=  407 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110000; // iC=-1936 
// vC = 14'b0000000111111100; // vC=  508 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010000; // iC=-2096 
// vC = 14'b0000001000011000; // vC=  536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b0000000111111000; // vC=  504 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000101; // iC=-1787 
// vC = 14'b0000001000110001; // vC=  561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010101; // iC=-2027 
// vC = 14'b0000000101101011; // vC=  363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b0000001001000011; // vC=  579 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b0000001001000011; // vC=  579 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010100; // iC=-2092 
// vC = 14'b0000000111101000; // vC=  488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b0000000111101101; // vC=  493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b0000000101000001; // vC=  321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b0000000101100011; // vC=  355 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000000101100111; // vC=  359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b0000000100010101; // vC=  277 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b0000001000000111; // vC=  519 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b0000000101110101; // vC=  373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b0000000110110100; // vC=  436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000000111001100; // vC=  460 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000000011101010; // vC=  234 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001110; // iC=-1906 
// vC = 14'b0000000100011010; // vC=  282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000101; // iC=-1851 
// vC = 14'b0000000110110100; // vC=  436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000111; // iC=-1913 
// vC = 14'b0000000110001110; // vC=  398 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001101; // iC=-2035 
// vC = 14'b0000000110110110; // vC=  438 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b0000000011110011; // vC=  243 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b0000000100001110; // vC=  270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b0000000110011111; // vC=  415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000000011011101; // vC=  221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111101; // iC=-1923 
// vC = 14'b0000000101011000; // vC=  344 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b0000000011100010; // vC=  226 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b0000000101110110; // vC=  374 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011011; // iC=-2085 
// vC = 14'b0000000101111010; // vC=  378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000000; // iC=-1792 
// vC = 14'b0000000100101111; // vC=  303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000010; // iC=-1854 
// vC = 14'b0000000101101011; // vC=  363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001001; // iC=-1847 
// vC = 14'b0000000010110010; // vC=  178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b0000000110010111; // vC=  407 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000000010110100; // vC=  180 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b0000000100010000; // vC=  272 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011011; // iC=-1829 
// vC = 14'b0000000011001001; // vC=  201 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b0000000101100011; // vC=  355 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011001; // iC=-1831 
// vC = 14'b0000000101000010; // vC=  322 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011100; // iC=-1892 
// vC = 14'b0000000010011001; // vC=  153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110011; // iC=-1997 
// vC = 14'b0000000101001001; // vC=  329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011000; // iC=-1896 
// vC = 14'b0000000000100110; // vC=   38 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010010; // iC=-1966 
// vC = 14'b0000000010101100; // vC=  172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110001; // iC=-1807 
// vC = 14'b0000000101010001; // vC=  337 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000000101001110; // vC=  334 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111100; // iC=-1988 
// vC = 14'b0000000100001110; // vC=  270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000110; // iC=-1786 
// vC = 14'b0000000010001011; // vC=  139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b0000000001100101; // vC=  101 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b1111111111110101; // vC=  -11 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b0000000010011111; // vC=  159 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b1111111111111011; // vC=   -5 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011000; // iC=-2088 
// vC = 14'b0000000000110010; // vC=   50 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b1111111111101010; // vC=  -22 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010100; // iC=-1772 
// vC = 14'b1111111111110000; // vC=  -16 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b1111111111100101; // vC=  -27 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010111; // iC=-1897 
// vC = 14'b0000000001100011; // vC=   99 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b0000000010111010; // vC=  186 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b1111111111000110; // vC=  -58 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011110; // iC=-2082 
// vC = 14'b1111111110100010; // vC=  -94 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b0000000010111111; // vC=  191 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110010; // iC=-1806 
// vC = 14'b0000000001110110; // vC=  118 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000110; // iC=-1914 
// vC = 14'b1111111110001101; // vC= -115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b1111111111000101; // vC=  -59 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010110; // iC=-1962 
// vC = 14'b0000000010001010; // vC=  138 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101111; // iC=-1937 
// vC = 14'b0000000001001011; // vC=   75 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b1111111110110000; // vC=  -80 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010111; // iC=-1897 
// vC = 14'b1111111101100000; // vC= -160 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110000; // iC=-1936 
// vC = 14'b0000000001001101; // vC=   77 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101010; // iC=-2070 
// vC = 14'b0000000000110000; // vC=   48 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000101; // iC=-2043 
// vC = 14'b0000000000111010; // vC=   58 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010010; // iC=-1774 
// vC = 14'b1111111101101010; // vC= -150 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110001; // iC=-2063 
// vC = 14'b1111111110001110; // vC= -114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b0000000000010111; // vC=   23 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101001; // iC=-1879 
// vC = 14'b1111111110011001; // vC= -103 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011000; // iC=-2024 
// vC = 14'b1111111110000011; // vC= -125 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000100; // iC=-2044 
// vC = 14'b1111111101011110; // vC= -162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b1111111111111101; // vC=   -3 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001111; // iC=-1777 
// vC = 14'b1111111101111010; // vC= -134 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b1111111111001110; // vC=  -50 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b1111111100110111; // vC= -201 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011111; // iC=-1825 
// vC = 14'b1111111011101000; // vC= -280 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b1111111101100001; // vC= -159 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010101; // iC=-1835 
// vC = 14'b0000000000000111; // vC=    7 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b1111111111111011; // vC=   -5 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110001; // iC=-1935 
// vC = 14'b1111111100111010; // vC= -198 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001001; // iC=-1847 
// vC = 14'b1111111011101000; // vC= -280 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101111; // iC=-1809 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110010; // iC=-1742 
// vC = 14'b1111111101100110; // vC= -154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100000; // iC=-2016 
// vC = 14'b1111111010100111; // vC= -345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b1111111110001111; // vC= -113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100010; // iC=-1758 
// vC = 14'b1111111110111110; // vC=  -66 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101001; // iC=-2007 
// vC = 14'b1111111010100011; // vC= -349 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000100; // iC=-1916 
// vC = 14'b1111111100110011; // vC= -205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b1111111100110011; // vC= -205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111001; // iC=-1735 
// vC = 14'b1111111100001111; // vC= -241 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111100; // iC=-1796 
// vC = 14'b1111111101111010; // vC= -134 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b1111111100100010; // vC= -222 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100111; // iC=-1753 
// vC = 14'b1111111010110001; // vC= -335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b1111111101000111; // vC= -185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b1111111100000100; // vC= -252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101111; // iC=-1873 
// vC = 14'b1111111001010111; // vC= -425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b1111111001100111; // vC= -409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100000; // iC=-1824 
// vC = 14'b1111111101011111; // vC= -161 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110011; // iC=-1869 
// vC = 14'b1111111101010001; // vC= -175 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b1111111100010100; // vC= -236 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000000; // iC=-1792 
// vC = 14'b1111111000011011; // vC= -485 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b1111111001101110; // vC= -402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011000; // iC=-1896 
// vC = 14'b1111111010011110; // vC= -354 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011111; // iC=-1953 
// vC = 14'b1111111000111100; // vC= -452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001000; // iC=-1784 
// vC = 14'b1111111100111000; // vC= -200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110101; // iC=-1803 
// vC = 14'b1111111100100010; // vC= -222 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b1111111000111111; // vC= -449 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111111010000111; // vC= -377 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b1111111000010101; // vC= -491 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100101; // iC=-1819 
// vC = 14'b1111111010100011; // vC= -349 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b1111110111011000; // vC= -552 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111011; // iC=-1733 
// vC = 14'b1111111011000001; // vC= -319 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101001; // iC=-1879 
// vC = 14'b1111111011001000; // vC= -312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100011; // iC=-1693 
// vC = 14'b1111110111111010; // vC= -518 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011011; // iC=-1765 
// vC = 14'b1111111010010111; // vC= -361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b1111111011011000; // vC= -296 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000001; // iC=-1791 
// vC = 14'b1111110110110010; // vC= -590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b1111110111101100; // vC= -532 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011010; // iC=-1894 
// vC = 14'b1111111001110101; // vC= -395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100111; // iC=-1881 
// vC = 14'b1111111000001011; // vC= -501 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101000; // iC=-1752 
// vC = 14'b1111111000100111; // vC= -473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101011; // iC=-1877 
// vC = 14'b1111110111101001; // vC= -535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000101; // iC=-1787 
// vC = 14'b1111110111011010; // vC= -550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b1111110110100010; // vC= -606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101000; // iC=-1688 
// vC = 14'b1111111000010101; // vC= -491 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000110; // iC=-1914 
// vC = 14'b1111110111000100; // vC= -572 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001011; // iC=-1717 
// vC = 14'b1111111000010100; // vC= -492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101010; // iC=-1878 
// vC = 14'b1111110111111101; // vC= -515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b1111110111101000; // vC= -536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010011; // iC=-1709 
// vC = 14'b1111110101000001; // vC= -703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010110; // iC=-1834 
// vC = 14'b1111110111000100; // vC= -572 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b1111110111010001; // vC= -559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010111; // iC=-1641 
// vC = 14'b1111110111101100; // vC= -532 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110101; // iC=-1611 
// vC = 14'b1111111000001101; // vC= -499 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b1111110111001011; // vC= -565 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000000; // iC=-1728 
// vC = 14'b1111111000111010; // vC= -454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100001; // iC=-1887 
// vC = 14'b1111110111110011; // vC= -525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101010; // iC=-1750 
// vC = 14'b1111110101011001; // vC= -679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111000; // iC=-1736 
// vC = 14'b1111110100010000; // vC= -752 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110110; // iC=-1802 
// vC = 14'b1111110100111000; // vC= -712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101111; // iC=-1681 
// vC = 14'b1111110100100010; // vC= -734 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001111; // iC=-1777 
// vC = 14'b1111110011110100; // vC= -780 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000111; // iC=-1785 
// vC = 14'b1111110111000010; // vC= -574 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b1111110111101111; // vC= -529 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000001; // iC=-1663 
// vC = 14'b1111110011111010; // vC= -774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101110; // iC=-1746 
// vC = 14'b1111110110100110; // vC= -602 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010100; // iC=-1772 
// vC = 14'b1111110110101010; // vC= -598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000000; // iC=-1792 
// vC = 14'b1111110110101010; // vC= -598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001100; // iC=-1652 
// vC = 14'b1111110011111001; // vC= -775 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110110; // iC=-1738 
// vC = 14'b1111110010110101; // vC= -843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110011; // iC=-1613 
// vC = 14'b1111110010100000; // vC= -864 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011010; // iC=-1638 
// vC = 14'b1111110110001010; // vC= -630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b1111110111001001; // vC= -567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111111; // iC=-1729 
// vC = 14'b1111110011110110; // vC= -778 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b1111110001111100; // vC= -900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010101; // iC=-1771 
// vC = 14'b1111110101001101; // vC= -691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011101; // iC=-1635 
// vC = 14'b1111110110011011; // vC= -613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110110; // iC=-1674 
// vC = 14'b1111110010000100; // vC= -892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110110; // iC=-1674 
// vC = 14'b1111110101111010; // vC= -646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000000; // iC=-1536 
// vC = 14'b1111110011011100; // vC= -804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b1111110001100011; // vC= -925 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b1111110001100011; // vC= -925 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100101; // iC=-1627 
// vC = 14'b1111110101101011; // vC= -661 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b1111110101010101; // vC= -683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011111; // iC=-1633 
// vC = 14'b1111110101000000; // vC= -704 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011110; // iC=-1698 
// vC = 14'b1111110010100011; // vC= -861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010101; // iC=-1643 
// vC = 14'b1111110101100111; // vC= -665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101001; // iC=-1559 
// vC = 14'b1111110100111000; // vC= -712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011111; // iC=-1761 
// vC = 14'b1111110101001100; // vC= -692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101111; // iC=-1681 
// vC = 14'b1111110011100111; // vC= -793 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110001; // iC=-1807 
// vC = 14'b1111110100000100; // vC= -764 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111000; // iC=-1736 
// vC = 14'b1111110000100101; // vC= -987 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111010; // iC=-1798 
// vC = 14'b1111110011010100; // vC= -812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111101; // iC=-1731 
// vC = 14'b1111110011001110; // vC= -818 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011110; // iC=-1762 
// vC = 14'b1111110100011011; // vC= -741 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100010; // iC=-1758 
// vC = 14'b1111110100000011; // vC= -765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110011; // iC=-1549 
// vC = 14'b1111101111101100; // vC=-1044 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000110; // iC=-1658 
// vC = 14'b1111110010000111; // vC= -889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110111; // iC=-1545 
// vC = 14'b1111101111010101; // vC=-1067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011001; // iC=-1511 
// vC = 14'b1111110011111011; // vC= -773 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100111; // iC=-1689 
// vC = 14'b1111101111010111; // vC=-1065 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011110; // iC=-1570 
// vC = 14'b1111110011000111; // vC= -825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b1111110001110100; // vC= -908 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111101; // iC=-1731 
// vC = 14'b1111101111001001; // vC=-1079 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011011; // iC=-1765 
// vC = 14'b1111110011001110; // vC= -818 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010011; // iC=-1581 
// vC = 14'b1111110000001111; // vC=-1009 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010101; // iC=-1643 
// vC = 14'b1111101111111100; // vC=-1028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101001; // iC=-1623 
// vC = 14'b1111110010101110; // vC= -850 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010010; // iC=-1582 
// vC = 14'b1111110001110000; // vC= -912 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010010; // iC=-1582 
// vC = 14'b1111110001010100; // vC= -940 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000000; // iC=-1472 
// vC = 14'b1111110010000001; // vC= -895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110001; // iC=-1487 
// vC = 14'b1111110001101100; // vC= -916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011000; // iC=-1512 
// vC = 14'b1111101110001010; // vC=-1142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001100; // iC=-1716 
// vC = 14'b1111110000001100; // vC=-1012 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011010; // iC=-1446 
// vC = 14'b1111110001110001; // vC= -911 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111101; // iC=-1411 
// vC = 14'b1111101110011110; // vC=-1122 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110100; // iC=-1676 
// vC = 14'b1111110001100000; // vC= -928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011001; // iC=-1447 
// vC = 14'b1111101111001100; // vC=-1076 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011000; // iC=-1576 
// vC = 14'b1111101101111110; // vC=-1154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011001; // iC=-1447 
// vC = 14'b1111101111010010; // vC=-1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001011; // iC=-1461 
// vC = 14'b1111101110000110; // vC=-1146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001110; // iC=-1394 
// vC = 14'b1111101111101100; // vC=-1044 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110001; // iC=-1615 
// vC = 14'b1111110001101010; // vC= -918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011100; // iC=-1572 
// vC = 14'b1111101111110111; // vC=-1033 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101010; // iC=-1686 
// vC = 14'b1111101101001110; // vC=-1202 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110001; // iC=-1679 
// vC = 14'b1111101111001010; // vC=-1078 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101010; // iC=-1558 
// vC = 14'b1111101110111000; // vC=-1096 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000001; // iC=-1471 
// vC = 14'b1111101100100010; // vC=-1246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011010; // iC=-1510 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100011; // iC=-1501 
// vC = 14'b1111101111001111; // vC=-1073 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101010; // iC=-1622 
// vC = 14'b1111101100010000; // vC=-1264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000010; // iC=-1342 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110101; // iC=-1419 
// vC = 14'b1111101110000001; // vC=-1151 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101001; // iC=-1559 
// vC = 14'b1111101110001101; // vC=-1139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111010; // iC=-1350 
// vC = 14'b1111101100111101; // vC=-1219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001111; // iC=-1521 
// vC = 14'b1111101011101010; // vC=-1302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100000; // iC=-1504 
// vC = 14'b1111101110011011; // vC=-1125 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000011; // iC=-1597 
// vC = 14'b1111101011011011; // vC=-1317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101111; // iC=-1361 
// vC = 14'b1111101011100110; // vC=-1306 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101001; // iC=-1431 
// vC = 14'b1111110000000001; // vC=-1023 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001111; // iC=-1393 
// vC = 14'b1111101111101001; // vC=-1047 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010110; // iC=-1322 
// vC = 14'b1111101100001010; // vC=-1270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100011; // iC=-1565 
// vC = 14'b1111101011011100; // vC=-1316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110001; // iC=-1359 
// vC = 14'b1111101110101110; // vC=-1106 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110111; // iC=-1609 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010111; // iC=-1321 
// vC = 14'b1111101101101011; // vC=-1173 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111110; // iC=-1538 
// vC = 14'b1111101011001011; // vC=-1333 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111101; // iC=-1347 
// vC = 14'b1111101110010011; // vC=-1133 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001001; // iC=-1399 
// vC = 14'b1111101111000010; // vC=-1086 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010011; // iC=-1517 
// vC = 14'b1111101100010001; // vC=-1263 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110001; // iC=-1295 
// vC = 14'b1111101100011101; // vC=-1251 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000001; // iC=-1343 
// vC = 14'b1111101110110110; // vC=-1098 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000011; // iC=-1469 
// vC = 14'b1111101110001000; // vC=-1144 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101001; // iC=-1495 
// vC = 14'b1111101011111111; // vC=-1281 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101101; // iC=-1427 
// vC = 14'b1111101101010010; // vC=-1198 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011001; // iC=-1511 
// vC = 14'b1111101010011001; // vC=-1383 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110000; // iC=-1296 
// vC = 14'b1111101001101111; // vC=-1425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000111; // iC=-1465 
// vC = 14'b1111101011011001; // vC=-1319 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100001; // iC=-1311 
// vC = 14'b1111101010000101; // vC=-1403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111001; // iC=-1415 
// vC = 14'b1111101001101001; // vC=-1431 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000100; // iC=-1468 
// vC = 14'b1111101010001101; // vC=-1395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011010; // iC=-1318 
// vC = 14'b1111101010000111; // vC=-1401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111110; // iC=-1282 
// vC = 14'b1111101010010001; // vC=-1391 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011111; // iC=-1505 
// vC = 14'b1111101011110110; // vC=-1290 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101110; // iC=-1490 
// vC = 14'b1111101100000101; // vC=-1275 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100011; // iC=-1245 
// vC = 14'b1111101010110000; // vC=-1360 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000000; // iC=-1280 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010110; // iC=-1322 
// vC = 14'b1111101001001100; // vC=-1460 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000010; // iC=-1406 
// vC = 14'b1111101000101011; // vC=-1493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110001; // iC=-1487 
// vC = 14'b1111101011000110; // vC=-1338 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110010; // iC=-1422 
// vC = 14'b1111101100011111; // vC=-1249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100101; // iC=-1179 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100101; // iC=-1307 
// vC = 14'b1111101011100101; // vC=-1307 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100011; // iC=-1181 
// vC = 14'b1111101000100011; // vC=-1501 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011000; // iC=-1448 
// vC = 14'b1111101011111011; // vC=-1285 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001001; // iC=-1463 
// vC = 14'b1111101010000101; // vC=-1403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001111; // iC=-1201 
// vC = 14'b1111101010111110; // vC=-1346 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000001; // iC=-1215 
// vC = 14'b1111101100010001; // vC=-1263 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011001; // iC=-1447 
// vC = 14'b1111101001111100; // vC=-1412 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010000; // iC=-1200 
// vC = 14'b1111101011100011; // vC=-1309 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010000; // iC=-1136 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111011; // iC=-1157 
// vC = 14'b1111101100010011; // vC=-1261 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011110; // iC=-1122 
// vC = 14'b1111101100000001; // vC=-1279 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011111; // iC=-1249 
// vC = 14'b1111101010100110; // vC=-1370 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010010; // iC=-1262 
// vC = 14'b1111101011111110; // vC=-1282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101001; // iC=-1303 
// vC = 14'b1111101010000011; // vC=-1405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111100; // iC=-1284 
// vC = 14'b1111101010011001; // vC=-1383 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000011; // iC=-1149 
// vC = 14'b1111100111111010; // vC=-1542 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100010; // iC=-1310 
// vC = 14'b1111101001010001; // vC=-1455 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110011; // iC=-1165 
// vC = 14'b1111101010111001; // vC=-1351 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101010; // iC=-1110 
// vC = 14'b1111101000111100; // vC=-1476 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101011; // iC=-1109 
// vC = 14'b1111100111111110; // vC=-1538 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010110; // iC=-1322 
// vC = 14'b1111101000010001; // vC=-1519 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001110; // iC=-1330 
// vC = 14'b1111101000101110; // vC=-1490 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110101; // iC=-1163 
// vC = 14'b1111101000001010; // vC=-1526 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011110; // iC=-1186 
// vC = 14'b1111101010110100; // vC=-1356 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111101; // iC=-1091 
// vC = 14'b1111101010011011; // vC=-1381 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000111; // iC=-1273 
// vC = 14'b1111100111000110; // vC=-1594 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001011; // iC=-1141 
// vC = 14'b1111100110010010; // vC=-1646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110101; // iC=-1227 
// vC = 14'b1111101001111100; // vC=-1412 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010001; // iC=-1135 
// vC = 14'b1111100110010011; // vC=-1645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001100; // iC=-1012 
// vC = 14'b1111100110010110; // vC=-1642 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001110; // iC=-1074 
// vC = 14'b1111100111101011; // vC=-1557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000110; // iC=-1210 
// vC = 14'b1111100101111011; // vC=-1669 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010001; // iC=-1263 
// vC = 14'b1111101000001000; // vC=-1528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100101; // iC=-1243 
// vC = 14'b1111101001010000; // vC=-1456 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010010; // iC=-1070 
// vC = 14'b1111100101101001; // vC=-1687 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010101; // iC=-1003 
// vC = 14'b1111101000110100; // vC=-1484 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100010; // iC=-1182 
// vC = 14'b1111101001101110; // vC=-1426 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111110; // iC=-1154 
// vC = 14'b1111101000101010; // vC=-1494 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100011; // iC=-1245 
// vC = 14'b1111100111100011; // vC=-1565 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101010; // iC=-1174 
// vC = 14'b1111100110011011; // vC=-1637 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011110; // iC=-1250 
// vC = 14'b1111100111000001; // vC=-1599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001100; // iC= -948 
// vC = 14'b1111100111000110; // vC=-1594 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111111; // iC=-1025 
// vC = 14'b1111100101100110; // vC=-1690 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101110; // iC=-1042 
// vC = 14'b1111101000000011; // vC=-1533 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111000; // iC=-1096 
// vC = 14'b1111101000111101; // vC=-1475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100000; // iC=-1248 
// vC = 14'b1111100101100000; // vC=-1696 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001010; // iC= -950 
// vC = 14'b1111100101010101; // vC=-1707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011011; // iC=-1189 
// vC = 14'b1111100110110000; // vC=-1616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001101; // iC= -947 
// vC = 14'b1111100110010100; // vC=-1644 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110001; // iC= -975 
// vC = 14'b1111100110000000; // vC=-1664 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110000; // iC=-1168 
// vC = 14'b1111100111101001; // vC=-1559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100111; // iC=-1177 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101111; // iC=-1169 
// vC = 14'b1111101001001011; // vC=-1461 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010110; // iC=-1002 
// vC = 14'b1111100111001100; // vC=-1588 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010001; // iC=-1199 
// vC = 14'b1111100110101101; // vC=-1619 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011011; // iC= -933 
// vC = 14'b1111100101000101; // vC=-1723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110011; // iC=-1101 
// vC = 14'b1111100110110001; // vC=-1615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101110; // iC=-1106 
// vC = 14'b1111100110010011; // vC=-1645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010111; // iC=-1065 
// vC = 14'b1111101000000100; // vC=-1532 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101001; // iC=-1047 
// vC = 14'b1111100101000110; // vC=-1722 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110011; // iC=-1037 
// vC = 14'b1111100100011110; // vC=-1762 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010001; // iC= -943 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100101; // iC= -923 
// vC = 14'b1111100111011101; // vC=-1571 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111100; // iC=-1028 
// vC = 14'b1111100101000001; // vC=-1727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110001; // iC= -847 
// vC = 14'b1111100011100001; // vC=-1823 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b1111100100110110; // vC=-1738 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111100; // iC= -836 
// vC = 14'b1111100111011111; // vC=-1569 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100000; // iC=-1120 
// vC = 14'b1111100101000001; // vC=-1727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011011; // iC= -933 
// vC = 14'b1111100100101100; // vC=-1748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010000; // iC= -944 
// vC = 14'b1111100110010001; // vC=-1647 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100000; // iC=-1056 
// vC = 14'b1111101000000111; // vC=-1529 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110000; // iC= -848 
// vC = 14'b1111100101000001; // vC=-1727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111001; // iC= -839 
// vC = 14'b1111100011001110; // vC=-1842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011001; // iC= -871 
// vC = 14'b1111100100010010; // vC=-1774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011010; // iC= -998 
// vC = 14'b1111100111011000; // vC=-1576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010100; // iC= -876 
// vC = 14'b1111100100100001; // vC=-1759 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b1111100011010010; // vC=-1838 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111001; // iC= -903 
// vC = 14'b1111100111110001; // vC=-1551 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100110; // iC= -794 
// vC = 14'b1111100101011100; // vC=-1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100011; // iC=-1053 
// vC = 14'b1111100010111000; // vC=-1864 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101010; // iC= -790 
// vC = 14'b1111100110011010; // vC=-1638 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001110; // iC= -946 
// vC = 14'b1111100111001100; // vC=-1588 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000101; // iC=-1019 
// vC = 14'b1111100011111100; // vC=-1796 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111110; // iC= -962 
// vC = 14'b1111100011101011; // vC=-1813 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101000; // iC= -984 
// vC = 14'b1111100010100011; // vC=-1885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010111; // iC= -809 
// vC = 14'b1111100110011000; // vC=-1640 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011001; // iC= -871 
// vC = 14'b1111100100101101; // vC=-1747 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000101; // iC= -763 
// vC = 14'b1111100100000110; // vC=-1786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100100; // iC= -732 
// vC = 14'b1111100011001110; // vC=-1842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110000; // iC= -912 
// vC = 14'b1111100101100001; // vC=-1695 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001011; // iC= -757 
// vC = 14'b1111100100101001; // vC=-1751 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101100; // iC= -724 
// vC = 14'b1111100101100010; // vC=-1694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111000; // iC= -776 
// vC = 14'b1111100011100011; // vC=-1821 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111000; // iC= -712 
// vC = 14'b1111100101100011; // vC=-1693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011000; // iC= -872 
// vC = 14'b1111100011001111; // vC=-1841 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111000; // iC= -648 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110111; // iC= -905 
// vC = 14'b1111100110101000; // vC=-1624 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101111; // iC= -913 
// vC = 14'b1111100100011000; // vC=-1768 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001001; // iC= -695 
// vC = 14'b1111100101111101; // vC=-1667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011001; // iC= -615 
// vC = 14'b1111100101010000; // vC=-1712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000000; // iC= -768 
// vC = 14'b1111100001110110; // vC=-1930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110101; // iC= -843 
// vC = 14'b1111100101110001; // vC=-1679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100001; // iC= -799 
// vC = 14'b1111100110010011; // vC=-1645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110100; // iC= -908 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111110; // iC= -770 
// vC = 14'b1111100010011111; // vC=-1889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101011; // iC= -853 
// vC = 14'b1111100001111111; // vC=-1921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010111; // iC= -681 
// vC = 14'b1111100010011100; // vC=-1892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010010; // iC= -878 
// vC = 14'b1111100101100010; // vC=-1694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001101; // iC= -755 
// vC = 14'b1111100001011001; // vC=-1959 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001000; // iC= -696 
// vC = 14'b1111100010001111; // vC=-1905 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000000; // iC= -832 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101001; // iC= -791 
// vC = 14'b1111100011101001; // vC=-1815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010001; // iC= -815 
// vC = 14'b1111100010110101; // vC=-1867 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011111; // iC= -545 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000001; // iC= -703 
// vC = 14'b1111100100010001; // vC=-1775 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011111; // iC= -609 
// vC = 14'b1111100100110111; // vC=-1737 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011010; // iC= -614 
// vC = 14'b1111100011001101; // vC=-1843 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100101; // iC= -795 
// vC = 14'b1111100101001010; // vC=-1718 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000000; // iC= -768 
// vC = 14'b1111100010111011; // vC=-1861 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111011; // iC= -645 
// vC = 14'b1111100011111010; // vC=-1798 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010000; // iC= -688 
// vC = 14'b1111100100111110; // vC=-1730 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011000; // iC= -808 
// vC = 14'b1111100001001000; // vC=-1976 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011011; // iC= -677 
// vC = 14'b1111100101010010; // vC=-1710 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100111; // iC= -473 
// vC = 14'b1111100001001111; // vC=-1969 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111010; // iC= -774 
// vC = 14'b1111100011011111; // vC=-1825 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011100; // iC= -612 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010000; // iC= -624 
// vC = 14'b1111100001011011; // vC=-1957 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110110; // iC= -458 
// vC = 14'b1111100001010100; // vC=-1964 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000100; // iC= -444 
// vC = 14'b1111100101011010; // vC=-1702 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011000; // iC= -488 
// vC = 14'b1111100010010111; // vC=-1897 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110001; // iC= -719 
// vC = 14'b1111100011010101; // vC=-1835 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000010; // iC= -446 
// vC = 14'b1111100011100110; // vC=-1818 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001110; // iC= -562 
// vC = 14'b1111100010110011; // vC=-1869 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001000; // iC= -568 
// vC = 14'b1111100000010011; // vC=-2029 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101001; // iC= -407 
// vC = 14'b1111100101000010; // vC=-1726 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010000; // iC= -432 
// vC = 14'b1111100000010011; // vC=-2029 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100000; // iC= -672 
// vC = 14'b1111100011100000; // vC=-1824 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001001; // iC= -439 
// vC = 14'b1111100001100000; // vC=-1952 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011100; // iC= -612 
// vC = 14'b1111100100111111; // vC=-1729 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010011; // iC= -429 
// vC = 14'b1111100100011101; // vC=-1763 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010101101; // iC= -339 
// vC = 14'b1111100100001110; // vC=-1778 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100111; // iC= -473 
// vC = 14'b1111100000101100; // vC=-2004 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111110; // iC= -386 
// vC = 14'b1111100010001111; // vC=-1905 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110110; // iC= -330 
// vC = 14'b1111011111111011; // vC=-2053 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011101; // iC= -291 
// vC = 14'b1111100001000111; // vC=-1977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001001; // iC= -567 
// vC = 14'b1111100010111111; // vC=-1857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111011; // iC= -389 
// vC = 14'b1111100001010010; // vC=-1966 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011101; // iC= -419 
// vC = 14'b1111100000110001; // vC=-1999 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000101; // iC= -251 
// vC = 14'b1111100100101110; // vC=-1746 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110010; // iC= -334 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011001; // iC= -423 
// vC = 14'b1111100001011001; // vC=-1959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110000; // iC= -464 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000110; // iC= -442 
// vC = 14'b1111100001100100; // vC=-1948 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000001; // iC= -383 
// vC = 14'b1111100000101000; // vC=-2008 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011010; // iC= -294 
// vC = 14'b1111100010000010; // vC=-1918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001100; // iC= -244 
// vC = 14'b1111100000110100; // vC=-1996 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001110; // iC= -114 
// vC = 14'b1111100011100010; // vC=-1822 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001011; // iC= -117 
// vC = 14'b1111100000111111; // vC=-1985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011100000; // iC= -288 
// vC = 14'b1111100001011010; // vC=-1958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011100; // iC= -292 
// vC = 14'b1111100011111100; // vC=-1796 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100110; // iC= -346 
// vC = 14'b1111100001011100; // vC=-1956 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000110; // iC= -314 
// vC = 14'b1111100001101111; // vC=-1937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001110; // iC=  -50 
// vC = 14'b1111100011101011; // vC=-1813 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101011011; // iC= -165 
// vC = 14'b1111100100001000; // vC=-1784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111111; // iC=  -65 
// vC = 14'b1111100011100000; // vC=-1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100100; // iC=   36 
// vC = 14'b1111100001000000; // vC=-1984 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100110; // iC=   38 
// vC = 14'b1111100011001010; // vC=-1846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000010; // iC= -190 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100000; // iC=  -32 
// vC = 14'b1111100100100000; // vC=-1760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000100; // iC= -124 
// vC = 14'b1111100001010001; // vC=-1967 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000111100; // iC=   60 
// vC = 14'b1111100011001001; // vC=-1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110001; // iC=  177 
// vC = 14'b1111011111101011; // vC=-2069 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011001; // iC= -103 
// vC = 14'b1111100100011010; // vC=-1766 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100000; // iC=  224 
// vC = 14'b1111100000101110; // vC=-2002 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100010; // iC=   98 
// vC = 14'b1111100001110011; // vC=-1933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101011; // iC=  171 
// vC = 14'b1111100000101000; // vC=-2008 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100101; // iC=   37 
// vC = 14'b1111100100000010; // vC=-1790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101000; // iC=  232 
// vC = 14'b1111100000110101; // vC=-1995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101100; // iC=  236 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111001; // iC=  313 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110110; // iC=  118 
// vC = 14'b1111100100010010; // vC=-1774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011011; // iC=  155 
// vC = 14'b1111100011111011; // vC=-1797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001010; // iC=  330 
// vC = 14'b1111100001010110; // vC=-1962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110010; // iC=  306 
// vC = 14'b1111100000101001; // vC=-2007 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010111; // iC=  343 
// vC = 14'b1111100010101011; // vC=-1877 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010101; // iC=  469 
// vC = 14'b1111100011101000; // vC=-1816 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001111; // iC=  399 
// vC = 14'b1111100100101101; // vC=-1747 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111111; // iC=  383 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000100; // iC=  324 
// vC = 14'b1111100010101010; // vC=-1878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010110; // iC=  342 
// vC = 14'b1111100011110100; // vC=-1804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100011; // iC=  611 
// vC = 14'b1111100001000101; // vC=-1979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111011; // iC=  379 
// vC = 14'b1111100001011001; // vC=-1959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001000; // iC=  456 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111010; // iC=  442 
// vC = 14'b1111100011111000; // vC=-1800 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110010; // iC=  626 
// vC = 14'b1111100010000000; // vC=-1920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101011; // iC=  683 
// vC = 14'b1111100011000001; // vC=-1855 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110111; // iC=  631 
// vC = 14'b1111100001000011; // vC=-1981 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010000; // iC=  592 
// vC = 14'b1111100001101000; // vC=-1944 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011110; // iC=  734 
// vC = 14'b1111100100001101; // vC=-1779 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100011; // iC=  547 
// vC = 14'b1111100100100110; // vC=-1754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101000; // iC=  552 
// vC = 14'b1111100000110110; // vC=-1994 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101011; // iC=  875 
// vC = 14'b1111100100010111; // vC=-1769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110010; // iC=  626 
// vC = 14'b1111100001011101; // vC=-1955 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001000; // iC=  712 
// vC = 14'b1111100101100111; // vC=-1689 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000011; // iC=  643 
// vC = 14'b1111100100101000; // vC=-1752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011000; // iC=  664 
// vC = 14'b1111100001101011; // vC=-1941 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010000; // iC=  720 
// vC = 14'b1111100101110110; // vC=-1674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010110; // iC=  918 
// vC = 14'b1111100011111000; // vC=-1800 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111001; // iC= 1017 
// vC = 14'b1111100100101100; // vC=-1748 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111001; // iC=  825 
// vC = 14'b1111100101011010; // vC=-1702 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101001; // iC= 1001 
// vC = 14'b1111100001100010; // vC=-1950 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000010; // iC= 1090 
// vC = 14'b1111100010010111; // vC=-1897 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101111; // iC=  815 
// vC = 14'b1111100110001100; // vC=-1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110110; // iC=  886 
// vC = 14'b1111100100101000; // vC=-1752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111111; // iC=  895 
// vC = 14'b1111100010000110; // vC=-1914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000000; // iC= 1024 
// vC = 14'b1111100100000010; // vC=-1790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101000; // iC=  936 
// vC = 14'b1111100101101100; // vC=-1684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100111; // iC=  935 
// vC = 14'b1111100010101000; // vC=-1880 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011100; // iC= 1116 
// vC = 14'b1111100101101011; // vC=-1685 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000001; // iC= 1025 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001110; // iC= 1102 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000010; // iC= 1218 
// vC = 14'b1111100010010001; // vC=-1903 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000000; // iC= 1216 
// vC = 14'b1111100100000010; // vC=-1790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110001; // iC= 1137 
// vC = 14'b1111100110101010; // vC=-1622 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011101; // iC= 1053 
// vC = 14'b1111100010111111; // vC=-1857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100100; // iC= 1124 
// vC = 14'b1111100010110011; // vC=-1869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011011; // iC= 1115 
// vC = 14'b1111100110010111; // vC=-1641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000100; // iC= 1412 
// vC = 14'b1111100110110001; // vC=-1615 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011010; // iC= 1114 
// vC = 14'b1111100110101111; // vC=-1617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001011; // iC= 1419 
// vC = 14'b1111100100010000; // vC=-1776 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001101; // iC= 1357 
// vC = 14'b1111100100001101; // vC=-1779 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101011; // iC= 1323 
// vC = 14'b1111100110001110; // vC=-1650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101110; // iC= 1454 
// vC = 14'b1111100101111111; // vC=-1665 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101100; // iC= 1324 
// vC = 14'b1111100111110110; // vC=-1546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100011; // iC= 1379 
// vC = 14'b1111100101100100; // vC=-1692 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101101; // iC= 1389 
// vC = 14'b1111100111011001; // vC=-1575 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101000; // iC= 1256 
// vC = 14'b1111100101000110; // vC=-1722 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101000; // iC= 1576 
// vC = 14'b1111100101111001; // vC=-1671 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010100; // iC= 1492 
// vC = 14'b1111100100011000; // vC=-1768 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010100; // iC= 1492 
// vC = 14'b1111100110011001; // vC=-1639 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101010; // iC= 1322 
// vC = 14'b1111100100001011; // vC=-1781 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100101; // iC= 1637 
// vC = 14'b1111100110001100; // vC=-1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001000; // iC= 1416 
// vC = 14'b1111100100010010; // vC=-1774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001101; // iC= 1421 
// vC = 14'b1111100111001010; // vC=-1590 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101011; // iC= 1579 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110000; // iC= 1584 
// vC = 14'b1111100110000101; // vC=-1659 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010101; // iC= 1493 
// vC = 14'b1111101001010111; // vC=-1449 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010110; // iC= 1558 
// vC = 14'b1111100111011110; // vC=-1570 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100000; // iC= 1440 
// vC = 14'b1111100101011011; // vC=-1701 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111001; // iC= 1657 
// vC = 14'b1111100111111110; // vC=-1538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110010; // iC= 1586 
// vC = 14'b1111100110100010; // vC=-1630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101000; // iC= 1512 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101010; // iC= 1578 
// vC = 14'b1111101001011011; // vC=-1445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101011; // iC= 1707 
// vC = 14'b1111101000000111; // vC=-1529 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100101; // iC= 1573 
// vC = 14'b1111100110000111; // vC=-1657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010110; // iC= 1750 
// vC = 14'b1111100110111101; // vC=-1603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110000; // iC= 1776 
// vC = 14'b1111101000001001; // vC=-1527 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010001; // iC= 1617 
// vC = 14'b1111101001010000; // vC=-1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101101; // iC= 1773 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011010; // iC= 1818 
// vC = 14'b1111100110101111; // vC=-1617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111101; // iC= 1789 
// vC = 14'b1111101010011100; // vC=-1380 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111110; // iC= 1598 
// vC = 14'b1111101010101110; // vC=-1362 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111011; // iC= 1659 
// vC = 14'b1111101001101001; // vC=-1431 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011111; // iC= 1631 
// vC = 14'b1111101010001011; // vC=-1397 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100111; // iC= 1895 
// vC = 14'b1111101001001101; // vC=-1459 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110000; // iC= 1712 
// vC = 14'b1111101000101110; // vC=-1490 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110000; // iC= 1712 
// vC = 14'b1111101000110100; // vC=-1484 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100010; // iC= 1698 
// vC = 14'b1111101010111110; // vC=-1346 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101001; // iC= 1833 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010101; // iC= 1749 
// vC = 14'b1111101001011001; // vC=-1447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011100; // iC= 1948 
// vC = 14'b1111101001100000; // vC=-1440 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010001; // iC= 1873 
// vC = 14'b1111101001001100; // vC=-1460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b1111101001111111; // vC=-1409 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101111; // iC= 1775 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111001; // iC= 1785 
// vC = 14'b1111101100100011; // vC=-1245 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b1111101010110011; // vC=-1357 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b1111101011101100; // vC=-1300 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000100; // iC= 1924 
// vC = 14'b1111101000101001; // vC=-1495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101110; // iC= 1838 
// vC = 14'b1111101011001110; // vC=-1330 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001100; // iC= 1740 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000101; // iC= 1861 
// vC = 14'b1111101010001011; // vC=-1397 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b1111101100011010; // vC=-1254 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111101011010110; // vC=-1322 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b1111101101000010; // vC=-1214 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000010; // iC= 1794 
// vC = 14'b1111101100101101; // vC=-1235 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100110; // iC= 1830 
// vC = 14'b1111101101000101; // vC=-1211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001101; // iC= 1869 
// vC = 14'b1111101001101011; // vC=-1429 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101110; // iC= 1966 
// vC = 14'b1111101110011101; // vC=-1123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110001; // iC= 1969 
// vC = 14'b1111101010101000; // vC=-1368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111100; // iC= 1852 
// vC = 14'b1111101110000011; // vC=-1149 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011100; // iC= 2012 
// vC = 14'b1111101110001001; // vC=-1143 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100011; // iC= 1891 
// vC = 14'b1111101011011001; // vC=-1319 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110110; // iC= 2038 
// vC = 14'b1111101101101010; // vC=-1174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010111; // iC= 1879 
// vC = 14'b1111101100000111; // vC=-1273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b1111101110101011; // vC=-1109 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010001; // iC= 1873 
// vC = 14'b1111101101101111; // vC=-1169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000000; // iC= 2048 
// vC = 14'b1111101011110100; // vC=-1292 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b1111101110110011; // vC=-1101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001100; // iC= 1868 
// vC = 14'b1111101100101000; // vC=-1240 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110110; // iC= 1974 
// vC = 14'b1111101101011110; // vC=-1186 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b1111110000001110; // vC=-1010 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111111; // iC= 1855 
// vC = 14'b1111110000010101; // vC=-1003 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b1111101011110111; // vC=-1289 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b1111101101100110; // vC=-1178 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110000; // iC= 1904 
// vC = 14'b1111101101101011; // vC=-1173 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111100; // iC= 1852 
// vC = 14'b1111101111001010; // vC=-1078 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010110; // iC= 1878 
// vC = 14'b1111101100111010; // vC=-1222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b1111101111001110; // vC=-1074 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111100; // iC= 2108 
// vC = 14'b1111101110110011; // vC=-1101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100101; // iC= 1957 
// vC = 14'b1111110000111110; // vC= -962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b1111101110001101; // vC=-1139 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100111; // iC= 2087 
// vC = 14'b1111101111001110; // vC=-1074 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011011; // iC= 2139 
// vC = 14'b1111101111100010; // vC=-1054 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100010; // iC= 2018 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b1111110001011011; // vC= -933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000010; // iC= 2114 
// vC = 14'b1111101111100100; // vC=-1052 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110001; // iC= 1841 
// vC = 14'b1111101111111011; // vC=-1029 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010011; // iC= 2067 
// vC = 14'b1111101110110110; // vC=-1098 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b1111110000111101; // vC= -963 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111100; // iC= 1852 
// vC = 14'b1111110001010011; // vC= -941 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101101; // iC= 2029 
// vC = 14'b1111110010010110; // vC= -874 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000010; // iC= 1858 
// vC = 14'b1111110001011101; // vC= -931 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b1111101110110010; // vC=-1102 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110110; // iC= 1974 
// vC = 14'b1111110000111110; // vC= -962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b1111110000010011; // vC=-1005 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010000; // iC= 2064 
// vC = 14'b1111101111010000; // vC=-1072 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011000; // iC= 2136 
// vC = 14'b1111110001110001; // vC= -911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001001; // iC= 1993 
// vC = 14'b1111101111110101; // vC=-1035 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b1111101111100111; // vC=-1049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110000; // iC= 1840 
// vC = 14'b1111101111011101; // vC=-1059 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110011; // iC= 1971 
// vC = 14'b1111110010111101; // vC= -835 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b1111110011100101; // vC= -795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000110; // iC= 2118 
// vC = 14'b1111110011000100; // vC= -828 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010001; // iC= 2129 
// vC = 14'b1111110001100001; // vC= -927 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010010; // iC= 1874 
// vC = 14'b1111110011100010; // vC= -798 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010010; // iC= 2002 
// vC = 14'b1111110000101101; // vC= -979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000010; // iC= 1922 
// vC = 14'b1111110100010011; // vC= -749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b1111110001101000; // vC= -920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100110; // iC= 2086 
// vC = 14'b1111110010000101; // vC= -891 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b1111110101010100; // vC= -684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b1111110001010101; // vC= -939 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110100; // iC= 2100 
// vC = 14'b1111110010100000; // vC= -864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b1111110101110110; // vC= -650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000010; // iC= 1858 
// vC = 14'b1111110001110010; // vC= -910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111110110000010; // vC= -638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b1111110100001000; // vC= -760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001011; // iC= 1867 
// vC = 14'b1111110100010011; // vC= -749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000000; // iC= 1856 
// vC = 14'b1111110001101000; // vC= -920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101011; // iC= 1963 
// vC = 14'b1111110100101010; // vC= -726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b1111110001111110; // vC= -898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100010; // iC= 2018 
// vC = 14'b1111110100010100; // vC= -748 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b1111110110110001; // vC= -591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000100; // iC= 1988 
// vC = 14'b1111110111011000; // vC= -552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110101; // iC= 1845 
// vC = 14'b1111110111001010; // vC= -566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100001; // iC= 2017 
// vC = 14'b1111110101111010; // vC= -646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110000; // iC= 2096 
// vC = 14'b1111110111001100; // vC= -564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b1111110010111110; // vC= -834 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b1111110110111101; // vC= -579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100111; // iC= 2087 
// vC = 14'b1111110101001111; // vC= -689 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100110; // iC= 1830 
// vC = 14'b1111111000010001; // vC= -495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b1111110110010000; // vC= -624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101000; // iC= 2152 
// vC = 14'b1111110110011101; // vC= -611 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101001; // iC= 1833 
// vC = 14'b1111110111010000; // vC= -560 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b1111110100011111; // vC= -737 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111110; // iC= 1918 
// vC = 14'b1111110110010101; // vC= -619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100111; // iC= 1831 
// vC = 14'b1111110101011011; // vC= -677 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101110; // iC= 2094 
// vC = 14'b1111110110011001; // vC= -615 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010010; // iC= 2002 
// vC = 14'b1111110110111100; // vC= -580 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100001; // iC= 1825 
// vC = 14'b1111111000001111; // vC= -497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111001; // iC= 2105 
// vC = 14'b1111110101111011; // vC= -645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011110; // iC= 2014 
// vC = 14'b1111111001010001; // vC= -431 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b1111110111100110; // vC= -538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100001; // iC= 2017 
// vC = 14'b1111111000111101; // vC= -451 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100000; // iC= 1888 
// vC = 14'b1111111010001100; // vC= -372 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111101; // iC= 2045 
// vC = 14'b1111110111010110; // vC= -554 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100100; // iC= 2020 
// vC = 14'b1111110110011001; // vC= -615 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110001; // iC= 2033 
// vC = 14'b1111110110001011; // vC= -629 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111000; // iC= 1848 
// vC = 14'b1111111001100010; // vC= -414 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101010; // iC= 2090 
// vC = 14'b1111111000000010; // vC= -510 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110010; // iC= 1842 
// vC = 14'b1111111000011101; // vC= -483 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100111; // iC= 2023 
// vC = 14'b1111111001001110; // vC= -434 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110011; // iC= 1971 
// vC = 14'b1111110110111100; // vC= -580 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001110; // iC= 2126 
// vC = 14'b1111111000110100; // vC= -460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101010; // iC= 1898 
// vC = 14'b1111111011010010; // vC= -302 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111111001000001; // vC= -447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b1111111010110000; // vC= -336 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000001; // iC= 1921 
// vC = 14'b1111111011000110; // vC= -314 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000110; // iC= 2118 
// vC = 14'b1111111001100101; // vC= -411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b1111111000011001; // vC= -487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000011; // iC= 2051 
// vC = 14'b1111111000101110; // vC= -466 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101111; // iC= 1839 
// vC = 14'b1111111001001100; // vC= -436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b1111111010111110; // vC= -322 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111101; // iC= 2109 
// vC = 14'b1111111001010000; // vC= -432 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010010; // iC= 1874 
// vC = 14'b1111111100010100; // vC= -236 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010100; // iC= 1876 
// vC = 14'b1111111011110111; // vC= -265 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000101; // iC= 1989 
// vC = 14'b1111111011100100; // vC= -284 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b1111111101010000; // vC= -176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b1111111001100101; // vC= -411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111111011101111; // vC= -273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110001; // iC= 2097 
// vC = 14'b1111111001110111; // vC= -393 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b1111111001110010; // vC= -398 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b1111111101101111; // vC= -145 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000000; // iC= 1984 
// vC = 14'b1111111101110011; // vC= -141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000111; // iC= 1799 
// vC = 14'b1111111100110011; // vC= -205 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b1111111011001100; // vC= -308 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111111011110011; // vC= -269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111111110000011; // vC= -125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b1111111101010101; // vC= -171 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000110; // iC= 1862 
// vC = 14'b1111111101011000; // vC= -168 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000000; // iC= 1920 
// vC = 14'b1111111101000001; // vC= -191 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001001; // iC= 1865 
// vC = 14'b1111111110110001; // vC=  -79 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111111010010111; // vC= -361 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110111; // iC= 1783 
// vC = 14'b1111111101111000; // vC= -136 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010010; // iC= 1874 
// vC = 14'b1111111110111111; // vC=  -65 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b1111111101101011; // vC= -149 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101111; // iC= 1839 
// vC = 14'b1111111111101100; // vC=  -20 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111111110111000; // vC=  -72 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011100; // iC= 1948 
// vC = 14'b1111111101110000; // vC= -144 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b1111111110100101; // vC=  -91 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001110; // iC= 1934 
// vC = 14'b1111111111011101; // vC=  -35 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011110; // iC= 2014 
// vC = 14'b1111111110111101; // vC=  -67 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010001; // iC= 1809 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001001; // iC= 2057 
// vC = 14'b0000000000000100; // vC=    4 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001001; // iC= 1865 
// vC = 14'b1111111101001011; // vC= -181 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010111; // iC= 1815 
// vC = 14'b1111111100110010; // vC= -206 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010010; // iC= 2066 
// vC = 14'b1111111100010111; // vC= -233 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111111100011000; // vC= -232 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000010; // iC= 1986 
// vC = 14'b0000000000000111; // vC=    7 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001000; // iC= 1800 
// vC = 14'b1111111110110100; // vC=  -76 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000000; // iC= 1792 
// vC = 14'b0000000000001111; // vC=   15 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b0000000000111111; // vC=   63 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000101; // iC= 1989 
// vC = 14'b1111111101111110; // vC= -130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101010; // iC= 1834 
// vC = 14'b0000000000010110; // vC=   22 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b1111111101011001; // vC= -167 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111000; // iC= 1784 
// vC = 14'b1111111110001010; // vC= -118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000100; // iC= 1924 
// vC = 14'b1111111101111010; // vC= -134 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b1111111101101110; // vC= -146 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001000; // iC= 1800 
// vC = 14'b0000000000011001; // vC=   25 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b1111111110000010; // vC= -126 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010010; // iC= 1746 
// vC = 14'b0000000001011010; // vC=   90 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111111111000100; // vC=  -60 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110000; // iC= 1904 
// vC = 14'b0000000001100010; // vC=   98 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001101; // iC= 1869 
// vC = 14'b0000000010010101; // vC=  149 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100000; // iC= 1824 
// vC = 14'b0000000000100101; // vC=   37 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011100; // iC= 1884 
// vC = 14'b0000000001010101; // vC=   85 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b0000000000011001; // vC=   25 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000011; // iC= 1859 
// vC = 14'b0000000000001000; // vC=    8 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b1111111111010000; // vC=  -48 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010101; // iC= 1749 
// vC = 14'b0000000010000000; // vC=  128 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101110; // iC= 1774 
// vC = 14'b0000000010000101; // vC=  133 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111000; // iC= 1720 
// vC = 14'b0000000010001111; // vC=  143 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100011; // iC= 1891 
// vC = 14'b0000000010000001; // vC=  129 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110100; // iC= 1844 
// vC = 14'b0000000000010111; // vC=   23 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100001; // iC= 1825 
// vC = 14'b0000000100011110; // vC=  286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011111; // iC= 1887 
// vC = 14'b1111111111101111; // vC=  -17 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101001; // iC= 1705 
// vC = 14'b0000000100111001; // vC=  313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101111; // iC= 1967 
// vC = 14'b0000000000101011; // vC=   43 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110101; // iC= 1845 
// vC = 14'b0000000010000100; // vC=  132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000000; // iC= 1984 
// vC = 14'b0000000100001101; // vC=  269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100101; // iC= 1957 
// vC = 14'b0000000011010011; // vC=  211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001101; // iC= 1677 
// vC = 14'b0000000010001110; // vC=  142 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111010; // iC= 1978 
// vC = 14'b0000000001110100; // vC=  116 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011011; // iC= 1691 
// vC = 14'b0000000010000010; // vC=  130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110100; // iC= 1716 
// vC = 14'b0000000011001110; // vC=  206 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011110; // iC= 1758 
// vC = 14'b0000000011001110; // vC=  206 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000100; // iC= 1732 
// vC = 14'b0000000110001110; // vC=  398 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b0000000101101000; // vC=  360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000100; // iC= 1796 
// vC = 14'b0000000100010010; // vC=  274 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000000; // iC= 1664 
// vC = 14'b0000000101111111; // vC=  383 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001100; // iC= 1804 
// vC = 14'b0000000010101000; // vC=  168 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111011; // iC= 1659 
// vC = 14'b0000000101101101; // vC=  365 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100111; // iC= 1831 
// vC = 14'b0000000110010010; // vC=  402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b0000000100001100; // vC=  268 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000011; // iC= 1923 
// vC = 14'b0000000100110111; // vC=  311 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011101; // iC= 1821 
// vC = 14'b0000000110100010; // vC=  418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010001; // iC= 1681 
// vC = 14'b0000000101000000; // vC=  320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001111; // iC= 1807 
// vC = 14'b0000000010101101; // vC=  173 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b0000000100100010; // vC=  290 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011000; // iC= 1816 
// vC = 14'b0000000111110001; // vC=  497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001111; // iC= 1871 
// vC = 14'b0000000100111001; // vC=  313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b0000000101010011; // vC=  339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111000; // iC= 1848 
// vC = 14'b0000000101000100; // vC=  324 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b0000000011100000; // vC=  224 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110000; // iC= 1904 
// vC = 14'b0000000110011011; // vC=  411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110001; // iC= 1841 
// vC = 14'b0000000110111101; // vC=  445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001101; // iC= 1741 
// vC = 14'b0000000100111010; // vC=  314 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b0000000111111111; // vC=  511 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011010; // iC= 1626 
// vC = 14'b0000000110101101; // vC=  429 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b0000000110010111; // vC=  407 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100101; // iC= 1765 
// vC = 14'b0000000111000101; // vC=  453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100011; // iC= 1699 
// vC = 14'b0000000110101010; // vC=  426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001111; // iC= 1743 
// vC = 14'b0000001000101110; // vC=  558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010100; // iC= 1684 
// vC = 14'b0000001000000011; // vC=  515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100100; // iC= 1572 
// vC = 14'b0000000110100100; // vC=  420 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011110; // iC= 1630 
// vC = 14'b0000000101001011; // vC=  331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010001; // iC= 1873 
// vC = 14'b0000000101110110; // vC=  374 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000001; // iC= 1729 
// vC = 14'b0000000110010010; // vC=  402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011101; // iC= 1693 
// vC = 14'b0000001001000001; // vC=  577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000001; // iC= 1665 
// vC = 14'b0000000111110100; // vC=  500 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011100; // iC= 1628 
// vC = 14'b0000000101001101; // vC=  333 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100101; // iC= 1637 
// vC = 14'b0000000111011111; // vC=  479 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111010; // iC= 1786 
// vC = 14'b0000000111011011; // vC=  475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000000; // iC= 1600 
// vC = 14'b0000000110001011; // vC=  395 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010000; // iC= 1808 
// vC = 14'b0000001000110110; // vC=  566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001101; // iC= 1677 
// vC = 14'b0000000110011010; // vC=  410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110111; // iC= 1719 
// vC = 14'b0000001001010001; // vC=  593 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100011; // iC= 1763 
// vC = 14'b0000000111010010; // vC=  466 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001011; // iC= 1739 
// vC = 14'b0000001000110100; // vC=  564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101000; // iC= 1640 
// vC = 14'b0000000111100111; // vC=  487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000010; // iC= 1794 
// vC = 14'b0000001000001001; // vC=  521 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000111; // iC= 1607 
// vC = 14'b0000000111100011; // vC=  483 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111011; // iC= 1659 
// vC = 14'b0000000110110111; // vC=  439 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000100; // iC= 1540 
// vC = 14'b0000001000001011; // vC=  523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011110; // iC= 1502 
// vC = 14'b0000001000111100; // vC=  572 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010110; // iC= 1750 
// vC = 14'b0000001001101011; // vC=  619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111100; // iC= 1660 
// vC = 14'b0000001000011110; // vC=  542 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000010; // iC= 1730 
// vC = 14'b0000000111011011; // vC=  475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010110; // iC= 1750 
// vC = 14'b0000001001011010; // vC=  602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001011; // iC= 1547 
// vC = 14'b0000001001110001; // vC=  625 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100001; // iC= 1697 
// vC = 14'b0000001010110100; // vC=  692 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010011; // iC= 1491 
// vC = 14'b0000001001010100; // vC=  596 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011100; // iC= 1564 
// vC = 14'b0000001010000101; // vC=  645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110110; // iC= 1718 
// vC = 14'b0000001011010110; // vC=  726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111100; // iC= 1468 
// vC = 14'b0000001010001000; // vC=  648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101100; // iC= 1516 
// vC = 14'b0000001100111011; // vC=  827 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101100; // iC= 1708 
// vC = 14'b0000001011101000; // vC=  744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110101; // iC= 1589 
// vC = 14'b0000001011011101; // vC=  733 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100100; // iC= 1572 
// vC = 14'b0000001100100001; // vC=  801 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010101; // iC= 1621 
// vC = 14'b0000001010101100; // vC=  684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101111; // iC= 1583 
// vC = 14'b0000001101010101; // vC=  853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000000; // iC= 1472 
// vC = 14'b0000001011010000; // vC=  720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001100; // iC= 1740 
// vC = 14'b0000001010100010; // vC=  674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000001; // iC= 1729 
// vC = 14'b0000001001100100; // vC=  612 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110000; // iC= 1520 
// vC = 14'b0000001011001010; // vC=  714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001001; // iC= 1481 
// vC = 14'b0000001100001110; // vC=  782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101000; // iC= 1448 
// vC = 14'b0000001101111000; // vC=  888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011011; // iC= 1691 
// vC = 14'b0000001010011010; // vC=  666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010111; // iC= 1559 
// vC = 14'b0000001011010110; // vC=  726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100111; // iC= 1639 
// vC = 14'b0000001100011101; // vC=  797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000111; // iC= 1415 
// vC = 14'b0000001110001111; // vC=  911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001101; // iC= 1421 
// vC = 14'b0000001011010000; // vC=  720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100010; // iC= 1506 
// vC = 14'b0000001110000111; // vC=  903 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100010; // iC= 1634 
// vC = 14'b0000001011001110; // vC=  718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101100; // iC= 1580 
// vC = 14'b0000001011100111; // vC=  743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111001; // iC= 1593 
// vC = 14'b0000001100001100; // vC=  780 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101111; // iC= 1391 
// vC = 14'b0000001011010111; // vC=  727 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011110; // iC= 1566 
// vC = 14'b0000001110000110; // vC=  902 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110000; // iC= 1456 
// vC = 14'b0000001011001101; // vC=  717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000001; // iC= 1409 
// vC = 14'b0000001101111110; // vC=  894 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101101; // iC= 1517 
// vC = 14'b0000001100111011; // vC=  827 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100011; // iC= 1443 
// vC = 14'b0000001110010000; // vC=  912 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100001; // iC= 1569 
// vC = 14'b0000001010110111; // vC=  695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001011; // iC= 1611 
// vC = 14'b0000001011010111; // vC=  727 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011110; // iC= 1438 
// vC = 14'b0000001011001101; // vC=  717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011010; // iC= 1562 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101111; // iC= 1583 
// vC = 14'b0000001011101000; // vC=  744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111000; // iC= 1528 
// vC = 14'b0000001101001101; // vC=  845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001100; // iC= 1356 
// vC = 14'b0000001100010011; // vC=  787 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101000; // iC= 1512 
// vC = 14'b0000010000010001; // vC= 1041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011011; // iC= 1499 
// vC = 14'b0000001101101110; // vC=  878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100100; // iC= 1316 
// vC = 14'b0000001111000000; // vC=  960 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111000; // iC= 1592 
// vC = 14'b0000001100100010; // vC=  802 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111111; // iC= 1599 
// vC = 14'b0000010000110001; // vC= 1073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010110; // iC= 1558 
// vC = 14'b0000001110100001; // vC=  929 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111111; // iC= 1343 
// vC = 14'b0000001110100111; // vC=  935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110000; // iC= 1328 
// vC = 14'b0000001101010100; // vC=  852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000100; // iC= 1412 
// vC = 14'b0000001110101101; // vC=  941 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101010; // iC= 1514 
// vC = 14'b0000001100101110; // vC=  814 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011011; // iC= 1563 
// vC = 14'b0000001111001111; // vC=  975 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100001; // iC= 1313 
// vC = 14'b0000001100011111; // vC=  799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101100; // iC= 1388 
// vC = 14'b0000001101001010; // vC=  842 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011101; // iC= 1501 
// vC = 14'b0000010000000000; // vC= 1024 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011000; // iC= 1368 
// vC = 14'b0000001110001001; // vC=  905 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101110; // iC= 1326 
// vC = 14'b0000001111110001; // vC= 1009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100111; // iC= 1511 
// vC = 14'b0000010001100111; // vC= 1127 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101011; // iC= 1323 
// vC = 14'b0000010000001000; // vC= 1032 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000001; // iC= 1473 
// vC = 14'b0000001110001010; // vC=  906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100011; // iC= 1443 
// vC = 14'b0000001110100010; // vC=  930 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011110; // iC= 1502 
// vC = 14'b0000001111111010; // vC= 1018 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111000; // iC= 1336 
// vC = 14'b0000010001011000; // vC= 1112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001111; // iC= 1231 
// vC = 14'b0000010010100001; // vC= 1185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101111; // iC= 1327 
// vC = 14'b0000010001001010; // vC= 1098 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010111; // iC= 1431 
// vC = 14'b0000010010011101; // vC= 1181 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010011; // iC= 1491 
// vC = 14'b0000001111101111; // vC= 1007 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100000; // iC= 1440 
// vC = 14'b0000010010110111; // vC= 1207 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011101; // iC= 1373 
// vC = 14'b0000001111100011; // vC=  995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010001; // iC= 1233 
// vC = 14'b0000010011000110; // vC= 1222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010111; // iC= 1303 
// vC = 14'b0000010001101011; // vC= 1131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000001; // iC= 1345 
// vC = 14'b0000010001000011; // vC= 1091 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110101; // iC= 1461 
// vC = 14'b0000010001000110; // vC= 1094 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111010; // iC= 1402 
// vC = 14'b0000001111111001; // vC= 1017 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111010; // iC= 1402 
// vC = 14'b0000010001101010; // vC= 1130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001111; // iC= 1423 
// vC = 14'b0000001110101001; // vC=  937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011110; // iC= 1310 
// vC = 14'b0000010001010011; // vC= 1107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110111; // iC= 1399 
// vC = 14'b0000010010001010; // vC= 1162 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110000; // iC= 1264 
// vC = 14'b0000001111110011; // vC= 1011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111001; // iC= 1145 
// vC = 14'b0000010001001000; // vC= 1096 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001110; // iC= 1230 
// vC = 14'b0000001111000001; // vC=  961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001101; // iC= 1229 
// vC = 14'b0000001111100010; // vC=  994 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000010; // iC= 1410 
// vC = 14'b0000010010110110; // vC= 1206 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011001; // iC= 1305 
// vC = 14'b0000010010000001; // vC= 1153 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110101; // iC= 1205 
// vC = 14'b0000010001100011; // vC= 1123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101111; // iC= 1327 
// vC = 14'b0000010001110110; // vC= 1142 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100111; // iC= 1127 
// vC = 14'b0000010010011000; // vC= 1176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110011; // iC= 1395 
// vC = 14'b0000010011111011; // vC= 1275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000000; // iC= 1280 
// vC = 14'b0000010000010001; // vC= 1041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010111; // iC= 1303 
// vC = 14'b0000010100000110; // vC= 1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010000; // iC= 1104 
// vC = 14'b0000010010111110; // vC= 1214 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001010; // iC= 1098 
// vC = 14'b0000010010000000; // vC= 1152 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101001; // iC= 1385 
// vC = 14'b0000010010010110; // vC= 1174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100100; // iC= 1124 
// vC = 14'b0000010001101110; // vC= 1134 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100100; // iC= 1316 
// vC = 14'b0000010000010110; // vC= 1046 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100111; // iC= 1191 
// vC = 14'b0000010010111010; // vC= 1210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010011; // iC= 1363 
// vC = 14'b0000010001111001; // vC= 1145 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110111; // iC= 1079 
// vC = 14'b0000010001010111; // vC= 1111 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010001; // iC= 1105 
// vC = 14'b0000010011011000; // vC= 1240 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101011; // iC= 1131 
// vC = 14'b0000010010011110; // vC= 1182 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011010; // iC= 1178 
// vC = 14'b0000010101000110; // vC= 1350 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001001; // iC= 1033 
// vC = 14'b0000010011110000; // vC= 1264 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101110; // iC= 1134 
// vC = 14'b0000010010000111; // vC= 1159 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110111; // iC= 1271 
// vC = 14'b0000010001010011; // vC= 1107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000110; // iC= 1030 
// vC = 14'b0000010001001001; // vC= 1097 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110100; // iC= 1140 
// vC = 14'b0000010001010001; // vC= 1105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011110; // iC= 1310 
// vC = 14'b0000010011111100; // vC= 1276 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000110; // iC= 1094 
// vC = 14'b0000010100110100; // vC= 1332 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101001; // iC= 1257 
// vC = 14'b0000010011110110; // vC= 1270 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100000; // iC= 1056 
// vC = 14'b0000010100001111; // vC= 1295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110110; // iC= 1014 
// vC = 14'b0000010110011011; // vC= 1435 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101001; // iC= 1193 
// vC = 14'b0000010010010010; // vC= 1170 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000100; // iC= 1220 
// vC = 14'b0000010100111011; // vC= 1339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011110; // iC= 1118 
// vC = 14'b0000010110000110; // vC= 1414 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010010; // iC= 1170 
// vC = 14'b0000010011101100; // vC= 1260 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101100; // iC= 1132 
// vC = 14'b0000010100001011; // vC= 1291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101111; // iC= 1007 
// vC = 14'b0000010100011010; // vC= 1306 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011101; // iC=  989 
// vC = 14'b0000010110110000; // vC= 1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111110; // iC= 1086 
// vC = 14'b0000010010011110; // vC= 1182 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101000; // iC= 1064 
// vC = 14'b0000010101100110; // vC= 1382 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000011; // iC= 1091 
// vC = 14'b0000010101111100; // vC= 1404 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000111; // iC= 1031 
// vC = 14'b0000010011000100; // vC= 1220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100101; // iC= 1189 
// vC = 14'b0000010011100001; // vC= 1249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010100; // iC=  916 
// vC = 14'b0000010110000110; // vC= 1414 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111010; // iC= 1146 
// vC = 14'b0000010011111011; // vC= 1275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100000; // iC= 1184 
// vC = 14'b0000010101011000; // vC= 1368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001110; // iC= 1038 
// vC = 14'b0000010101001000; // vC= 1352 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001001; // iC= 1161 
// vC = 14'b0000010100000011; // vC= 1283 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011111; // iC=  927 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010010; // iC= 1042 
// vC = 14'b0000010110001000; // vC= 1416 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011100; // iC=  988 
// vC = 14'b0000010101101001; // vC= 1385 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001011; // iC= 1035 
// vC = 14'b0000010101101011; // vC= 1387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101010; // iC=  938 
// vC = 14'b0000010110101101; // vC= 1453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010001; // iC= 1041 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111111; // iC= 1023 
// vC = 14'b0000010100001000; // vC= 1288 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110000; // iC= 1008 
// vC = 14'b0000010110000111; // vC= 1415 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111101; // iC= 1085 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101101; // iC= 1133 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111101; // iC= 1149 
// vC = 14'b0000010011110000; // vC= 1264 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010001; // iC=  913 
// vC = 14'b0000010111110011; // vC= 1523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001001; // iC= 1097 
// vC = 14'b0000010110111111; // vC= 1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010110; // iC=  982 
// vC = 14'b0000010101111010; // vC= 1402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000011; // iC= 1091 
// vC = 14'b0000010100011010; // vC= 1306 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001100; // iC=  844 
// vC = 14'b0000010100000101; // vC= 1285 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011110; // iC=  990 
// vC = 14'b0000011000101001; // vC= 1577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010010; // iC=  914 
// vC = 14'b0000010110001010; // vC= 1418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010001; // iC= 1105 
// vC = 14'b0000010110010111; // vC= 1431 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100101; // iC=  805 
// vC = 14'b0000010101100101; // vC= 1381 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100100; // iC=  868 
// vC = 14'b0000010111001110; // vC= 1486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001000; // iC= 1096 
// vC = 14'b0000010100111111; // vC= 1343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010000; // iC=  912 
// vC = 14'b0000010100100010; // vC= 1314 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111110; // iC= 1022 
// vC = 14'b0000011000000010; // vC= 1538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b0000010110111101; // vC= 1469 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010000; // iC=  912 
// vC = 14'b0000011000011010; // vC= 1562 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111010; // iC=  890 
// vC = 14'b0000011000001100; // vC= 1548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001101; // iC=  845 
// vC = 14'b0000011001001101; // vC= 1613 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001000; // iC= 1032 
// vC = 14'b0000010111000101; // vC= 1477 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001101; // iC=  845 
// vC = 14'b0000010101101010; // vC= 1386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101011; // iC=  747 
// vC = 14'b0000010101000100; // vC= 1348 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101010; // iC=  810 
// vC = 14'b0000010110001101; // vC= 1421 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110001; // iC= 1009 
// vC = 14'b0000011001001000; // vC= 1608 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101101; // iC=  813 
// vC = 14'b0000011001000011; // vC= 1603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100111; // iC=  935 
// vC = 14'b0000010111001011; // vC= 1483 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000110; // iC=  902 
// vC = 14'b0000010111110100; // vC= 1524 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111110; // iC=  766 
// vC = 14'b0000010110010100; // vC= 1428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001001; // iC=  905 
// vC = 14'b0000010110011110; // vC= 1438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110100; // iC=  820 
// vC = 14'b0000011001000000; // vC= 1600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b0000010101111111; // vC= 1407 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011010; // iC=  730 
// vC = 14'b0000011001001101; // vC= 1613 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100101; // iC=  933 
// vC = 14'b0000010110010001; // vC= 1425 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110011; // iC=  947 
// vC = 14'b0000010101110000; // vC= 1392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000111; // iC=  711 
// vC = 14'b0000010111011001; // vC= 1497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111000; // iC=  696 
// vC = 14'b0000011000000011; // vC= 1539 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100110; // iC=  806 
// vC = 14'b0000011000000100; // vC= 1540 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101001; // iC=  745 
// vC = 14'b0000010101110011; // vC= 1395 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110111; // iC=  887 
// vC = 14'b0000010101010101; // vC= 1365 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011111; // iC=  863 
// vC = 14'b0000010110111110; // vC= 1470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100110; // iC=  806 
// vC = 14'b0000010111001001; // vC= 1481 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101011; // iC=  747 
// vC = 14'b0000011001110001; // vC= 1649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010110; // iC=  790 
// vC = 14'b0000011000111000; // vC= 1592 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011110; // iC=  734 
// vC = 14'b0000010111110010; // vC= 1522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011001; // iC=  857 
// vC = 14'b0000011001010101; // vC= 1621 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100110; // iC=  742 
// vC = 14'b0000010101101111; // vC= 1391 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110011; // iC=  755 
// vC = 14'b0000011010100010; // vC= 1698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111000; // iC=  568 
// vC = 14'b0000010101101110; // vC= 1390 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100010; // iC=  738 
// vC = 14'b0000010110011010; // vC= 1434 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100000; // iC=  800 
// vC = 14'b0000010110001001; // vC= 1417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100101; // iC=  677 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001111; // iC=  719 
// vC = 14'b0000010110001011; // vC= 1419 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100000; // iC=  608 
// vC = 14'b0000011001100101; // vC= 1637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000111; // iC=  839 
// vC = 14'b0000010110110111; // vC= 1463 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100100; // iC=  740 
// vC = 14'b0000010111111110; // vC= 1534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111000; // iC=  760 
// vC = 14'b0000011000000000; // vC= 1536 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010001; // iC=  721 
// vC = 14'b0000011001110111; // vC= 1655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001010; // iC=  714 
// vC = 14'b0000010110010010; // vC= 1426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110100; // iC=  756 
// vC = 14'b0000010111110010; // vC= 1522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001000; // iC=  520 
// vC = 14'b0000010110010100; // vC= 1428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110011; // iC=  627 
// vC = 14'b0000011010000110; // vC= 1670 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100101; // iC=  549 
// vC = 14'b0000011000100100; // vC= 1572 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100011; // iC=  611 
// vC = 14'b0000010110010110; // vC= 1430 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100101; // iC=  485 
// vC = 14'b0000011010100101; // vC= 1701 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100000; // iC=  544 
// vC = 14'b0000011001001101; // vC= 1613 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010000; // iC=  784 
// vC = 14'b0000011001001001; // vC= 1609 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101111; // iC=  495 
// vC = 14'b0000010110100001; // vC= 1441 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100101; // iC=  549 
// vC = 14'b0000011000101101; // vC= 1581 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110001; // iC=  689 
// vC = 14'b0000010111001110; // vC= 1486 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100010; // iC=  738 
// vC = 14'b0000011010011001; // vC= 1689 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011010; // iC=  602 
// vC = 14'b0000011000000100; // vC= 1540 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000100; // iC=  708 
// vC = 14'b0000011000111001; // vC= 1593 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000000; // iC=  704 
// vC = 14'b0000011010111101; // vC= 1725 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011101; // iC=  733 
// vC = 14'b0000011001101001; // vC= 1641 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010100; // iC=  596 
// vC = 14'b0000011001111110; // vC= 1662 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000101; // iC=  581 
// vC = 14'b0000011001011101; // vC= 1629 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001010; // iC=  586 
// vC = 14'b0000010111110010; // vC= 1522 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110101; // iC=  437 
// vC = 14'b0000011001001000; // vC= 1608 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000011; // iC=  579 
// vC = 14'b0000011010011111; // vC= 1695 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111010; // iC=  634 
// vC = 14'b0000011010100100; // vC= 1700 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010011; // iC=  467 
// vC = 14'b0000011100000100; // vC= 1796 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001001; // iC=  393 
// vC = 14'b0000011010001000; // vC= 1672 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000111; // iC=  391 
// vC = 14'b0000010111010011; // vC= 1491 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101110; // iC=  494 
// vC = 14'b0000011000111111; // vC= 1599 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010001; // iC=  593 
// vC = 14'b0000011011111001; // vC= 1785 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100010; // iC=  546 
// vC = 14'b0000011011010110; // vC= 1750 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111011; // iC=  507 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001011; // iC=  395 
// vC = 14'b0000011000101000; // vC= 1576 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011101; // iC=  285 
// vC = 14'b0000011000101011; // vC= 1579 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001001; // iC=  393 
// vC = 14'b0000010111100000; // vC= 1504 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101000; // iC=  360 
// vC = 14'b0000011011001001; // vC= 1737 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111110; // iC=  318 
// vC = 14'b0000010111011010; // vC= 1498 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000011; // iC=  259 
// vC = 14'b0000011000001111; // vC= 1551 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101100; // iC=  300 
// vC = 14'b0000011001001101; // vC= 1613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111011; // iC=  315 
// vC = 14'b0000011011110011; // vC= 1779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010010; // iC=  338 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001000; // iC=  392 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100110; // iC=  166 
// vC = 14'b0000011100001110; // vC= 1806 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000001; // iC=  449 
// vC = 14'b0000011011100101; // vC= 1765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001010; // iC=  138 
// vC = 14'b0000011010001000; // vC= 1672 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110111; // iC=  119 
// vC = 14'b0000011010100001; // vC= 1697 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011011; // iC=  347 
// vC = 14'b0000011100011010; // vC= 1818 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011011010; // iC=  218 
// vC = 14'b0000011000001111; // vC= 1551 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000111; // iC=  327 
// vC = 14'b0000011011000111; // vC= 1735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001101; // iC=  141 
// vC = 14'b0000011000011000; // vC= 1560 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001110; // iC=  334 
// vC = 14'b0000011011000000; // vC= 1728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110110; // iC=  246 
// vC = 14'b0000010111110101; // vC= 1525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010111; // iC=  151 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001001; // iC=  265 
// vC = 14'b0000011011110011; // vC= 1779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110011; // iC=  243 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011111; // iC=  159 
// vC = 14'b0000011000001101; // vC= 1549 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001010; // iC=   74 
// vC = 14'b0000011000010001; // vC= 1553 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000111101; // iC=   61 
// vC = 14'b0000011011011010; // vC= 1754 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110101; // iC=  181 
// vC = 14'b0000011001000001; // vC= 1601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111011; // iC=  123 
// vC = 14'b0000011011110100; // vC= 1780 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000110010; // iC=   50 
// vC = 14'b0000011000011100; // vC= 1564 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000110; // iC=    6 
// vC = 14'b0000011001000011; // vC= 1603 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111001; // iC=  -71 
// vC = 14'b0000011010101101; // vC= 1709 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100000; // iC=  -96 
// vC = 14'b0000011000001011; // vC= 1547 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100101; // iC=  -27 
// vC = 14'b0000011011001010; // vC= 1738 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101110100; // iC= -140 
// vC = 14'b0000011000011110; // vC= 1566 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111111; // iC=   -1 
// vC = 14'b0000010111100110; // vC= 1510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011111; // iC= -225 
// vC = 14'b0000011000100010; // vC= 1570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001101; // iC= -115 
// vC = 14'b0000011010011001; // vC= 1689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110110101; // iC=  -75 
// vC = 14'b0000011001001010; // vC= 1610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000111; // iC= -249 
// vC = 14'b0000010111011110; // vC= 1502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010100; // iC= -364 
// vC = 14'b0000011001001111; // vC= 1615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010100; // iC= -108 
// vC = 14'b0000011000001110; // vC= 1550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101111; // iC= -273 
// vC = 14'b0000010111011110; // vC= 1502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010101010; // iC= -342 
// vC = 14'b0000011010111101; // vC= 1725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110001; // iC= -463 
// vC = 14'b0000011010110110; // vC= 1718 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000001; // iC= -447 
// vC = 14'b0000011010110000; // vC= 1712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011011; // iC= -485 
// vC = 14'b0000011000110111; // vC= 1591 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000011; // iC= -381 
// vC = 14'b0000011001111101; // vC= 1661 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001111; // iC= -305 
// vC = 14'b0000011010000110; // vC= 1670 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100001; // iC= -351 
// vC = 14'b0000011001011100; // vC= 1628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100100; // iC= -348 
// vC = 14'b0000011000010001; // vC= 1553 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001100; // iC= -564 
// vC = 14'b0000010111110111; // vC= 1527 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010101111; // iC= -337 
// vC = 14'b0000011010011011; // vC= 1691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101011; // iC= -405 
// vC = 14'b0000011011110110; // vC= 1782 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001110; // iC= -434 
// vC = 14'b0000011001111110; // vC= 1662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001111; // iC= -433 
// vC = 14'b0000010111111111; // vC= 1535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001100; // iC= -628 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010101; // iC= -555 
// vC = 14'b0000010111110010; // vC= 1522 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100101; // iC= -603 
// vC = 14'b0000011011011010; // vC= 1754 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011001; // iC= -679 
// vC = 14'b0000011001111010; // vC= 1658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100101; // iC= -603 
// vC = 14'b0000011010000101; // vC= 1669 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101011; // iC= -789 
// vC = 14'b0000011011101100; // vC= 1772 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001000; // iC= -568 
// vC = 14'b0000011001011110; // vC= 1630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011010; // iC= -870 
// vC = 14'b0000010111111100; // vC= 1532 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000110; // iC= -762 
// vC = 14'b0000011010111001; // vC= 1721 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111110; // iC= -834 
// vC = 14'b0000010110111011; // vC= 1467 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000101; // iC= -827 
// vC = 14'b0000010110011101; // vC= 1437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101011; // iC= -981 
// vC = 14'b0000011001000001; // vC= 1601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011011; // iC= -741 
// vC = 14'b0000011010011111; // vC= 1695 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000110; // iC= -954 
// vC = 14'b0000010111101001; // vC= 1513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100101; // iC= -923 
// vC = 14'b0000011010010101; // vC= 1685 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000010; // iC= -958 
// vC = 14'b0000011001001111; // vC= 1615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011110; // iC= -866 
// vC = 14'b0000011010101011; // vC= 1707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101101; // iC= -851 
// vC = 14'b0000010111001010; // vC= 1482 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100000; // iC= -992 
// vC = 14'b0000010110010010; // vC= 1426 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b0000011000010111; // vC= 1559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100010; // iC= -926 
// vC = 14'b0000011000110000; // vC= 1584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010110; // iC=-1130 
// vC = 14'b0000010110001111; // vC= 1423 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010000; // iC= -944 
// vC = 14'b0000011010001100; // vC= 1676 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001000; // iC=-1208 
// vC = 14'b0000010101100101; // vC= 1381 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010110; // iC=-1066 
// vC = 14'b0000011010011110; // vC= 1694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011100; // iC=-1252 
// vC = 14'b0000010110100111; // vC= 1447 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100100; // iC=-1116 
// vC = 14'b0000011010001100; // vC= 1676 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011111; // iC= -993 
// vC = 14'b0000011010001011; // vC= 1675 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100111; // iC=-1305 
// vC = 14'b0000010111011101; // vC= 1501 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101101; // iC=-1171 
// vC = 14'b0000010110100010; // vC= 1442 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111111; // iC=-1089 
// vC = 14'b0000010110000111; // vC= 1415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010110; // iC=-1066 
// vC = 14'b0000010111111101; // vC= 1533 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101011; // iC=-1173 
// vC = 14'b0000011001001110; // vC= 1614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101110; // iC=-1362 
// vC = 14'b0000010110001000; // vC= 1416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001001; // iC=-1335 
// vC = 14'b0000010101100101; // vC= 1381 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010111; // iC=-1193 
// vC = 14'b0000010110110101; // vC= 1461 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011100; // iC=-1188 
// vC = 14'b0000010101000011; // vC= 1347 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001111; // iC=-1265 
// vC = 14'b0000010111111000; // vC= 1528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111000; // iC=-1288 
// vC = 14'b0000010100100111; // vC= 1319 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100010; // iC=-1310 
// vC = 14'b0000010110111001; // vC= 1465 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110111; // iC=-1225 
// vC = 14'b0000010100111000; // vC= 1336 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100110; // iC=-1498 
// vC = 14'b0000010111110100; // vC= 1524 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111001; // iC=-1287 
// vC = 14'b0000010111000100; // vC= 1476 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110001; // iC=-1487 
// vC = 14'b0000010100001001; // vC= 1289 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001010; // iC=-1590 
// vC = 14'b0000010110011111; // vC= 1439 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110010; // iC=-1486 
// vC = 14'b0000010100001111; // vC= 1295 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001101; // iC=-1587 
// vC = 14'b0000010101001001; // vC= 1353 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111000; // iC=-1416 
// vC = 14'b0000010111100101; // vC= 1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011010; // iC=-1638 
// vC = 14'b0000010111011100; // vC= 1500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010101; // iC=-1579 
// vC = 14'b0000010011010000; // vC= 1232 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011101; // iC=-1571 
// vC = 14'b0000011000000011; // vC= 1539 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001011; // iC=-1653 
// vC = 14'b0000010011110000; // vC= 1264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100011; // iC=-1565 
// vC = 14'b0000010100110101; // vC= 1333 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110110; // iC=-1674 
// vC = 14'b0000010100110001; // vC= 1329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000111; // iC=-1593 
// vC = 14'b0000010100111100; // vC= 1340 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b0000010110000000; // vC= 1408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100110; // iC=-1434 
// vC = 14'b0000010100000111; // vC= 1287 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100000; // iC=-1568 
// vC = 14'b0000010101100010; // vC= 1378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000011; // iC=-1725 
// vC = 14'b0000010100100000; // vC= 1312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110101; // iC=-1611 
// vC = 14'b0000010100111000; // vC= 1336 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111101; // iC=-1731 
// vC = 14'b0000010110100100; // vC= 1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110111; // iC=-1673 
// vC = 14'b0000010110101001; // vC= 1449 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b0000010010010110; // vC= 1174 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011010; // iC=-1638 
// vC = 14'b0000010001111110; // vC= 1150 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010010; // iC=-1774 
// vC = 14'b0000010001101110; // vC= 1134 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000001; // iC=-1855 
// vC = 14'b0000010001110100; // vC= 1140 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110000; // iC=-1744 
// vC = 14'b0000010101011011; // vC= 1371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111110; // iC=-1666 
// vC = 14'b0000010011110010; // vC= 1266 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010110; // iC=-1706 
// vC = 14'b0000010101000111; // vC= 1351 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011000; // iC=-1640 
// vC = 14'b0000010101000001; // vC= 1345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011011; // iC=-1765 
// vC = 14'b0000010101001101; // vC= 1357 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100001; // iC=-1631 
// vC = 14'b0000010010001010; // vC= 1162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000101; // iC=-1659 
// vC = 14'b0000010011101110; // vC= 1262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011110; // iC=-1698 
// vC = 14'b0000010100100100; // vC= 1316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110101; // iC=-1803 
// vC = 14'b0000010011110111; // vC= 1271 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110000; // iC=-1872 
// vC = 14'b0000010010111001; // vC= 1209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111000; // iC=-1736 
// vC = 14'b0000010010100111; // vC= 1191 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000010011011100; // vC= 1244 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110111; // iC=-1865 
// vC = 14'b0000010001111000; // vC= 1144 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001111; // iC=-1713 
// vC = 14'b0000010000101111; // vC= 1071 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011001; // iC=-1895 
// vC = 14'b0000010011100000; // vC= 1248 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000110; // iC=-1978 
// vC = 14'b0000010010011100; // vC= 1180 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011011; // iC=-1765 
// vC = 14'b0000010011011111; // vC= 1247 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111101; // iC=-1923 
// vC = 14'b0000010001101100; // vC= 1132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b0000010010111010; // vC= 1210 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110100; // iC=-1676 
// vC = 14'b0000010001111110; // vC= 1150 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000010011001110; // vC= 1230 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101000; // iC=-1688 
// vC = 14'b0000010001110001; // vC= 1137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110000; // iC=-1744 
// vC = 14'b0000001110011000; // vC=  920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101111; // iC=-2001 
// vC = 14'b0000010000101111; // vC= 1071 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110011; // iC=-1997 
// vC = 14'b0000001111001101; // vC=  973 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110001; // iC=-1999 
// vC = 14'b0000010010001110; // vC= 1166 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011000; // iC=-1832 
// vC = 14'b0000010010101000; // vC= 1192 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001111; // iC=-1841 
// vC = 14'b0000001110001010; // vC=  906 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010101; // iC=-1707 
// vC = 14'b0000010001110111; // vC= 1143 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b0000001110111101; // vC=  957 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011000; // iC=-1768 
// vC = 14'b0000001110101010; // vC=  938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010011; // iC=-1773 
// vC = 14'b0000001111100001; // vC=  993 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110010; // iC=-1870 
// vC = 14'b0000001101101111; // vC=  879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101011; // iC=-1877 
// vC = 14'b0000001101010010; // vC=  850 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b0000001110010101; // vC=  917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b0000001110111100; // vC=  956 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b0000001110010011; // vC=  915 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b0000001100110011; // vC=  819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b0000001110000101; // vC=  901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000001100011111; // vC=  799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011010; // iC=-1894 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101010; // iC=-1878 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b0000010000100001; // vC= 1057 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011001; // iC=-1767 
// vC = 14'b0000010000010011; // vC= 1043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001100; // iC=-1780 
// vC = 14'b0000001101001001; // vC=  841 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110111; // iC=-1801 
// vC = 14'b0000010000011100; // vC= 1052 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b0000001100011110; // vC=  798 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010111; // iC=-1897 
// vC = 14'b0000010000000111; // vC= 1031 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000101; // iC=-1787 
// vC = 14'b0000001011110100; // vC=  756 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b0000001111010001; // vC=  977 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001111; // iC=-1905 
// vC = 14'b0000001101110010; // vC=  882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000001110011000; // vC=  920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011111; // iC=-1825 
// vC = 14'b0000001100011101; // vC=  797 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111101; // iC=-1795 
// vC = 14'b0000001100111010; // vC=  826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b0000001010101100; // vC=  684 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011000; // iC=-2024 
// vC = 14'b0000001010100111; // vC=  679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b0000001100111010; // vC=  826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010100; // iC=-1772 
// vC = 14'b0000001110010111; // vC=  919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b0000001010110010; // vC=  690 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b0000001110100110; // vC=  934 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b0000001101000001; // vC=  833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001001; // iC=-2039 
// vC = 14'b0000001011011001; // vC=  729 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b0000001010010011; // vC=  659 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b0000001011001111; // vC=  719 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000001011110010; // vC=  754 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b0000001011000111; // vC=  711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b0000001011110000; // vC=  752 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b0000001010100100; // vC=  676 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000100; // iC=-1788 
// vC = 14'b0000001011010100; // vC=  724 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b0000001101010101; // vC=  853 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111001; // iC=-1799 
// vC = 14'b0000001010111111; // vC=  703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111101; // iC=-1795 
// vC = 14'b0000001001101001; // vC=  617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000010; // iC=-1790 
// vC = 14'b0000001000101001; // vC=  553 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100010; // iC=-2014 
// vC = 14'b0000001100100110; // vC=  806 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b0000001010000000; // vC=  640 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b0000001010000110; // vC=  646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b0000001001110011; // vC=  627 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b0000001000010010; // vC=  530 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001110; // iC=-1842 
// vC = 14'b0000000111110011; // vC=  499 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b0000001010100010; // vC=  674 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011111; // iC=-1825 
// vC = 14'b0000000110111010; // vC=  442 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001010; // iC=-1910 
// vC = 14'b0000001000100001; // vC=  545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b0000001010011111; // vC=  671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b0000001010001000; // vC=  648 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110000; // iC=-2000 
// vC = 14'b0000000111101010; // vC=  490 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b0000001001110010; // vC=  626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b0000000110010011; // vC=  403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010100; // iC=-1900 
// vC = 14'b0000000111011101; // vC=  477 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b0000000111111110; // vC=  510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010001; // iC=-2031 
// vC = 14'b0000001010010100; // vC=  660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b0000001001101111; // vC=  623 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000011; // iC=-1853 
// vC = 14'b0000000101111001; // vC=  377 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110101; // iC=-1867 
// vC = 14'b0000000101111100; // vC=  380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b0000001001000000; // vC=  576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b0000001001101000; // vC=  616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b0000000111111111; // vC=  511 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000000100111010; // vC=  314 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010001; // iC=-1775 
// vC = 14'b0000000111110110; // vC=  502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b0000000110101100; // vC=  428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b0000000100110100; // vC=  308 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111101; // iC=-1923 
// vC = 14'b0000000100111001; // vC=  313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b0000000110101111; // vC=  431 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111010; // iC=-1862 
// vC = 14'b0000000101100111; // vC=  359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110011; // iC=-1805 
// vC = 14'b0000000111111101; // vC=  509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000000111011001; // vC=  473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b0000001000100011; // vC=  547 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b0000000101011101; // vC=  349 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101100; // iC=-2068 
// vC = 14'b0000000100011110; // vC=  286 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b0000000110001001; // vC=  393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b0000000100000111; // vC=  263 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000000110001110; // vC=  398 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b0000000100011011; // vC=  283 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000000110011000; // vC=  408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b0000000100011010; // vC=  282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100100; // iC=-1820 
// vC = 14'b0000000011010010; // vC=  210 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000000110100110; // vC=  422 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000110; // iC=-1978 
// vC = 14'b0000000100110000; // vC=  304 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b0000000110011111; // vC=  415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b0000000110011000; // vC=  408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110001; // iC=-1743 
// vC = 14'b0000000101010101; // vC=  341 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b0000000110011101; // vC=  413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000000011010000; // vC=  208 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b0000000110010101; // vC=  405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b0000000010111001; // vC=  185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b0000000100110110; // vC=  310 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100010; // iC=-1758 
// vC = 14'b0000000010011100; // vC=  156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b0000000101101001; // vC=  361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b0000000001100100; // vC=  100 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011010; // iC=-1766 
// vC = 14'b0000000000110010; // vC=   50 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111100; // iC=-1860 
// vC = 14'b0000000001001011; // vC=   75 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101100; // iC=-1748 
// vC = 14'b0000000011000110; // vC=  198 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100111; // iC=-1881 
// vC = 14'b0000000011111101; // vC=  253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011111; // iC=-1825 
// vC = 14'b0000000011110100; // vC=  244 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001110; // iC=-1842 
// vC = 14'b0000000001001011; // vC=   75 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000101; // iC=-1851 
// vC = 14'b0000000000011111; // vC=   31 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101001; // iC=-2007 
// vC = 14'b0000000011101110; // vC=  238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b1111111111111011; // vC=   -5 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110100; // iC=-1740 
// vC = 14'b0000000000110100; // vC=   52 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001111; // iC=-1905 
// vC = 14'b0000000000111111; // vC=   63 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b0000000011110111; // vC=  247 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011000; // iC=-1832 
// vC = 14'b0000000010010100; // vC=  148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000001; // iC=-1855 
// vC = 14'b0000000001001001; // vC=   73 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b0000000001101110; // vC=  110 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000110; // iC=-1914 
// vC = 14'b0000000000110110; // vC=   54 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100011; // iC=-1757 
// vC = 14'b0000000010011000; // vC=  152 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110100; // iC=-1932 
// vC = 14'b1111111110110110; // vC=  -74 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000110; // iC=-1978 
// vC = 14'b0000000000111111; // vC=   63 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110000; // iC=-2000 
// vC = 14'b0000000001001101; // vC=   77 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b1111111111010011; // vC=  -45 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000010; // iC=-1918 
// vC = 14'b0000000000110001; // vC=   49 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b0000000000010000; // vC=   16 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010110; // iC=-1770 
// vC = 14'b0000000001100000; // vC=   96 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b0000000010001011; // vC=  139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111110; // iC=-1794 
// vC = 14'b1111111110101001; // vC=  -87 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b0000000000110011; // vC=   51 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011111; // iC=-1761 
// vC = 14'b0000000001111011; // vC=  123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b1111111101111100; // vC= -132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b0000000000001100; // vC=   12 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b1111111111100111; // vC=  -25 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b0000000000010101; // vC=   21 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101010; // iC=-1750 
// vC = 14'b1111111101101100; // vC= -148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b1111111110001111; // vC= -113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011110; // iC=-1698 
// vC = 14'b1111111111010011; // vC=  -45 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b1111111110100000; // vC=  -96 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001011; // iC=-1781 
// vC = 14'b1111111100101100; // vC= -212 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b1111111101101100; // vC= -148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010010; // iC=-1710 
// vC = 14'b1111111111110001; // vC=  -15 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b1111111101111011; // vC= -133 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100000; // iC=-1952 
// vC = 14'b1111111110110001; // vC=  -79 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100111; // iC=-1817 
// vC = 14'b1111111110001110; // vC= -114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b1111111100100111; // vC= -217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b1111111100011111; // vC= -225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b1111111011010110; // vC= -298 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101011; // iC=-1749 
// vC = 14'b1111111101000000; // vC= -192 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100001; // iC=-1887 
// vC = 14'b1111111100100011; // vC= -221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000111; // iC=-1721 
// vC = 14'b1111111010111111; // vC= -321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b1111111011010100; // vC= -300 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111111; // iC=-1729 
// vC = 14'b1111111100011000; // vC= -232 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100011; // iC=-1757 
// vC = 14'b1111111011000110; // vC= -314 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111110; // iC=-1794 
// vC = 14'b1111111111001110; // vC=  -50 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110000; // iC=-1936 
// vC = 14'b1111111111000001; // vC=  -63 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101010; // iC=-1878 
// vC = 14'b1111111011111000; // vC= -264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b1111111110001100; // vC= -116 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b1111111101111011; // vC= -133 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b1111111100000011; // vC= -253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001000; // iC=-1656 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100000; // iC=-1696 
// vC = 14'b1111111110000111; // vC= -121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011001; // iC=-1767 
// vC = 14'b1111111010111101; // vC= -323 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b1111111001011011; // vC= -421 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111111011101111; // vC= -273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000001; // iC=-1791 
// vC = 14'b1111111011111110; // vC= -258 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b1111111101010011; // vC= -173 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110010; // iC=-1678 
// vC = 14'b1111111010010001; // vC= -367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000011; // iC=-1725 
// vC = 14'b1111111011100001; // vC= -287 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101111; // iC=-1617 
// vC = 14'b1111111000111001; // vC= -455 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000010; // iC=-1726 
// vC = 14'b1111111001100001; // vC= -415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000101; // iC=-1851 
// vC = 14'b1111111001011110; // vC= -418 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010110; // iC=-1898 
// vC = 14'b1111111010001111; // vC= -369 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100111; // iC=-1689 
// vC = 14'b1111111100111101; // vC= -195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010101; // iC=-1771 
// vC = 14'b1111110111111101; // vC= -515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110100; // iC=-1804 
// vC = 14'b1111111010011001; // vC= -359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010110; // iC=-1898 
// vC = 14'b1111111100100100; // vC= -220 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000101; // iC=-1659 
// vC = 14'b1111111011100100; // vC= -284 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010011; // iC=-1709 
// vC = 14'b1111111001000010; // vC= -446 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010011; // iC=-1773 
// vC = 14'b1111110111101110; // vC= -530 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b1111111011001110; // vC= -306 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b1111111001011000; // vC= -424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001010; // iC=-1782 
// vC = 14'b1111111001110110; // vC= -394 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100101; // iC=-1755 
// vC = 14'b1111111001111001; // vC= -391 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011000; // iC=-1640 
// vC = 14'b1111111000111011; // vC= -453 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010100; // iC=-1772 
// vC = 14'b1111111001001110; // vC= -434 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b1111111011010010; // vC= -302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000101; // iC=-1659 
// vC = 14'b1111110110011010; // vC= -614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111111; // iC=-1601 
// vC = 14'b1111110111111000; // vC= -520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011000; // iC=-1704 
// vC = 14'b1111110110101111; // vC= -593 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100111; // iC=-1817 
// vC = 14'b1111110111111000; // vC= -520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111101; // iC=-1731 
// vC = 14'b1111111001010011; // vC= -429 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011010; // iC=-1830 
// vC = 14'b1111110101110101; // vC= -651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110111; // iC=-1609 
// vC = 14'b1111111001011000; // vC= -424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001101; // iC=-1715 
// vC = 14'b1111110101101110; // vC= -658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101110; // iC=-1810 
// vC = 14'b1111111001101010; // vC= -406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100101; // iC=-1691 
// vC = 14'b1111110110110110; // vC= -586 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011010; // iC=-1638 
// vC = 14'b1111111001010000; // vC= -432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101111; // iC=-1681 
// vC = 14'b1111110110101000; // vC= -600 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111111; // iC=-1537 
// vC = 14'b1111111001111000; // vC= -392 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110011; // iC=-1549 
// vC = 14'b1111110101111010; // vC= -646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001001; // iC=-1655 
// vC = 14'b1111111001101101; // vC= -403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010100; // iC=-1644 
// vC = 14'b1111110110111101; // vC= -579 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111110; // iC=-1666 
// vC = 14'b1111110111110110; // vC= -522 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001111; // iC=-1713 
// vC = 14'b1111110111111000; // vC= -520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001001; // iC=-1655 
// vC = 14'b1111110111000011; // vC= -573 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011000; // iC=-1768 
// vC = 14'b1111110110110000; // vC= -592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b1111110101000101; // vC= -699 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101100; // iC=-1556 
// vC = 14'b1111110100000101; // vC= -763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000011; // iC=-1533 
// vC = 14'b1111110111100011; // vC= -541 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000110; // iC=-1594 
// vC = 14'b1111110101101001; // vC= -663 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101000; // iC=-1560 
// vC = 14'b1111110110110011; // vC= -589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100100; // iC=-1500 
// vC = 14'b1111110100010100; // vC= -748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000111; // iC=-1721 
// vC = 14'b1111110100001011; // vC= -757 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011000; // iC=-1768 
// vC = 14'b1111110101110110; // vC= -650 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000101; // iC=-1659 
// vC = 14'b1111110101011101; // vC= -675 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000010; // iC=-1662 
// vC = 14'b1111110101000110; // vC= -698 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100000; // iC=-1632 
// vC = 14'b1111110100000001; // vC= -767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011010; // iC=-1574 
// vC = 14'b1111110100011000; // vC= -744 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001101; // iC=-1651 
// vC = 14'b1111110011100001; // vC= -799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110100; // iC=-1484 
// vC = 14'b1111110101101000; // vC= -664 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000100; // iC=-1596 
// vC = 14'b1111110110110111; // vC= -585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100000; // iC=-1568 
// vC = 14'b1111110011101100; // vC= -788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000110; // iC=-1594 
// vC = 14'b1111110100100011; // vC= -733 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101011; // iC=-1749 
// vC = 14'b1111110100010001; // vC= -751 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000111; // iC=-1593 
// vC = 14'b1111110011101000; // vC= -792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010100; // iC=-1772 
// vC = 14'b1111110110110101; // vC= -587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100000; // iC=-1696 
// vC = 14'b1111110010011010; // vC= -870 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111110; // iC=-1474 
// vC = 14'b1111110110110010; // vC= -590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011010; // iC=-1638 
// vC = 14'b1111110101100101; // vC= -667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110101; // iC=-1675 
// vC = 14'b1111110010010101; // vC= -875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010010; // iC=-1518 
// vC = 14'b1111110100110110; // vC= -714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010000; // iC=-1648 
// vC = 14'b1111110101010011; // vC= -685 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100110; // iC=-1434 
// vC = 14'b1111110110001110; // vC= -626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011101; // iC=-1443 
// vC = 14'b1111110001101001; // vC= -919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000111; // iC=-1465 
// vC = 14'b1111110101001001; // vC= -695 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100110; // iC=-1562 
// vC = 14'b1111110101101100; // vC= -660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111010; // iC=-1606 
// vC = 14'b1111110010111111; // vC= -833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000011; // iC=-1597 
// vC = 14'b1111110010101000; // vC= -856 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001111; // iC=-1713 
// vC = 14'b1111110100101001; // vC= -727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010100; // iC=-1452 
// vC = 14'b1111110011011111; // vC= -801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101001; // iC=-1495 
// vC = 14'b1111110100111110; // vC= -706 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100110; // iC=-1498 
// vC = 14'b1111110010101111; // vC= -849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011010; // iC=-1574 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100111; // iC=-1433 
// vC = 14'b1111110100110110; // vC= -714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010001; // iC=-1391 
// vC = 14'b1111110100101101; // vC= -723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001000; // iC=-1400 
// vC = 14'b1111110100110011; // vC= -717 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000011; // iC=-1469 
// vC = 14'b1111110001100101; // vC= -923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110000; // iC=-1488 
// vC = 14'b1111110001111010; // vC= -902 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110011; // iC=-1549 
// vC = 14'b1111110001111100; // vC= -900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010101; // iC=-1451 
// vC = 14'b1111110000100011; // vC= -989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011010; // iC=-1510 
// vC = 14'b1111110001111001; // vC= -903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110110; // iC=-1546 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000001; // iC=-1535 
// vC = 14'b1111110010011000; // vC= -872 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000010; // iC=-1470 
// vC = 14'b1111110000001011; // vC=-1013 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111100; // iC=-1604 
// vC = 14'b1111101111000101; // vC=-1083 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110101; // iC=-1355 
// vC = 14'b1111101110111110; // vC=-1090 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100001; // iC=-1375 
// vC = 14'b1111110010010000; // vC= -880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000001; // iC=-1599 
// vC = 14'b1111101111001010; // vC=-1078 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001001; // iC=-1335 
// vC = 14'b1111110001011010; // vC= -934 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011010; // iC=-1638 
// vC = 14'b1111110011000101; // vC= -827 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001000; // iC=-1336 
// vC = 14'b1111110010001101; // vC= -883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101100; // iC=-1556 
// vC = 14'b1111110010000100; // vC= -892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110111; // iC=-1609 
// vC = 14'b1111101111110000; // vC=-1040 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010110; // iC=-1578 
// vC = 14'b1111110011000010; // vC= -830 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101001; // iC=-1431 
// vC = 14'b1111110000110001; // vC= -975 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110010; // iC=-1358 
// vC = 14'b1111101111011100; // vC=-1060 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110111; // iC=-1609 
// vC = 14'b1111110010100101; // vC= -859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111010; // iC=-1350 
// vC = 14'b1111101110011011; // vC=-1125 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001001; // iC=-1335 
// vC = 14'b1111110001010100; // vC= -940 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111010; // iC=-1414 
// vC = 14'b1111110001101101; // vC= -915 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101100; // iC=-1556 
// vC = 14'b1111101111111110; // vC=-1026 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110011; // iC=-1485 
// vC = 14'b1111110000101010; // vC= -982 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010011; // iC=-1389 
// vC = 14'b1111101110101111; // vC=-1105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100111; // iC=-1497 
// vC = 14'b1111101101101000; // vC=-1176 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011110; // iC=-1442 
// vC = 14'b1111110000110001; // vC= -975 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011111; // iC=-1505 
// vC = 14'b1111110001011010; // vC= -934 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001001; // iC=-1271 
// vC = 14'b1111101111000010; // vC=-1086 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001100; // iC=-1332 
// vC = 14'b1111101111001001; // vC=-1079 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110000; // iC=-1360 
// vC = 14'b1111101101011111; // vC=-1185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000001; // iC=-1343 
// vC = 14'b1111101110110011; // vC=-1101 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111111; // iC=-1537 
// vC = 14'b1111110000110001; // vC= -975 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111010; // iC=-1286 
// vC = 14'b1111110001100001; // vC= -927 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011010; // iC=-1382 
// vC = 14'b1111110001011000; // vC= -936 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101010; // iC=-1302 
// vC = 14'b1111110000110110; // vC= -970 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000010; // iC=-1406 
// vC = 14'b1111110001001000; // vC= -952 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110101; // iC=-1291 
// vC = 14'b1111101100100100; // vC=-1244 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000100; // iC=-1276 
// vC = 14'b1111101100100011; // vC=-1245 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000001; // iC=-1471 
// vC = 14'b1111101110100010; // vC=-1118 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010001; // iC=-1391 
// vC = 14'b1111101111111100; // vC=-1028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001011; // iC=-1461 
// vC = 14'b1111101100010101; // vC=-1259 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000110; // iC=-1274 
// vC = 14'b1111110000101111; // vC= -977 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110111; // iC=-1289 
// vC = 14'b1111101110010010; // vC=-1134 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011100; // iC=-1444 
// vC = 14'b1111101111100111; // vC=-1049 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010011; // iC=-1261 
// vC = 14'b1111101111010000; // vC=-1072 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001011; // iC=-1269 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101110; // iC=-1426 
// vC = 14'b1111110000010100; // vC=-1004 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011000; // iC=-1192 
// vC = 14'b1111101101001101; // vC=-1203 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101111; // iC=-1169 
// vC = 14'b1111101011001011; // vC=-1333 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110110; // iC=-1354 
// vC = 14'b1111101100010100; // vC=-1260 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101100; // iC=-1236 
// vC = 14'b1111101111011000; // vC=-1064 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110001; // iC=-1167 
// vC = 14'b1111101011001011; // vC=-1333 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101011; // iC=-1173 
// vC = 14'b1111101101110111; // vC=-1161 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101000; // iC=-1176 
// vC = 14'b1111101011010011; // vC=-1325 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010110; // iC=-1258 
// vC = 14'b1111101110111000; // vC=-1096 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010111; // iC=-1257 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010001; // iC=-1391 
// vC = 14'b1111101101000100; // vC=-1212 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110101; // iC=-1419 
// vC = 14'b1111101011001100; // vC=-1332 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101100; // iC=-1236 
// vC = 14'b1111101011000110; // vC=-1338 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011110; // iC=-1122 
// vC = 14'b1111101011010101; // vC=-1323 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101111; // iC=-1361 
// vC = 14'b1111101110100110; // vC=-1114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010011; // iC=-1133 
// vC = 14'b1111101101111001; // vC=-1159 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101011; // iC=-1173 
// vC = 14'b1111101100110001; // vC=-1231 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111110; // iC=-1154 
// vC = 14'b1111101100101011; // vC=-1237 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011101; // iC=-1379 
// vC = 14'b1111101010000101; // vC=-1403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100100; // iC=-1116 
// vC = 14'b1111101100010110; // vC=-1258 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101001; // iC=-1175 
// vC = 14'b1111101010000111; // vC=-1401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001010; // iC=-1142 
// vC = 14'b1111101010110110; // vC=-1354 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100000; // iC=-1248 
// vC = 14'b1111101011001101; // vC=-1331 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000011; // iC=-1085 
// vC = 14'b1111101010010101; // vC=-1387 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100111; // iC=-1305 
// vC = 14'b1111101110001100; // vC=-1140 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110100; // iC=-1292 
// vC = 14'b1111101100111011; // vC=-1221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010011; // iC=-1325 
// vC = 14'b1111101011110111; // vC=-1289 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101010; // iC=-1302 
// vC = 14'b1111101011001110; // vC=-1330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011111; // iC=-1121 
// vC = 14'b1111101100111000; // vC=-1224 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010111; // iC=-1257 
// vC = 14'b1111101001111110; // vC=-1410 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110000; // iC=-1104 
// vC = 14'b1111101011100011; // vC=-1309 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001001; // iC=-1143 
// vC = 14'b1111101011010001; // vC=-1327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001110; // iC=-1074 
// vC = 14'b1111101011100110; // vC=-1306 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010011; // iC=-1197 
// vC = 14'b1111101001111001; // vC=-1415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011010; // iC=-1190 
// vC = 14'b1111101011111001; // vC=-1287 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011001; // iC=-1063 
// vC = 14'b1111101011011100; // vC=-1316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001111; // iC=-1201 
// vC = 14'b1111101011011011; // vC=-1317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100111; // iC=-1049 
// vC = 14'b1111101010001010; // vC=-1398 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101101; // iC=-1107 
// vC = 14'b1111101011101001; // vC=-1303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011101; // iC=-1059 
// vC = 14'b1111101001010010; // vC=-1454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001101; // iC=-1075 
// vC = 14'b1111101011011111; // vC=-1313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111010; // iC=-1094 
// vC = 14'b1111101011001000; // vC=-1336 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010001; // iC=-1007 
// vC = 14'b1111101000000001; // vC=-1535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101100; // iC= -980 
// vC = 14'b1111101000111101; // vC=-1475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101100; // iC=-1108 
// vC = 14'b1111101010111111; // vC=-1345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110110; // iC=-1162 
// vC = 14'b1111101010010000; // vC=-1392 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111001; // iC=-1159 
// vC = 14'b1111101100110010; // vC=-1230 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111011; // iC= -965 
// vC = 14'b1111101000111111; // vC=-1473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011001; // iC=-1127 
// vC = 14'b1111101000100000; // vC=-1504 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010100; // iC=-1068 
// vC = 14'b1111101000100100; // vC=-1500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010001; // iC=-1071 
// vC = 14'b1111101100011101; // vC=-1251 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001101; // iC=-1011 
// vC = 14'b1111100111110010; // vC=-1550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010001; // iC=-1007 
// vC = 14'b1111101001011000; // vC=-1448 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010110; // iC=-1130 
// vC = 14'b1111101000100100; // vC=-1500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101011; // iC=-1109 
// vC = 14'b1111101000111101; // vC=-1475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110001; // iC= -975 
// vC = 14'b1111101010110111; // vC=-1353 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111111; // iC=-1025 
// vC = 14'b1111101011000100; // vC=-1340 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011000; // iC= -936 
// vC = 14'b1111101010001111; // vC=-1393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011000; // iC=-1128 
// vC = 14'b1111101000000100; // vC=-1532 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100111; // iC= -985 
// vC = 14'b1111101011011011; // vC=-1317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110101; // iC= -971 
// vC = 14'b1111101001100010; // vC=-1438 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010010; // iC=-1006 
// vC = 14'b1111100110110111; // vC=-1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110111; // iC=-1097 
// vC = 14'b1111100110101010; // vC=-1622 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110001; // iC=-1167 
// vC = 14'b1111101000101111; // vC=-1489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001011; // iC=-1013 
// vC = 14'b1111101010000000; // vC=-1408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b1111101010101111; // vC=-1361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011011; // iC=-1125 
// vC = 14'b1111101000011110; // vC=-1506 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111101; // iC= -899 
// vC = 14'b1111100110100100; // vC=-1628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b1111101010101011; // vC=-1365 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111100; // iC= -900 
// vC = 14'b1111100110001100; // vC=-1652 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110110; // iC= -842 
// vC = 14'b1111100111101011; // vC=-1557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000001; // iC=-1087 
// vC = 14'b1111100111110111; // vC=-1545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011101; // iC= -867 
// vC = 14'b1111101001110010; // vC=-1422 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100010; // iC=-1118 
// vC = 14'b1111101010101011; // vC=-1365 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010100; // iC= -876 
// vC = 14'b1111101001001011; // vC=-1461 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010101; // iC= -939 
// vC = 14'b1111101010001111; // vC=-1393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101010; // iC=-1046 
// vC = 14'b1111101010010110; // vC=-1386 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101101; // iC= -979 
// vC = 14'b1111100110111111; // vC=-1601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111000; // iC= -776 
// vC = 14'b1111101010010111; // vC=-1385 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101000; // iC= -984 
// vC = 14'b1111100111011010; // vC=-1574 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000111; // iC= -825 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111011; // iC= -837 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111100; // iC= -836 
// vC = 14'b1111101010001101; // vC=-1395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b1111101001011010; // vC=-1446 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001101; // iC= -819 
// vC = 14'b1111101001100101; // vC=-1435 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101111; // iC= -977 
// vC = 14'b1111100101111010; // vC=-1670 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111000; // iC= -840 
// vC = 14'b1111101000001001; // vC=-1527 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101011; // iC= -917 
// vC = 14'b1111100110011001; // vC=-1639 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000111; // iC= -825 
// vC = 14'b1111101001011011; // vC=-1445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001111; // iC= -881 
// vC = 14'b1111101000000101; // vC=-1531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010111; // iC= -937 
// vC = 14'b1111100101000111; // vC=-1721 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000010; // iC= -766 
// vC = 14'b1111101001011110; // vC=-1442 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010011; // iC= -877 
// vC = 14'b1111100111100010; // vC=-1566 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110001; // iC= -719 
// vC = 14'b1111100111100001; // vC=-1567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010110; // iC= -746 
// vC = 14'b1111100111010111; // vC=-1577 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101010; // iC= -854 
// vC = 14'b1111101000111010; // vC=-1478 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110010; // iC= -974 
// vC = 14'b1111101000110011; // vC=-1485 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101110; // iC= -978 
// vC = 14'b1111101000111010; // vC=-1478 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001101; // iC= -883 
// vC = 14'b1111100101100100; // vC=-1692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101111; // iC= -721 
// vC = 14'b1111101000010111; // vC=-1513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011100; // iC= -868 
// vC = 14'b1111100111111010; // vC=-1542 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110011; // iC= -845 
// vC = 14'b1111100100111101; // vC=-1731 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011111; // iC= -865 
// vC = 14'b1111100111101011; // vC=-1557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000100; // iC= -764 
// vC = 14'b1111101001010100; // vC=-1452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100001; // iC= -863 
// vC = 14'b1111100101111011; // vC=-1669 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001010; // iC= -822 
// vC = 14'b1111100111110111; // vC=-1545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011111; // iC= -673 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001011; // iC= -693 
// vC = 14'b1111101000000101; // vC=-1531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100010; // iC= -798 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011101; // iC= -867 
// vC = 14'b1111100111101010; // vC=-1558 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101011; // iC= -789 
// vC = 14'b1111100100110111; // vC=-1737 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110111; // iC= -713 
// vC = 14'b1111101000011001; // vC=-1511 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001100; // iC= -820 
// vC = 14'b1111100101000111; // vC=-1721 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101001; // iC= -727 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100001; // iC= -671 
// vC = 14'b1111100101000011; // vC=-1725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011110; // iC= -802 
// vC = 14'b1111100100100000; // vC=-1760 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010110; // iC= -682 
// vC = 14'b1111100110011100; // vC=-1636 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100101; // iC= -667 
// vC = 14'b1111100110110100; // vC=-1612 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101011; // iC= -789 
// vC = 14'b1111100110110011; // vC=-1613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100101; // iC= -603 
// vC = 14'b1111100110110101; // vC=-1611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010011; // iC= -621 
// vC = 14'b1111100110011001; // vC=-1639 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100100; // iC= -732 
// vC = 14'b1111100110010010; // vC=-1646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001101; // iC= -691 
// vC = 14'b1111100011101001; // vC=-1815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100110; // iC= -538 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011100; // iC= -676 
// vC = 14'b1111100101011111; // vC=-1697 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001110; // iC= -626 
// vC = 14'b1111100100111100; // vC=-1732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101111; // iC= -721 
// vC = 14'b1111101000001111; // vC=-1521 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100011; // iC= -797 
// vC = 14'b1111100100000110; // vC=-1786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100111; // iC= -793 
// vC = 14'b1111100100000011; // vC=-1789 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100101; // iC= -603 
// vC = 14'b1111100111001000; // vC=-1592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111000; // iC= -648 
// vC = 14'b1111101000010000; // vC=-1520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011000; // iC= -616 
// vC = 14'b1111100011100000; // vC=-1824 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111001; // iC= -711 
// vC = 14'b1111100111010010; // vC=-1582 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001011; // iC= -629 
// vC = 14'b1111100011011110; // vC=-1826 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011011; // iC= -549 
// vC = 14'b1111100100010011; // vC=-1773 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000000; // iC= -704 
// vC = 14'b1111100100000011; // vC=-1789 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011101; // iC= -739 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011011; // iC= -677 
// vC = 14'b1111100101110111; // vC=-1673 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011011; // iC= -677 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110100; // iC= -652 
// vC = 14'b1111100111101111; // vC=-1553 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100011; // iC= -541 
// vC = 14'b1111100010111011; // vC=-1861 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000000000; // iC= -512 
// vC = 14'b1111100101111000; // vC=-1672 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010010; // iC= -494 
// vC = 14'b1111100111001101; // vC=-1587 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010100; // iC= -684 
// vC = 14'b1111100111100101; // vC=-1563 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110001; // iC= -655 
// vC = 14'b1111100011101000; // vC=-1816 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010001; // iC= -623 
// vC = 14'b1111100011001111; // vC=-1841 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101011; // iC= -469 
// vC = 14'b1111100101011010; // vC=-1702 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000110; // iC= -442 
// vC = 14'b1111100110010010; // vC=-1646 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000101; // iC= -635 
// vC = 14'b1111100110010101; // vC=-1643 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101101; // iC= -531 
// vC = 14'b1111100110111001; // vC=-1607 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000000010; // iC= -510 
// vC = 14'b1111100100111010; // vC=-1734 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010010; // iC= -494 
// vC = 14'b1111100110000000; // vC=-1664 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111111; // iC= -513 
// vC = 14'b1111100011100000; // vC=-1824 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001111; // iC= -625 
// vC = 14'b1111100101000100; // vC=-1724 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111000; // iC= -328 
// vC = 14'b1111100011110111; // vC=-1801 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100100; // iC= -540 
// vC = 14'b1111100110101011; // vC=-1621 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011110; // iC= -546 
// vC = 14'b1111100010101111; // vC=-1873 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111110; // iC= -386 
// vC = 14'b1111100010110000; // vC=-1872 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010010; // iC= -302 
// vC = 14'b1111100011011100; // vC=-1828 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111110011; // iC= -525 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010010; // iC= -366 
// vC = 14'b1111100100011011; // vC=-1765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111100; // iC= -452 
// vC = 14'b1111100100111011; // vC=-1733 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000100; // iC= -252 
// vC = 14'b1111100101011100; // vC=-1700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011100100; // iC= -284 
// vC = 14'b1111100010101011; // vC=-1877 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010010; // iC= -494 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101111; // iC= -273 
// vC = 14'b1111100011100000; // vC=-1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111100; // iC= -196 
// vC = 14'b1111100100111010; // vC=-1734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101000; // iC= -216 
// vC = 14'b1111100100101010; // vC=-1750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010101; // iC= -427 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011100; // iC= -292 
// vC = 14'b1111100011100101; // vC=-1819 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010101; // iC= -171 
// vC = 14'b1111100010100100; // vC=-1884 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110111; // iC= -393 
// vC = 14'b1111100010010111; // vC=-1897 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100111; // iC= -345 
// vC = 14'b1111100011101001; // vC=-1815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111011000; // iC=  -40 
// vC = 14'b1111100010110010; // vC=-1870 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101110011; // iC= -141 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110110001; // iC=  -79 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100101; // iC=  -27 
// vC = 14'b1111100010000011; // vC=-1917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111111; // iC=   -1 
// vC = 14'b1111100110101101; // vC=-1619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111001; // iC=   -7 
// vC = 14'b1111100010111000; // vC=-1864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011000; // iC= -232 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111001; // iC=   -7 
// vC = 14'b1111100110010110; // vC=-1642 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111101; // iC= -131 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001101; // iC=   77 
// vC = 14'b1111100011000100; // vC=-1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010110; // iC= -106 
// vC = 14'b1111100101000000; // vC=-1728 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100000; // iC= -160 
// vC = 14'b1111100010000100; // vC=-1916 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010101; // iC=   21 
// vC = 14'b1111100101101110; // vC=-1682 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010100; // iC= -108 
// vC = 14'b1111100110101110; // vC=-1618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100100; // iC=  228 
// vC = 14'b1111100110011011; // vC=-1637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100010; // iC=   34 
// vC = 14'b1111100100100001; // vC=-1759 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101001; // iC=  105 
// vC = 14'b1111100101101100; // vC=-1684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111001; // iC=  249 
// vC = 14'b1111100100011110; // vC=-1762 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010101; // iC=   21 
// vC = 14'b1111100110010100; // vC=-1644 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100100; // iC=  292 
// vC = 14'b1111100101001111; // vC=-1713 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011111; // iC=   95 
// vC = 14'b1111100101011010; // vC=-1702 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110101; // iC=  181 
// vC = 14'b1111100100001100; // vC=-1780 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001101; // iC=  269 
// vC = 14'b1111100101111111; // vC=-1665 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010101; // iC=  405 
// vC = 14'b1111100101000001; // vC=-1727 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101111; // iC=  367 
// vC = 14'b1111100100001000; // vC=-1784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101011; // iC=  299 
// vC = 14'b1111100101000001; // vC=-1727 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100000; // iC=  288 
// vC = 14'b1111100110000000; // vC=-1664 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110001; // iC=  241 
// vC = 14'b1111100111001000; // vC=-1592 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100001; // iC=  225 
// vC = 14'b1111100111000110; // vC=-1594 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111010; // iC=  570 
// vC = 14'b1111100101100001; // vC=-1695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101011; // iC=  427 
// vC = 14'b1111100010111000; // vC=-1864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111010; // iC=  506 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001000; // iC=  456 
// vC = 14'b1111100101100011; // vC=-1693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011001; // iC=  537 
// vC = 14'b1111100010110000; // vC=-1872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101011; // iC=  619 
// vC = 14'b1111100010110000; // vC=-1872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101011; // iC=  491 
// vC = 14'b1111100100101111; // vC=-1745 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100010; // iC=  610 
// vC = 14'b1111100110011010; // vC=-1638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110010; // iC=  562 
// vC = 14'b1111100100001001; // vC=-1783 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101110; // iC=  686 
// vC = 14'b1111100011101110; // vC=-1810 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010001; // iC=  785 
// vC = 14'b1111100100110010; // vC=-1742 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111010; // iC=  762 
// vC = 14'b1111100101011001; // vC=-1703 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111001; // iC=  825 
// vC = 14'b1111100101110100; // vC=-1676 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011110; // iC=  798 
// vC = 14'b1111100100100100; // vC=-1756 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100101; // iC=  741 
// vC = 14'b1111100111111001; // vC=-1543 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011001; // iC=  665 
// vC = 14'b1111100110101111; // vC=-1617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100010; // iC=  930 
// vC = 14'b1111100110101101; // vC=-1619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110111; // iC=  823 
// vC = 14'b1111100100100000; // vC=-1760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101101; // iC=  877 
// vC = 14'b1111100101011000; // vC=-1704 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011011; // iC=  987 
// vC = 14'b1111100100100010; // vC=-1758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001001; // iC= 1033 
// vC = 14'b1111100110000010; // vC=-1662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010111; // iC=  983 
// vC = 14'b1111100101100000; // vC=-1696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010011; // iC=  787 
// vC = 14'b1111100011100010; // vC=-1822 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100110; // iC=  806 
// vC = 14'b1111101000001001; // vC=-1527 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101111; // iC=  879 
// vC = 14'b1111100111101110; // vC=-1554 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100000; // iC= 1056 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111000; // iC= 1016 
// vC = 14'b1111100110000010; // vC=-1662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101101; // iC=  941 
// vC = 14'b1111100111010011; // vC=-1581 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011100; // iC= 1052 
// vC = 14'b1111100110111010; // vC=-1606 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110001; // iC=  945 
// vC = 14'b1111100111111111; // vC=-1537 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100000; // iC=  928 
// vC = 14'b1111100100010001; // vC=-1775 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001101; // iC= 1101 
// vC = 14'b1111100111001101; // vC=-1587 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010110; // iC= 1046 
// vC = 14'b1111101001000101; // vC=-1467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101010; // iC= 1066 
// vC = 14'b1111101000000101; // vC=-1531 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000011; // iC= 1091 
// vC = 14'b1111100110100000; // vC=-1632 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110101; // iC= 1205 
// vC = 14'b1111100110100010; // vC=-1630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001111; // iC= 1295 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100101; // iC= 1061 
// vC = 14'b1111101000101001; // vC=-1495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100111; // iC= 1255 
// vC = 14'b1111101001011010; // vC=-1446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010011; // iC= 1299 
// vC = 14'b1111101000011001; // vC=-1511 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000100; // iC= 1412 
// vC = 14'b1111101001110000; // vC=-1424 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101110; // iC= 1326 
// vC = 14'b1111100110010011; // vC=-1645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111110; // iC= 1342 
// vC = 14'b1111101001010010; // vC=-1454 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010010; // iC= 1298 
// vC = 14'b1111101000100111; // vC=-1497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100011; // iC= 1379 
// vC = 14'b1111100101101111; // vC=-1681 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110100; // iC= 1396 
// vC = 14'b1111101001111110; // vC=-1410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101001; // iC= 1449 
// vC = 14'b1111101000110000; // vC=-1488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110100; // iC= 1396 
// vC = 14'b1111101000100100; // vC=-1500 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100011; // iC= 1507 
// vC = 14'b1111101010100111; // vC=-1369 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110010; // iC= 1266 
// vC = 14'b1111100110011010; // vC=-1638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000101; // iC= 1541 
// vC = 14'b1111100110001110; // vC=-1650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101000; // iC= 1576 
// vC = 14'b1111101001111101; // vC=-1411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011010; // iC= 1370 
// vC = 14'b1111101001100101; // vC=-1435 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000000; // iC= 1408 
// vC = 14'b1111101010010001; // vC=-1391 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110010; // iC= 1394 
// vC = 14'b1111101010111110; // vC=-1346 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100000; // iC= 1568 
// vC = 14'b1111101000000111; // vC=-1529 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010111; // iC= 1623 
// vC = 14'b1111100111011011; // vC=-1573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101000; // iC= 1448 
// vC = 14'b1111101011100110; // vC=-1306 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000100; // iC= 1604 
// vC = 14'b1111101011100111; // vC=-1305 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111111; // iC= 1535 
// vC = 14'b1111101011110001; // vC=-1295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100010; // iC= 1634 
// vC = 14'b1111101011110011; // vC=-1293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110000; // iC= 1456 
// vC = 14'b1111101010110101; // vC=-1355 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100011; // iC= 1635 
// vC = 14'b1111101001011110; // vC=-1442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000011; // iC= 1667 
// vC = 14'b1111101001000010; // vC=-1470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110110; // iC= 1590 
// vC = 14'b1111101000010000; // vC=-1520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110001; // iC= 1777 
// vC = 14'b1111100111111001; // vC=-1543 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111001; // iC= 1593 
// vC = 14'b1111101011111110; // vC=-1282 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101110; // iC= 1646 
// vC = 14'b1111101001000000; // vC=-1472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111011; // iC= 1659 
// vC = 14'b1111101100011100; // vC=-1252 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111100; // iC= 1660 
// vC = 14'b1111101001010110; // vC=-1450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101111; // iC= 1647 
// vC = 14'b1111101000110110; // vC=-1482 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010111; // iC= 1687 
// vC = 14'b1111101000101111; // vC=-1489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100100; // iC= 1636 
// vC = 14'b1111101100110000; // vC=-1232 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010001; // iC= 1617 
// vC = 14'b1111101101010011; // vC=-1197 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001010; // iC= 1802 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000111; // iC= 1735 
// vC = 14'b1111101100001110; // vC=-1266 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100111; // iC= 1703 
// vC = 14'b1111101100001001; // vC=-1271 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001011; // iC= 1867 
// vC = 14'b1111101010001101; // vC=-1395 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011110; // iC= 1630 
// vC = 14'b1111101010111001; // vC=-1351 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b1111101001010010; // vC=-1454 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111010; // iC= 1914 
// vC = 14'b1111101011000011; // vC=-1341 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b1111101110010110; // vC=-1130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110010; // iC= 1650 
// vC = 14'b1111101110001011; // vC=-1141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101110; // iC= 1710 
// vC = 14'b1111101110001001; // vC=-1143 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010101; // iC= 1685 
// vC = 14'b1111101011111111; // vC=-1281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b1111101100011011; // vC=-1253 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010001; // iC= 1681 
// vC = 14'b1111101100101001; // vC=-1239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010100; // iC= 1748 
// vC = 14'b1111101101011001; // vC=-1191 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000010; // iC= 1730 
// vC = 14'b1111101011010111; // vC=-1321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101101; // iC= 1773 
// vC = 14'b1111101100010011; // vC=-1261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111101110010000; // vC=-1136 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100010; // iC= 1698 
// vC = 14'b1111101110111110; // vC=-1090 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001011; // iC= 1803 
// vC = 14'b1111101101011011; // vC=-1189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001010; // iC= 1802 
// vC = 14'b1111101111010010; // vC=-1070 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110001; // iC= 2033 
// vC = 14'b1111101111111100; // vC=-1028 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010010; // iC= 1874 
// vC = 14'b1111101100111000; // vC=-1224 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b1111101111110010; // vC=-1038 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100110; // iC= 2022 
// vC = 14'b1111101111000100; // vC=-1084 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b1111101110100111; // vC=-1113 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010101; // iC= 1877 
// vC = 14'b1111101101011111; // vC=-1185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001001; // iC= 2057 
// vC = 14'b1111110000100101; // vC= -987 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b1111101111111110; // vC=-1026 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b1111110000001000; // vC=-1016 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110011; // iC= 1907 
// vC = 14'b1111110000001111; // vC=-1009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b1111101101100101; // vC=-1179 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001101; // iC= 1869 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111001; // iC= 1785 
// vC = 14'b1111110000111100; // vC= -964 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010001; // iC= 2001 
// vC = 14'b1111101100111101; // vC=-1219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110100; // iC= 2036 
// vC = 14'b1111101111000111; // vC=-1081 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b1111110010000100; // vC= -892 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b1111110001001000; // vC= -952 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110110; // iC= 1782 
// vC = 14'b1111110000110101; // vC= -971 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001100; // iC= 1804 
// vC = 14'b1111101111101001; // vC=-1047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110000; // iC= 1904 
// vC = 14'b1111110000000100; // vC=-1020 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000001; // iC= 1857 
// vC = 14'b1111101110111111; // vC=-1089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000101; // iC= 1989 
// vC = 14'b1111101111000001; // vC=-1087 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b1111110010000000; // vC= -896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110101; // iC= 2037 
// vC = 14'b1111101111010111; // vC=-1065 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b1111101111110001; // vC=-1039 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101011; // iC= 1963 
// vC = 14'b1111110010010001; // vC= -879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b1111110010101010; // vC= -854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110000; // iC= 2032 
// vC = 14'b1111110010001010; // vC= -886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000010; // iC= 1922 
// vC = 14'b1111110001001000; // vC= -952 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101100; // iC= 1900 
// vC = 14'b1111101111011000; // vC=-1064 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100010; // iC= 1954 
// vC = 14'b1111110001000001; // vC= -959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100110; // iC= 2086 
// vC = 14'b1111110001010110; // vC= -938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110110; // iC= 2038 
// vC = 14'b1111110001001111; // vC= -945 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b1111110001011110; // vC= -930 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111110011111000; // vC= -776 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100001; // iC= 2081 
// vC = 14'b1111110001001011; // vC= -949 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b1111110011010011; // vC= -813 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011111; // iC= 2015 
// vC = 14'b1111110100001000; // vC= -760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000000; // iC= 1856 
// vC = 14'b1111110011000000; // vC= -832 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100101; // iC= 1829 
// vC = 14'b1111110010110001; // vC= -847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111010; // iC= 2106 
// vC = 14'b1111110001110111; // vC= -905 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010101; // iC= 2005 
// vC = 14'b1111110001011111; // vC= -929 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011011; // iC= 1819 
// vC = 14'b1111110010101101; // vC= -851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111110100101111; // vC= -721 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000100; // iC= 1796 
// vC = 14'b1111110011001110; // vC= -818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010011; // iC= 2067 
// vC = 14'b1111110101101111; // vC= -657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b1111110110000101; // vC= -635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010110; // iC= 1814 
// vC = 14'b1111110100110010; // vC= -718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000000; // iC= 2048 
// vC = 14'b1111110011101111; // vC= -785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b1111110100110001; // vC= -719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100101; // iC= 1957 
// vC = 14'b1111110011111111; // vC= -769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011110; // iC= 2014 
// vC = 14'b1111110100110001; // vC= -719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b1111110010100001; // vC= -863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b1111110110111001; // vC= -583 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b1111110010110001; // vC= -847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101101; // iC= 1837 
// vC = 14'b1111110100101100; // vC= -724 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111010; // iC= 1914 
// vC = 14'b1111110110010001; // vC= -623 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b1111110100010100; // vC= -748 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011111; // iC= 1823 
// vC = 14'b1111110101100000; // vC= -672 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000101; // iC= 1925 
// vC = 14'b1111110111100010; // vC= -542 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011000; // iC= 1880 
// vC = 14'b1111110100000011; // vC= -765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010110; // iC= 1814 
// vC = 14'b1111110110010001; // vC= -623 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101010; // iC= 1834 
// vC = 14'b1111110110001010; // vC= -630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100110; // iC= 1830 
// vC = 14'b1111110011100101; // vC= -795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110110; // iC= 2038 
// vC = 14'b1111110111010110; // vC= -554 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111110100111110; // vC= -706 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b1111110111100010; // vC= -542 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001001; // iC= 1801 
// vC = 14'b1111110111000000; // vC= -576 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b1111111000000011; // vC= -509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111000; // iC= 2104 
// vC = 14'b1111110110010000; // vC= -624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001101; // iC= 1997 
// vC = 14'b1111110101000101; // vC= -699 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b1111110111001110; // vC= -562 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101001; // iC= 1833 
// vC = 14'b1111111000100100; // vC= -476 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b1111110110101001; // vC= -599 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111011; // iC= 1851 
// vC = 14'b1111110110100111; // vC= -601 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b1111110101011001; // vC= -679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010011; // iC= 1811 
// vC = 14'b1111110111111001; // vC= -519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b1111110111011011; // vC= -549 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001110; // iC= 1934 
// vC = 14'b1111111000110001; // vC= -463 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011101; // iC= 1885 
// vC = 14'b1111110101101010; // vC= -662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100010; // iC= 2018 
// vC = 14'b1111111000101101; // vC= -467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111101; // iC= 2109 
// vC = 14'b1111111001011111; // vC= -417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111111000010000; // vC= -496 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010100; // iC= 1876 
// vC = 14'b1111110110111101; // vC= -579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000101; // iC= 1861 
// vC = 14'b1111110111111100; // vC= -516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b1111110111001001; // vC= -567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010101; // iC= 1813 
// vC = 14'b1111111000100110; // vC= -474 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001100; // iC= 1804 
// vC = 14'b1111110111100001; // vC= -543 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000010; // iC= 2050 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100101; // iC= 1893 
// vC = 14'b1111110111010011; // vC= -557 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011101; // iC= 1821 
// vC = 14'b1111111001110000; // vC= -400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b1111110111011111; // vC= -545 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b1111111000010010; // vC= -494 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101110; // iC= 2030 
// vC = 14'b1111111011000100; // vC= -316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b1111111011111000; // vC= -264 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000101; // iC= 1797 
// vC = 14'b1111111011100001; // vC= -287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b1111111011000101; // vC= -315 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010000; // iC= 1808 
// vC = 14'b1111111100110101; // vC= -203 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001001; // iC= 1801 
// vC = 14'b1111111100000000; // vC= -256 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b1111111100011110; // vC= -226 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000001; // iC= 1793 
// vC = 14'b1111111101000011; // vC= -189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b1111111100010100; // vC= -236 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110011; // iC= 1971 
// vC = 14'b1111111010010001; // vC= -367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111000; // iC= 1976 
// vC = 14'b1111111101000100; // vC= -188 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101111; // iC= 2095 
// vC = 14'b1111111001101010; // vC= -406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000101; // iC= 1989 
// vC = 14'b1111111011011101; // vC= -291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111111101110101; // vC= -139 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000111; // iC= 1799 
// vC = 14'b1111111010011111; // vC= -353 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b1111111100111000; // vC= -200 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b1111111010111100; // vC= -324 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b1111111001111001; // vC= -391 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b1111111101111101; // vC= -131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010000; // iC= 2064 
// vC = 14'b1111111011000001; // vC= -319 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000011; // iC= 1859 
// vC = 14'b1111111011001110; // vC= -306 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111010; // iC= 1850 
// vC = 14'b1111111101100010; // vC= -158 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111010; // iC= 1786 
// vC = 14'b1111111101110011; // vC= -141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010001; // iC= 1809 
// vC = 14'b1111111100011111; // vC= -225 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111111011100111; // vC= -281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b1111111110111000; // vC=  -72 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010001; // iC= 1809 
// vC = 14'b1111111010111111; // vC= -321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111111011101111; // vC= -273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101110; // iC= 1902 
// vC = 14'b1111111101000011; // vC= -189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b1111111111110000; // vC=  -16 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011000; // iC= 1816 
// vC = 14'b1111111110110000; // vC=  -80 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111010; // iC= 1786 
// vC = 14'b1111111101111010; // vC= -134 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100101; // iC= 1893 
// vC = 14'b1111111101000110; // vC= -186 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111110; // iC= 1854 
// vC = 14'b1111111011101011; // vC= -277 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100000; // iC= 1760 
// vC = 14'b0000000000001000; // vC=    8 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b1111111100011010; // vC= -230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010011; // iC= 1875 
// vC = 14'b0000000001001001; // vC=   73 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100000; // iC= 1760 
// vC = 14'b1111111110001101; // vC= -115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010000; // iC= 1808 
// vC = 14'b1111111111000110; // vC=  -58 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110100; // iC= 1780 
// vC = 14'b1111111111010111; // vC=  -41 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001000; // iC= 1928 
// vC = 14'b1111111111110111; // vC=   -9 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b1111111101101111; // vC= -145 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101011; // iC= 1899 
// vC = 14'b1111111100111101; // vC= -195 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010001; // iC= 1745 
// vC = 14'b1111111111110101; // vC=  -11 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010101; // iC= 2005 
// vC = 14'b1111111101100111; // vC= -153 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000101; // iC= 1797 
// vC = 14'b0000000001110101; // vC=  117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110000; // iC= 1968 
// vC = 14'b1111111111101011; // vC=  -21 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111111110100011; // vC=  -93 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b0000000000101000; // vC=   40 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010111; // iC= 1879 
// vC = 14'b0000000001110010; // vC=  114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b0000000010111011; // vC=  187 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b1111111110011101; // vC=  -99 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110100; // iC= 1844 
// vC = 14'b1111111110111100; // vC=  -68 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000100; // iC= 1988 
// vC = 14'b1111111111111011; // vC=   -5 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111101; // iC= 1725 
// vC = 14'b1111111111010111; // vC=  -41 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000101; // iC= 1733 
// vC = 14'b0000000001100011; // vC=   99 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111110; // iC= 1854 
// vC = 14'b0000000010111110; // vC=  190 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101010; // iC= 1770 
// vC = 14'b0000000000100101; // vC=   37 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101010; // iC= 1834 
// vC = 14'b1111111111100000; // vC=  -32 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001110; // iC= 1806 
// vC = 14'b1111111111001001; // vC=  -55 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101100; // iC= 1708 
// vC = 14'b0000000011001001; // vC=  201 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b1111111111011010; // vC=  -38 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b1111111111100010; // vC=  -30 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b0000000000011010; // vC=   26 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101100; // iC= 1708 
// vC = 14'b0000000011111111; // vC=  255 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110110; // iC= 1718 
// vC = 14'b0000000011011011; // vC=  219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b0000000010011000; // vC=  152 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b0000000001000101; // vC=   69 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101101; // iC= 1837 
// vC = 14'b0000000011010101; // vC=  213 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111001; // iC= 1849 
// vC = 14'b0000000010010100; // vC=  148 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100101; // iC= 1893 
// vC = 14'b0000000010101110; // vC=  174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011100; // iC= 1948 
// vC = 14'b0000000101011011; // vC=  347 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b0000000010111111; // vC=  191 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110101; // iC= 1845 
// vC = 14'b0000000011100111; // vC=  231 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b0000000011001111; // vC=  207 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010100; // iC= 1684 
// vC = 14'b0000000001111000; // vC=  120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011100; // iC= 1820 
// vC = 14'b0000000100010110; // vC=  278 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000110; // iC= 1862 
// vC = 14'b0000000100111110; // vC=  318 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b0000000011111000; // vC=  248 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001010; // iC= 1738 
// vC = 14'b0000000011010010; // vC=  210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b0000000011110111; // vC=  247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000000; // iC= 1728 
// vC = 14'b0000000110010110; // vC=  406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011111; // iC= 1887 
// vC = 14'b0000000100111101; // vC=  317 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100100; // iC= 1764 
// vC = 14'b0000000011010111; // vC=  215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b0000000110101000; // vC=  424 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b0000000100100001; // vC=  289 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b0000000010111101; // vC=  189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011101; // iC= 1885 
// vC = 14'b0000000110100101; // vC=  421 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b0000000011000011; // vC=  195 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000001; // iC= 1729 
// vC = 14'b0000000011111010; // vC=  250 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001010; // iC= 1866 
// vC = 14'b0000001000000000; // vC=  512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010110; // iC= 1878 
// vC = 14'b0000000110111010; // vC=  442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111000; // iC= 1656 
// vC = 14'b0000000110101101; // vC=  429 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011001; // iC= 1689 
// vC = 14'b0000000011011100; // vC=  220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101011; // iC= 1899 
// vC = 14'b0000000111110111; // vC=  503 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000010; // iC= 1730 
// vC = 14'b0000001000010010; // vC=  530 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100001; // iC= 1761 
// vC = 14'b0000001000000001; // vC=  513 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101100; // iC= 1772 
// vC = 14'b0000000011111000; // vC=  248 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000001; // iC= 1729 
// vC = 14'b0000000011110111; // vC=  247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110100; // iC= 1716 
// vC = 14'b0000000100000110; // vC=  262 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110100; // iC= 1652 
// vC = 14'b0000000100011000; // vC=  280 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101010; // iC= 1834 
// vC = 14'b0000001000110011; // vC=  563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b0000000110111100; // vC=  444 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100100; // iC= 1700 
// vC = 14'b0000000111101101; // vC=  493 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100101; // iC= 1637 
// vC = 14'b0000000101001101; // vC=  333 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000110; // iC= 1670 
// vC = 14'b0000001001101110; // vC=  622 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010100; // iC= 1748 
// vC = 14'b0000000110101110; // vC=  430 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100011; // iC= 1763 
// vC = 14'b0000000111001011; // vC=  459 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111101; // iC= 1597 
// vC = 14'b0000000111111011; // vC=  507 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100101; // iC= 1893 
// vC = 14'b0000000110000001; // vC=  385 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010011; // iC= 1811 
// vC = 14'b0000000111101011; // vC=  491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b0000000101111101; // vC=  381 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111111; // iC= 1663 
// vC = 14'b0000000111001111; // vC=  463 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011001; // iC= 1817 
// vC = 14'b0000001000110111; // vC=  567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111010; // iC= 1658 
// vC = 14'b0000000111011000; // vC=  472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101000; // iC= 1768 
// vC = 14'b0000001001010100; // vC=  596 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b0000001010100110; // vC=  678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101001; // iC= 1705 
// vC = 14'b0000000111010110; // vC=  470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011010; // iC= 1754 
// vC = 14'b0000000110011110; // vC=  414 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110111; // iC= 1591 
// vC = 14'b0000001001001100; // vC=  588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000001; // iC= 1857 
// vC = 14'b0000000110101101; // vC=  429 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001111; // iC= 1679 
// vC = 14'b0000001000111001; // vC=  569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100110; // iC= 1702 
// vC = 14'b0000001010000001; // vC=  641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b0000000111100101; // vC=  485 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101101; // iC= 1773 
// vC = 14'b0000001000110011; // vC=  563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111010; // iC= 1658 
// vC = 14'b0000001000101100; // vC=  556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110101; // iC= 1717 
// vC = 14'b0000001001101001; // vC=  617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001011; // iC= 1675 
// vC = 14'b0000001000001110; // vC=  526 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010100; // iC= 1556 
// vC = 14'b0000001001001100; // vC=  588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000011; // iC= 1667 
// vC = 14'b0000001000100111; // vC=  551 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000110; // iC= 1798 
// vC = 14'b0000000111111100; // vC=  508 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010010; // iC= 1618 
// vC = 14'b0000001011101111; // vC=  751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110110; // iC= 1782 
// vC = 14'b0000001100110110; // vC=  822 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010111; // iC= 1815 
// vC = 14'b0000001011101111; // vC=  751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110110; // iC= 1718 
// vC = 14'b0000001000010001; // vC=  529 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110110; // iC= 1718 
// vC = 14'b0000001011001111; // vC=  719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101000; // iC= 1512 
// vC = 14'b0000001011110100; // vC=  756 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011100; // iC= 1756 
// vC = 14'b0000001001111001; // vC=  633 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001111; // iC= 1551 
// vC = 14'b0000001011011111; // vC=  735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001001; // iC= 1545 
// vC = 14'b0000001001001110; // vC=  590 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010111; // iC= 1687 
// vC = 14'b0000001001001110; // vC=  590 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000010; // iC= 1794 
// vC = 14'b0000001010010011; // vC=  659 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001010; // iC= 1674 
// vC = 14'b0000001001011100; // vC=  604 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010101; // iC= 1621 
// vC = 14'b0000001001110001; // vC=  625 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010100; // iC= 1684 
// vC = 14'b0000001010110010; // vC=  690 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011110; // iC= 1694 
// vC = 14'b0000001100010010; // vC=  786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101101; // iC= 1517 
// vC = 14'b0000001101010010; // vC=  850 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010100; // iC= 1556 
// vC = 14'b0000001100100010; // vC=  802 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110001; // iC= 1521 
// vC = 14'b0000001101001000; // vC=  840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100001; // iC= 1505 
// vC = 14'b0000001010011110; // vC=  670 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011011; // iC= 1691 
// vC = 14'b0000001001111010; // vC=  634 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110100; // iC= 1524 
// vC = 14'b0000001100001001; // vC=  777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111000; // iC= 1720 
// vC = 14'b0000001101010011; // vC=  851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001011; // iC= 1739 
// vC = 14'b0000001111000010; // vC=  962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001000; // iC= 1672 
// vC = 14'b0000001101101110; // vC=  878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100000; // iC= 1696 
// vC = 14'b0000001101010010; // vC=  850 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110011; // iC= 1523 
// vC = 14'b0000001101011000; // vC=  856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110000; // iC= 1712 
// vC = 14'b0000001011000001; // vC=  705 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000000; // iC= 1536 
// vC = 14'b0000001011101011; // vC=  747 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001011; // iC= 1483 
// vC = 14'b0000001101101111; // vC=  879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110111; // iC= 1591 
// vC = 14'b0000001110000001; // vC=  897 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010001; // iC= 1681 
// vC = 14'b0000001101101111; // vC=  879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010101; // iC= 1621 
// vC = 14'b0000001111101110; // vC= 1006 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100110; // iC= 1510 
// vC = 14'b0000001110111011; // vC=  955 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100110; // iC= 1446 
// vC = 14'b0000001011011111; // vC=  735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001001; // iC= 1417 
// vC = 14'b0000001100100111; // vC=  807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100010; // iC= 1378 
// vC = 14'b0000010000011001; // vC= 1049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011101; // iC= 1501 
// vC = 14'b0000001101100001; // vC=  865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100001; // iC= 1505 
// vC = 14'b0000010000011101; // vC= 1053 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011110; // iC= 1630 
// vC = 14'b0000001101101111; // vC=  879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011100; // iC= 1436 
// vC = 14'b0000001111010001; // vC=  977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000011; // iC= 1667 
// vC = 14'b0000001100000010; // vC=  770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101110; // iC= 1390 
// vC = 14'b0000001101001001; // vC=  841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100011; // iC= 1571 
// vC = 14'b0000001100010011; // vC=  787 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000101; // iC= 1413 
// vC = 14'b0000001110001101; // vC=  909 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001100; // iC= 1484 
// vC = 14'b0000001111000011; // vC=  963 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110011; // iC= 1651 
// vC = 14'b0000001111010011; // vC=  979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111111; // iC= 1599 
// vC = 14'b0000010000000101; // vC= 1029 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001110; // iC= 1358 
// vC = 14'b0000001101011001; // vC=  857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110000; // iC= 1520 
// vC = 14'b0000010000010111; // vC= 1047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001011; // iC= 1355 
// vC = 14'b0000010001010001; // vC= 1105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101100; // iC= 1452 
// vC = 14'b0000001110110001; // vC=  945 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111110; // iC= 1342 
// vC = 14'b0000001110111000; // vC=  952 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010000; // iC= 1424 
// vC = 14'b0000001101111001; // vC=  889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001001; // iC= 1609 
// vC = 14'b0000001111000101; // vC=  965 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011011; // iC= 1499 
// vC = 14'b0000001110110110; // vC=  950 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010010; // iC= 1426 
// vC = 14'b0000010010001011; // vC= 1163 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001100; // iC= 1356 
// vC = 14'b0000001101101000; // vC=  872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011110; // iC= 1502 
// vC = 14'b0000001110111010; // vC=  954 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101110; // iC= 1518 
// vC = 14'b0000001110100100; // vC=  932 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000111; // iC= 1287 
// vC = 14'b0000001110110101; // vC=  949 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111010; // iC= 1530 
// vC = 14'b0000001110101101; // vC=  941 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100110; // iC= 1510 
// vC = 14'b0000010000011101; // vC= 1053 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011100; // iC= 1308 
// vC = 14'b0000010010100010; // vC= 1186 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000011; // iC= 1411 
// vC = 14'b0000001110111110; // vC=  958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101101; // iC= 1517 
// vC = 14'b0000001111001101; // vC=  973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001101; // iC= 1549 
// vC = 14'b0000010010100000; // vC= 1184 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000101; // iC= 1349 
// vC = 14'b0000001110110110; // vC=  950 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100000; // iC= 1568 
// vC = 14'b0000001110111110; // vC=  958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011001; // iC= 1433 
// vC = 14'b0000001111001000; // vC=  968 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010011; // iC= 1491 
// vC = 14'b0000010011000100; // vC= 1220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000110; // iC= 1350 
// vC = 14'b0000010010010000; // vC= 1168 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011010; // iC= 1370 
// vC = 14'b0000001111010110; // vC=  982 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111111; // iC= 1279 
// vC = 14'b0000010011001111; // vC= 1231 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101101; // iC= 1517 
// vC = 14'b0000010001111000; // vC= 1144 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000110; // iC= 1286 
// vC = 14'b0000010001001010; // vC= 1098 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110101; // iC= 1525 
// vC = 14'b0000010001100100; // vC= 1124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110011; // iC= 1267 
// vC = 14'b0000001111011001; // vC=  985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011001; // iC= 1497 
// vC = 14'b0000010011101010; // vC= 1258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111101; // iC= 1341 
// vC = 14'b0000010011010100; // vC= 1236 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100110; // iC= 1382 
// vC = 14'b0000001111101110; // vC= 1006 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100110; // iC= 1446 
// vC = 14'b0000010001000001; // vC= 1089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101110; // iC= 1198 
// vC = 14'b0000010010111011; // vC= 1211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111001; // iC= 1337 
// vC = 14'b0000010001001100; // vC= 1100 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101110; // iC= 1262 
// vC = 14'b0000010001011101; // vC= 1117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011010; // iC= 1306 
// vC = 14'b0000010000000010; // vC= 1026 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001001; // iC= 1289 
// vC = 14'b0000010100011110; // vC= 1310 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110010; // iC= 1330 
// vC = 14'b0000010100011101; // vC= 1309 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000110; // iC= 1222 
// vC = 14'b0000010100000110; // vC= 1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001010; // iC= 1162 
// vC = 14'b0000010100101101; // vC= 1325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000110; // iC= 1350 
// vC = 14'b0000010010111000; // vC= 1208 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001000; // iC= 1352 
// vC = 14'b0000010011001001; // vC= 1225 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100111; // iC= 1255 
// vC = 14'b0000010011101010; // vC= 1258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111000; // iC= 1336 
// vC = 14'b0000010010010110; // vC= 1174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101001; // iC= 1385 
// vC = 14'b0000010001100010; // vC= 1122 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001111; // iC= 1231 
// vC = 14'b0000010001111010; // vC= 1146 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100100; // iC= 1252 
// vC = 14'b0000010101000010; // vC= 1346 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101111; // iC= 1391 
// vC = 14'b0000010010110110; // vC= 1206 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101010; // iC= 1386 
// vC = 14'b0000010011000001; // vC= 1217 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010011; // iC= 1235 
// vC = 14'b0000010011111101; // vC= 1277 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000100; // iC= 1092 
// vC = 14'b0000010001100101; // vC= 1125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111101; // iC= 1341 
// vC = 14'b0000010010101011; // vC= 1195 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000110; // iC= 1222 
// vC = 14'b0000010110010110; // vC= 1430 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000101; // iC= 1349 
// vC = 14'b0000010001101011; // vC= 1131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011010; // iC= 1242 
// vC = 14'b0000010010011111; // vC= 1183 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110111; // iC= 1271 
// vC = 14'b0000010011011110; // vC= 1246 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110100; // iC= 1268 
// vC = 14'b0000010011010100; // vC= 1236 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110000; // iC= 1200 
// vC = 14'b0000010001110001; // vC= 1137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011110; // iC= 1374 
// vC = 14'b0000010010010001; // vC= 1169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000100; // iC= 1284 
// vC = 14'b0000010100001110; // vC= 1294 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101001; // iC= 1129 
// vC = 14'b0000010100110000; // vC= 1328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111001; // iC= 1337 
// vC = 14'b0000010011000101; // vC= 1221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011101; // iC= 1309 
// vC = 14'b0000010011101100; // vC= 1260 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111011; // iC= 1147 
// vC = 14'b0000010100001101; // vC= 1293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001000; // iC= 1160 
// vC = 14'b0000010011100111; // vC= 1255 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100010; // iC= 1250 
// vC = 14'b0000010110100101; // vC= 1445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011001; // iC= 1049 
// vC = 14'b0000010101111110; // vC= 1406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101000; // iC= 1064 
// vC = 14'b0000010110001000; // vC= 1416 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011000; // iC= 1304 
// vC = 14'b0000010110111011; // vC= 1467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001100; // iC= 1228 
// vC = 14'b0000010111001011; // vC= 1483 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100100; // iC= 1188 
// vC = 14'b0000010100111011; // vC= 1339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111100; // iC= 1084 
// vC = 14'b0000010011000011; // vC= 1219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011001; // iC=  985 
// vC = 14'b0000010110001010; // vC= 1418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111001; // iC= 1209 
// vC = 14'b0000010110100101; // vC= 1445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011111; // iC= 1119 
// vC = 14'b0000010101111010; // vC= 1402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111101; // iC= 1277 
// vC = 14'b0000010111101000; // vC= 1512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010110; // iC= 1110 
// vC = 14'b0000011000001010; // vC= 1546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101100; // iC= 1196 
// vC = 14'b0000010110100101; // vC= 1445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101001; // iC= 1257 
// vC = 14'b0000010100011110; // vC= 1310 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010010; // iC= 1106 
// vC = 14'b0000010101001000; // vC= 1352 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101011; // iC= 1131 
// vC = 14'b0000010111011001; // vC= 1497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101001; // iC= 1129 
// vC = 14'b0000010111100000; // vC= 1504 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010101; // iC= 1173 
// vC = 14'b0000010100100011; // vC= 1315 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010000; // iC= 1104 
// vC = 14'b0000010011101010; // vC= 1258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001011; // iC= 1227 
// vC = 14'b0000011000101011; // vC= 1579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000110; // iC= 1030 
// vC = 14'b0000010111001101; // vC= 1485 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111100; // iC= 1020 
// vC = 14'b0000010110000000; // vC= 1408 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111111; // iC= 1023 
// vC = 14'b0000010011111011; // vC= 1275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011010; // iC= 1050 
// vC = 14'b0000010111001010; // vC= 1482 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101100; // iC= 1196 
// vC = 14'b0000010111001100; // vC= 1484 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010100; // iC= 1108 
// vC = 14'b0000010110000111; // vC= 1415 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010000; // iC= 1168 
// vC = 14'b0000011000010011; // vC= 1555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001100; // iC=  908 
// vC = 14'b0000010101011000; // vC= 1368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101101; // iC= 1069 
// vC = 14'b0000010100110001; // vC= 1329 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110001; // iC= 1009 
// vC = 14'b0000010101111001; // vC= 1401 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101010; // iC= 1066 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101101; // iC=  877 
// vC = 14'b0000011000010110; // vC= 1558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000110; // iC= 1158 
// vC = 14'b0000010101001101; // vC= 1357 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100001; // iC=  929 
// vC = 14'b0000010111010101; // vC= 1493 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110111; // iC= 1143 
// vC = 14'b0000011000110000; // vC= 1584 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011101; // iC=  861 
// vC = 14'b0000010101110001; // vC= 1393 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010111; // iC=  983 
// vC = 14'b0000011000111101; // vC= 1597 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010011; // iC=  851 
// vC = 14'b0000011001010001; // vC= 1617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111100; // iC=  892 
// vC = 14'b0000011000101100; // vC= 1580 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101111; // iC=  879 
// vC = 14'b0000010101001100; // vC= 1356 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000010; // iC=  962 
// vC = 14'b0000010101111100; // vC= 1404 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100111; // iC=  935 
// vC = 14'b0000011000011111; // vC= 1567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101001; // iC=  873 
// vC = 14'b0000010110011001; // vC= 1433 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100110; // iC=  934 
// vC = 14'b0000011001111111; // vC= 1663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000101; // iC=  901 
// vC = 14'b0000011010010010; // vC= 1682 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001000; // iC= 1032 
// vC = 14'b0000011000101101; // vC= 1581 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010110; // iC=  918 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100101; // iC= 1061 
// vC = 14'b0000010111011011; // vC= 1499 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011000; // iC=  984 
// vC = 14'b0000011000100111; // vC= 1575 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011000; // iC=  792 
// vC = 14'b0000011010000010; // vC= 1666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010100; // iC=  980 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110000; // iC= 1008 
// vC = 14'b0000011001001101; // vC= 1613 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111010; // iC=  826 
// vC = 14'b0000011001001001; // vC= 1609 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000010; // iC=  770 
// vC = 14'b0000011010010111; // vC= 1687 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110000; // iC=  944 
// vC = 14'b0000010110010001; // vC= 1425 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000000; // iC=  896 
// vC = 14'b0000011010110110; // vC= 1718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110000; // iC=  880 
// vC = 14'b0000011001001101; // vC= 1613 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011011; // iC=  923 
// vC = 14'b0000010110110000; // vC= 1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001000; // iC=  904 
// vC = 14'b0000011000000110; // vC= 1542 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001011; // iC=  971 
// vC = 14'b0000010111100100; // vC= 1508 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111111; // iC=  703 
// vC = 14'b0000010110101011; // vC= 1451 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010001; // iC=  785 
// vC = 14'b0000011000011111; // vC= 1567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110010; // iC=  690 
// vC = 14'b0000011000010001; // vC= 1553 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001000; // iC=  712 
// vC = 14'b0000011011000110; // vC= 1734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000011; // iC=  899 
// vC = 14'b0000010111011010; // vC= 1498 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110010; // iC=  754 
// vC = 14'b0000011000010110; // vC= 1558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001011; // iC=  779 
// vC = 14'b0000011011100000; // vC= 1760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001110; // iC=  910 
// vC = 14'b0000010111011111; // vC= 1503 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111110; // iC=  766 
// vC = 14'b0000010111010111; // vC= 1495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001011; // iC=  843 
// vC = 14'b0000011000010111; // vC= 1559 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101001; // iC=  809 
// vC = 14'b0000010111010110; // vC= 1494 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101001; // iC=  873 
// vC = 14'b0000011001110101; // vC= 1653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101010; // iC=  682 
// vC = 14'b0000011001010101; // vC= 1621 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010101; // iC=  789 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110001; // iC=  753 
// vC = 14'b0000011010001111; // vC= 1679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001101; // iC=  653 
// vC = 14'b0000011001111111; // vC= 1663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111011; // iC=  827 
// vC = 14'b0000011000011000; // vC= 1560 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100110; // iC=  614 
// vC = 14'b0000011001011011; // vC= 1627 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111110; // iC=  702 
// vC = 14'b0000010111111010; // vC= 1530 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000101; // iC=  773 
// vC = 14'b0000011001100011; // vC= 1635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001100; // iC=  780 
// vC = 14'b0000011011111011; // vC= 1787 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111111; // iC=  767 
// vC = 14'b0000011001001111; // vC= 1615 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101010; // iC=  746 
// vC = 14'b0000011011100001; // vC= 1761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001111; // iC=  591 
// vC = 14'b0000010111100010; // vC= 1506 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011111; // iC=  543 
// vC = 14'b0000011100011000; // vC= 1816 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b0000011011010101; // vC= 1749 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100101; // iC=  741 
// vC = 14'b0000011011011000; // vC= 1752 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010001; // iC=  785 
// vC = 14'b0000011011000010; // vC= 1730 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000010; // iC=  642 
// vC = 14'b0000010111110100; // vC= 1524 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101011; // iC=  811 
// vC = 14'b0000011011001110; // vC= 1742 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011110; // iC=  606 
// vC = 14'b0000011011011000; // vC= 1752 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000101; // iC=  773 
// vC = 14'b0000011010001011; // vC= 1675 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001101; // iC=  781 
// vC = 14'b0000011010101000; // vC= 1704 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001000; // iC=  584 
// vC = 14'b0000011011101010; // vC= 1770 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000111; // iC=  711 
// vC = 14'b0000011011000111; // vC= 1735 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100101; // iC=  805 
// vC = 14'b0000011010001111; // vC= 1679 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010000; // iC=  592 
// vC = 14'b0000011010111100; // vC= 1724 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100100; // iC=  676 
// vC = 14'b0000011100111101; // vC= 1853 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000110; // iC=  646 
// vC = 14'b0000011010110110; // vC= 1718 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011101; // iC=  733 
// vC = 14'b0000011010010000; // vC= 1680 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000011; // iC=  771 
// vC = 14'b0000011011000011; // vC= 1731 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000000; // iC=  512 
// vC = 14'b0000011101000110; // vC= 1862 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111100; // iC=  444 
// vC = 14'b0000011001111101; // vC= 1661 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011000; // iC=  600 
// vC = 14'b0000011100100110; // vC= 1830 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101100; // iC=  556 
// vC = 14'b0000011100101000; // vC= 1832 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010000; // iC=  720 
// vC = 14'b0000011011100101; // vC= 1765 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011100; // iC=  668 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011011; // iC=  411 
// vC = 14'b0000011101001010; // vC= 1866 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110010; // iC=  562 
// vC = 14'b0000011011001011; // vC= 1739 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111010; // iC=  378 
// vC = 14'b0000011000111110; // vC= 1598 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011100; // iC=  668 
// vC = 14'b0000011100010110; // vC= 1814 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100011; // iC=  419 
// vC = 14'b0000011010101100; // vC= 1708 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100110; // iC=  486 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111100; // iC=  572 
// vC = 14'b0000011010100111; // vC= 1703 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000010; // iC=  514 
// vC = 14'b0000011011010111; // vC= 1751 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100001; // iC=  481 
// vC = 14'b0000011101000000; // vC= 1856 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011001; // iC=  281 
// vC = 14'b0000011101100010; // vC= 1890 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101011; // iC=  363 
// vC = 14'b0000011100000110; // vC= 1798 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001100; // iC=  396 
// vC = 14'b0000011011110011; // vC= 1779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101010; // iC=  490 
// vC = 14'b0000011011011011; // vC= 1755 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110101; // iC=  373 
// vC = 14'b0000011010000101; // vC= 1669 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100011; // iC=  419 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101110; // iC=  302 
// vC = 14'b0000011101010100; // vC= 1876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001001; // iC=  329 
// vC = 14'b0000011000111000; // vC= 1592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110011; // iC=  435 
// vC = 14'b0000011100000110; // vC= 1798 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010000; // iC=  144 
// vC = 14'b0000011001111110; // vC= 1662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110100; // iC=  372 
// vC = 14'b0000011001010000; // vC= 1616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000100; // iC=  260 
// vC = 14'b0000011100100111; // vC= 1831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001010; // iC=  394 
// vC = 14'b0000011101000100; // vC= 1860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101111; // iC=  175 
// vC = 14'b0000011100011011; // vC= 1819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011000; // iC=  280 
// vC = 14'b0000011010001111; // vC= 1679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010010; // iC=  338 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101001; // iC=  297 
// vC = 14'b0000011010110001; // vC= 1713 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011101; // iC=   93 
// vC = 14'b0000011010100100; // vC= 1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010010; // iC=  274 
// vC = 14'b0000011011000101; // vC= 1733 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110000; // iC=  176 
// vC = 14'b0000011100111001; // vC= 1849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100011; // iC=   99 
// vC = 14'b0000011101011011; // vC= 1883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001101; // iC=   77 
// vC = 14'b0000011101010001; // vC= 1873 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111010; // iC=  -70 
// vC = 14'b0000011010000111; // vC= 1671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011010; // iC=   26 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011111; // iC=   31 
// vC = 14'b0000011011010100; // vC= 1748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101111; // iC=  -17 
// vC = 14'b0000011011110000; // vC= 1776 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001000011; // iC=   67 
// vC = 14'b0000011001001000; // vC= 1608 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011101; // iC=   29 
// vC = 14'b0000011011110010; // vC= 1778 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111100; // iC= -132 
// vC = 14'b0000011010101110; // vC= 1710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010100; // iC=   84 
// vC = 14'b0000011100110101; // vC= 1845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100001; // iC=   33 
// vC = 14'b0000011001100101; // vC= 1637 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100000; // iC= -224 
// vC = 14'b0000011010100111; // vC= 1703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000110; // iC= -250 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101001; // iC= -215 
// vC = 14'b0000011101000110; // vC= 1862 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010100; // iC= -236 
// vC = 14'b0000011001001100; // vC= 1612 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001011; // iC= -181 
// vC = 14'b0000011100001010; // vC= 1802 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011010; // iC= -358 
// vC = 14'b0000011001001111; // vC= 1615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101011010; // iC= -166 
// vC = 14'b0000011100100001; // vC= 1825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100100; // iC= -220 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010011; // iC= -237 
// vC = 14'b0000011101011100; // vC= 1884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010010; // iC= -430 
// vC = 14'b0000011001101000; // vC= 1640 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001101; // iC= -307 
// vC = 14'b0000011100001001; // vC= 1801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001100; // iC= -500 
// vC = 14'b0000011001110110; // vC= 1654 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001100; // iC= -308 
// vC = 14'b0000011010111011; // vC= 1723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101100; // iC= -404 
// vC = 14'b0000011100100010; // vC= 1826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010000; // iC= -432 
// vC = 14'b0000011011010100; // vC= 1748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111101; // iC= -451 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111010; // iC= -326 
// vC = 14'b0000011001000100; // vC= 1604 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111011; // iC= -517 
// vC = 14'b0000011001011100; // vC= 1628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010010; // iC= -430 
// vC = 14'b0000011000110001; // vC= 1585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000110; // iC= -698 
// vC = 14'b0000011100000000; // vC= 1792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001001; // iC= -631 
// vC = 14'b0000011100111010; // vC= 1850 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111100; // iC= -580 
// vC = 14'b0000011010111111; // vC= 1727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111001; // iC= -583 
// vC = 14'b0000011001011110; // vC= 1630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111000; // iC= -520 
// vC = 14'b0000011100101101; // vC= 1837 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001110; // iC= -562 
// vC = 14'b0000011010111000; // vC= 1720 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111000; // iC= -712 
// vC = 14'b0000011010101101; // vC= 1709 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001000; // iC= -696 
// vC = 14'b0000011010011110; // vC= 1694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011000; // iC= -872 
// vC = 14'b0000011011011110; // vC= 1758 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101110; // iC= -786 
// vC = 14'b0000011001001111; // vC= 1615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000000; // iC= -896 
// vC = 14'b0000011001000011; // vC= 1603 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001010; // iC= -822 
// vC = 14'b0000011001101100; // vC= 1644 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100110; // iC= -922 
// vC = 14'b0000011000001111; // vC= 1551 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100101; // iC= -859 
// vC = 14'b0000011000000011; // vC= 1539 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010101; // iC= -747 
// vC = 14'b0000011000110100; // vC= 1588 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010001; // iC= -751 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011111; // iC= -929 
// vC = 14'b0000011010111111; // vC= 1727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101011; // iC=-1045 
// vC = 14'b0000011011011000; // vC= 1752 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110011; // iC= -973 
// vC = 14'b0000010111111110; // vC= 1534 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001110; // iC=-1074 
// vC = 14'b0000010111111000; // vC= 1528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001010; // iC=-1014 
// vC = 14'b0000011011011001; // vC= 1753 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010010; // iC=-1070 
// vC = 14'b0000011000111011; // vC= 1595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011001; // iC= -935 
// vC = 14'b0000011000111111; // vC= 1599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101111; // iC= -977 
// vC = 14'b0000011010110101; // vC= 1717 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111011; // iC=-1029 
// vC = 14'b0000011001100001; // vC= 1633 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100111; // iC=-1049 
// vC = 14'b0000011001000001; // vC= 1601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110001; // iC= -975 
// vC = 14'b0000011011011101; // vC= 1757 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001001; // iC= -951 
// vC = 14'b0000011001101110; // vC= 1646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011001; // iC=-1127 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000101; // iC=-1083 
// vC = 14'b0000011010000010; // vC= 1666 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011000; // iC=-1128 
// vC = 14'b0000011010101011; // vC= 1707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001011; // iC=-1205 
// vC = 14'b0000011011001110; // vC= 1742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000101; // iC=-1211 
// vC = 14'b0000010111001111; // vC= 1487 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101000; // iC=-1240 
// vC = 14'b0000011010110100; // vC= 1716 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101111; // iC=-1169 
// vC = 14'b0000011010011100; // vC= 1692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101011; // iC=-1109 
// vC = 14'b0000011000101111; // vC= 1583 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000110; // iC=-1146 
// vC = 14'b0000010111010011; // vC= 1491 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010000; // iC=-1392 
// vC = 14'b0000010111100010; // vC= 1506 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111101; // iC=-1347 
// vC = 14'b0000010111010010; // vC= 1490 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011010; // iC=-1382 
// vC = 14'b0000010101110010; // vC= 1394 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101001; // iC=-1303 
// vC = 14'b0000011001011101; // vC= 1629 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010101; // iC=-1387 
// vC = 14'b0000011001011000; // vC= 1624 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000001; // iC=-1343 
// vC = 14'b0000011001011101; // vC= 1629 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000110; // iC=-1274 
// vC = 14'b0000010110011110; // vC= 1438 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100000; // iC=-1440 
// vC = 14'b0000011001001001; // vC= 1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010001; // iC=-1327 
// vC = 14'b0000011010000000; // vC= 1664 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011111; // iC=-1441 
// vC = 14'b0000010110101101; // vC= 1453 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110010; // iC=-1422 
// vC = 14'b0000011001011110; // vC= 1630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101001; // iC=-1623 
// vC = 14'b0000010110101101; // vC= 1453 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000001; // iC=-1343 
// vC = 14'b0000010100100111; // vC= 1319 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110001; // iC=-1551 
// vC = 14'b0000011001001001; // vC= 1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001111; // iC=-1649 
// vC = 14'b0000010101000110; // vC= 1350 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010111; // iC=-1641 
// vC = 14'b0000010110010011; // vC= 1427 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100001; // iC=-1567 
// vC = 14'b0000010100100101; // vC= 1317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110100; // iC=-1612 
// vC = 14'b0000010101011101; // vC= 1373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011110; // iC=-1442 
// vC = 14'b0000010111111110; // vC= 1534 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111111; // iC=-1537 
// vC = 14'b0000010101111001; // vC= 1401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100011; // iC=-1437 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101011; // iC=-1557 
// vC = 14'b0000010101011110; // vC= 1374 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101100; // iC=-1620 
// vC = 14'b0000010011111110; // vC= 1278 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110101; // iC=-1547 
// vC = 14'b0000010111000001; // vC= 1473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101100; // iC=-1492 
// vC = 14'b0000010101111111; // vC= 1407 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001001; // iC=-1655 
// vC = 14'b0000010101010010; // vC= 1362 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100100; // iC=-1564 
// vC = 14'b0000010101000110; // vC= 1350 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011111; // iC=-1825 
// vC = 14'b0000010010111001; // vC= 1209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010000; // iC=-1712 
// vC = 14'b0000010101110001; // vC= 1393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010110; // iC=-1834 
// vC = 14'b0000010110110010; // vC= 1458 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100100; // iC=-1564 
// vC = 14'b0000010101010001; // vC= 1361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b0000010110100100; // vC= 1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101000; // iC=-1688 
// vC = 14'b0000010111010101; // vC= 1493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001000; // iC=-1656 
// vC = 14'b0000010010101010; // vC= 1194 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101010; // iC=-1622 
// vC = 14'b0000010100010110; // vC= 1302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b0000010101110011; // vC= 1395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111110; // iC=-1794 
// vC = 14'b0000010101100110; // vC= 1382 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b0000010100110011; // vC= 1331 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b0000010101110011; // vC= 1395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110111; // iC=-1673 
// vC = 14'b0000010010101101; // vC= 1197 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010100; // iC=-1708 
// vC = 14'b0000010011000100; // vC= 1220 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111101; // iC=-1731 
// vC = 14'b0000010101000010; // vC= 1346 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011001; // iC=-1895 
// vC = 14'b0000010001100011; // vC= 1123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100011; // iC=-1821 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b0000010010011000; // vC= 1176 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110111; // iC=-1673 
// vC = 14'b0000010010001110; // vC= 1166 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110011; // iC=-1869 
// vC = 14'b0000010100100011; // vC= 1315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111010; // iC=-1862 
// vC = 14'b0000010010110101; // vC= 1205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111110; // iC=-1922 
// vC = 14'b0000010001101110; // vC= 1134 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000010010111100; // vC= 1212 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001010; // iC=-1910 
// vC = 14'b0000010010010001; // vC= 1169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b0000010100000000; // vC= 1280 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000111; // iC=-1721 
// vC = 14'b0000010001101111; // vC= 1135 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b0000010010101001; // vC= 1193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b0000010000000111; // vC= 1031 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010111; // iC=-1833 
// vC = 14'b0000010010011100; // vC= 1180 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000010010101101; // vC= 1197 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b0000010000011011; // vC= 1051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000010001000011; // vC= 1091 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b0000001111011001; // vC=  985 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b0000010001110100; // vC= 1140 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b0000001111100110; // vC=  998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b0000001111010100; // vC=  980 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001011; // iC=-1973 
// vC = 14'b0000001111110010; // vC= 1010 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011110; // iC=-1762 
// vC = 14'b0000010010010111; // vC= 1175 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010101; // iC=-1771 
// vC = 14'b0000010001110010; // vC= 1138 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111111; // iC=-1921 
// vC = 14'b0000001110011010; // vC=  922 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b0000010001011011; // vC= 1115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111010; // iC=-1798 
// vC = 14'b0000010010100000; // vC= 1184 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001000; // iC=-2040 
// vC = 14'b0000001101111001; // vC=  889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b0000010000100100; // vC= 1060 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b0000010001100001; // vC= 1121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001111; // iC=-1777 
// vC = 14'b0000010000010111; // vC= 1047 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011010; // iC=-2022 
// vC = 14'b0000001101110101; // vC=  885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010010; // iC=-1966 
// vC = 14'b0000010000001101; // vC= 1037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101110; // iC=-1810 
// vC = 14'b0000001111111010; // vC= 1018 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b0000010000101101; // vC= 1069 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111101; // iC=-1859 
// vC = 14'b0000001100110101; // vC=  821 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101010; // iC=-2070 
// vC = 14'b0000001101010010; // vC=  850 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b0000001101100010; // vC=  866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001001; // iC=-2039 
// vC = 14'b0000001111110001; // vC= 1009 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011101; // iC=-1827 
// vC = 14'b0000010001000100; // vC= 1092 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110101; // iC=-1803 
// vC = 14'b0000001110011000; // vC=  920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010001; // iC=-2031 
// vC = 14'b0000001111011101; // vC=  989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000010000000111; // vC= 1031 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001111; // iC=-2097 
// vC = 14'b0000001110101011; // vC=  939 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b0000001101010101; // vC=  853 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110111; // iC=-1865 
// vC = 14'b0000001101010100; // vC=  852 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b0000001110100101; // vC=  933 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011101; // iC=-2083 
// vC = 14'b0000001100101110; // vC=  814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000001011001010; // vC=  714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b0000001110010101; // vC=  917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b0000001111011100; // vC=  988 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000001101000001; // vC=  833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100111; // iC=-2009 
// vC = 14'b0000001011110111; // vC=  759 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000001011010110; // vC=  726 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b0000001110111000; // vC=  952 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b0000001010101110; // vC=  686 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b0000001010000011; // vC=  643 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001010; // iC=-1910 
// vC = 14'b0000001010101111; // vC=  687 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b0000001100111110; // vC=  830 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b0000001101010100; // vC=  852 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b0000001010011101; // vC=  669 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000100; // iC=-2108 
// vC = 14'b0000001101100001; // vC=  865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101000; // iC=-1880 
// vC = 14'b0000001100010001; // vC=  785 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111101; // iC=-1795 
// vC = 14'b0000001010011111; // vC=  671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111100; // iC=-1988 
// vC = 14'b0000001100111100; // vC=  828 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000100; // iC=-1916 
// vC = 14'b0000001001011110; // vC=  606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b0000001011010100; // vC=  724 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b0000001100100110; // vC=  806 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b0000001001110111; // vC=  631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b0000001011111101; // vC=  765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000001001010111; // vC=  599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b0000001000011110; // vC=  542 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b0000001011111000; // vC=  760 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000001001101000; // vC=  616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b0000001011010011; // vC=  723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b0000001011100100; // vC=  740 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110011; // iC=-1805 
// vC = 14'b0000001011010111; // vC=  727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b0000001001101010; // vC=  618 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100111; // iC=-1817 
// vC = 14'b0000001000001110; // vC=  526 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010110; // iC=-2090 
// vC = 14'b0000001001000110; // vC=  582 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000111; // iC=-2105 
// vC = 14'b0000001000110000; // vC=  560 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101001; // iC=-2071 
// vC = 14'b0000000110001100; // vC=  396 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001001; // iC=-1847 
// vC = 14'b0000000110011100; // vC=  412 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b0000001001111011; // vC=  635 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101111; // iC=-1809 
// vC = 14'b0000001000001110; // vC=  526 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000000110101010; // vC=  426 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010110; // iC=-2090 
// vC = 14'b0000000111011111; // vC=  479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010111; // iC=-1897 
// vC = 14'b0000001001010001; // vC=  593 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b0000001000110011; // vC=  563 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010001; // iC=-2095 
// vC = 14'b0000000110010101; // vC=  405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110000; // iC=-2000 
// vC = 14'b0000001001101101; // vC=  621 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001111; // iC=-1905 
// vC = 14'b0000000111010100; // vC=  468 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101101; // iC=-2067 
// vC = 14'b0000001001000100; // vC=  580 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b0000000111001110; // vC=  462 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b0000000110111011; // vC=  443 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b0000001000111011; // vC=  571 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b0000000111101001; // vC=  489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b0000001000101100; // vC=  556 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b0000000101000110; // vC=  326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000000101000111; // vC=  327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b0000000100000110; // vC=  262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001101; // iC=-1907 
// vC = 14'b0000000100000010; // vC=  258 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101111; // iC=-1873 
// vC = 14'b0000000100110000; // vC=  304 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000101; // iC=-2043 
// vC = 14'b0000000110110100; // vC=  436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101001; // iC=-2071 
// vC = 14'b0000000011011110; // vC=  222 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b0000000111000010; // vC=  450 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000001; // iC=-1791 
// vC = 14'b0000000011010011; // vC=  211 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000100; // iC=-1916 
// vC = 14'b0000000100100110; // vC=  294 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011011; // iC=-2085 
// vC = 14'b0000000100011010; // vC=  282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b0000000101001111; // vC=  335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000000101111010; // vC=  378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111110; // iC=-1794 
// vC = 14'b0000000111001101; // vC=  461 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b0000000110010011; // vC=  403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000000011001000; // vC=  200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111111; // iC=-2049 
// vC = 14'b0000000010011110; // vC=  158 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101111; // iC=-1937 
// vC = 14'b0000000101000000; // vC=  320 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b0000000110010010; // vC=  402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101110; // iC=-1874 
// vC = 14'b0000000011100011; // vC=  227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111010; // iC=-1862 
// vC = 14'b0000000011010110; // vC=  214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000000100100110; // vC=  294 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000001; // iC=-1791 
// vC = 14'b0000000101101110; // vC=  366 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000000; // iC=-1856 
// vC = 14'b0000000001101100; // vC=  108 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101110; // iC=-1874 
// vC = 14'b0000000100100000; // vC=  288 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100111; // iC=-2009 
// vC = 14'b0000000100100110; // vC=  294 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011110; // iC=-2018 
// vC = 14'b0000000100011100; // vC=  284 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b0000000010000110; // vC=  134 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110010; // iC=-1934 
// vC = 14'b0000000000011101; // vC=   29 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b0000000011100110; // vC=  230 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000000000101110; // vC=   46 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000110; // iC=-1914 
// vC = 14'b0000000001000101; // vC=   69 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000000001001111; // vC=   79 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b0000000000100101; // vC=   37 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b0000000000101001; // vC=   41 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011000; // iC=-1768 
// vC = 14'b1111111111001001; // vC=  -55 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000000011101011; // vC=  235 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b0000000000100101; // vC=   37 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100010; // iC=-2014 
// vC = 14'b0000000011101000; // vC=  232 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b1111111111000101; // vC=  -59 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b0000000001001100; // vC=   76 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000000001110000; // vC=  112 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111001; // iC=-1991 
// vC = 14'b0000000000001101; // vC=   13 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101011; // iC=-1749 
// vC = 14'b1111111110001110; // vC= -114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b0000000000010100; // vC=   20 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000000000010110; // vC=   22 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b0000000000001110; // vC=   14 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100111; // iC=-1753 
// vC = 14'b0000000010001000; // vC=  136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010111; // iC=-2025 
// vC = 14'b1111111111100100; // vC=  -28 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011010; // iC=-1894 
// vC = 14'b1111111110011101; // vC=  -99 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b0000000000000100; // vC=    4 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b1111111110001100; // vC= -116 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000001; // iC=-1727 
// vC = 14'b0000000001110010; // vC=  114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b0000000000101011; // vC=   43 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000001; // iC=-1983 
// vC = 14'b1111111111010111; // vC=  -41 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b1111111101000100; // vC= -188 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110101; // iC=-1867 
// vC = 14'b1111111111111100; // vC=   -4 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100001; // iC=-1887 
// vC = 14'b1111111101011001; // vC= -167 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110011; // iC=-1741 
// vC = 14'b1111111110101001; // vC=  -87 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101000; // iC=-1816 
// vC = 14'b1111111111101101; // vC=  -19 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111110; // iC=-1922 
// vC = 14'b1111111100000001; // vC= -255 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100010; // iC=-1886 
// vC = 14'b1111111100011101; // vC= -227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111101; // iC=-1795 
// vC = 14'b1111111101101110; // vC= -146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011110; // iC=-1762 
// vC = 14'b0000000000000111; // vC=    7 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001101; // iC=-1779 
// vC = 14'b1111111011100011; // vC= -285 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000110; // iC=-1850 
// vC = 14'b1111111111001010; // vC=  -54 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b1111111110010110; // vC= -106 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b1111111101000001; // vC= -191 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100100; // iC=-1884 
// vC = 14'b1111111110110011; // vC=  -77 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b1111111110001110; // vC= -114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011111; // iC=-1953 
// vC = 14'b1111111100110001; // vC= -207 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b1111111101001010; // vC= -182 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b1111111111000111; // vC=  -57 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b1111111100000111; // vC= -249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b1111111011011000; // vC= -296 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b1111111100001010; // vC= -246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000001; // iC=-1919 
// vC = 14'b1111111010010100; // vC= -364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001011; // iC=-1973 
// vC = 14'b1111111110110110; // vC=  -74 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010000; // iC=-1712 
// vC = 14'b1111111110100010; // vC=  -94 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111111; // iC=-1985 
// vC = 14'b1111111011101111; // vC= -273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010110; // iC=-1898 
// vC = 14'b1111111101011100; // vC= -164 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b1111111010110100; // vC= -332 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011110; // iC=-1698 
// vC = 14'b1111111001010011; // vC= -429 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100010; // iC=-1694 
// vC = 14'b1111111011011010; // vC= -294 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111110; // iC=-1666 
// vC = 14'b1111111101111101; // vC= -131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000100; // iC=-1980 
// vC = 14'b1111111000110111; // vC= -457 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011110; // iC=-1762 
// vC = 14'b1111111100010010; // vC= -238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b1111111000111100; // vC= -452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001010; // iC=-1654 
// vC = 14'b1111111011001001; // vC= -311 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b1111111011010110; // vC= -298 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011010; // iC=-1766 
// vC = 14'b1111111000110101; // vC= -459 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110011; // iC=-1933 
// vC = 14'b1111111011001100; // vC= -308 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111010; // iC=-1862 
// vC = 14'b1111111000001101; // vC= -499 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b1111111100101100; // vC= -212 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111001; // iC=-1799 
// vC = 14'b1111111000101101; // vC= -467 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b1111111011111010; // vC= -262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b1111111100010010; // vC= -238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b1111111011101001; // vC= -279 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010101; // iC=-1771 
// vC = 14'b1111111010010100; // vC= -364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111011; // iC=-1733 
// vC = 14'b1111111010010001; // vC= -367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101111; // iC=-1937 
// vC = 14'b1111110111101000; // vC= -536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b1111111011100011; // vC= -285 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010101; // iC=-1835 
// vC = 14'b1111110111110000; // vC= -528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b1111111010011101; // vC= -355 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110111; // iC=-1801 
// vC = 14'b1111111000111101; // vC= -451 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010100; // iC=-1644 
// vC = 14'b1111110111101010; // vC= -534 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011010; // iC=-1894 
// vC = 14'b1111111001100010; // vC= -414 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100101; // iC=-1627 
// vC = 14'b1111110110111111; // vC= -577 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011101; // iC=-1699 
// vC = 14'b1111110110010110; // vC= -618 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000000; // iC=-1792 
// vC = 14'b1111110111001111; // vC= -561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000110; // iC=-1658 
// vC = 14'b1111110110111000; // vC= -584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b1111111010100001; // vC= -351 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110110; // iC=-1674 
// vC = 14'b1111111001000100; // vC= -444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110011; // iC=-1677 
// vC = 14'b1111111000000010; // vC= -510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000011; // iC=-1597 
// vC = 14'b1111111010010111; // vC= -361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100110; // iC=-1690 
// vC = 14'b1111110101010100; // vC= -684 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100000; // iC=-1632 
// vC = 14'b1111111000010101; // vC= -491 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110101; // iC=-1739 
// vC = 14'b1111111000110001; // vC= -463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010110; // iC=-1706 
// vC = 14'b1111111000100010; // vC= -478 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110000; // iC=-1680 
// vC = 14'b1111110101100111; // vC= -665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011011; // iC=-1765 
// vC = 14'b1111110111111111; // vC= -513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b1111111001010111; // vC= -425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011101; // iC=-1635 
// vC = 14'b1111111001100000; // vC= -416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110011; // iC=-1805 
// vC = 14'b1111111001011010; // vC= -422 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b1111110101111100; // vC= -644 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010111; // iC=-1577 
// vC = 14'b1111110111111111; // vC= -513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101100; // iC=-1556 
// vC = 14'b1111110101101100; // vC= -660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111010; // iC=-1670 
// vC = 14'b1111110111101000; // vC= -536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001100; // iC=-1780 
// vC = 14'b1111110100000110; // vC= -762 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000000; // iC=-1856 
// vC = 14'b1111110110001000; // vC= -632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110010; // iC=-1806 
// vC = 14'b1111110011101101; // vC= -787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100111; // iC=-1561 
// vC = 14'b1111110101111110; // vC= -642 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011001; // iC=-1767 
// vC = 14'b1111110111011111; // vC= -545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111000; // iC=-1608 
// vC = 14'b1111110100100111; // vC= -729 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111001; // iC=-1799 
// vC = 14'b1111110111100010; // vC= -542 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111100; // iC=-1796 
// vC = 14'b1111110110101101; // vC= -595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101111; // iC=-1617 
// vC = 14'b1111110011001001; // vC= -823 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011101; // iC=-1827 
// vC = 14'b1111110110001100; // vC= -628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011111; // iC=-1825 
// vC = 14'b1111110110011001; // vC= -615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001000; // iC=-1528 
// vC = 14'b1111110011011001; // vC= -807 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110011; // iC=-1805 
// vC = 14'b1111110101001001; // vC= -695 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101100; // iC=-1748 
// vC = 14'b1111110101011010; // vC= -678 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000101; // iC=-1595 
// vC = 14'b1111110100100100; // vC= -732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010110; // iC=-1578 
// vC = 14'b1111110011010001; // vC= -815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001111; // iC=-1585 
// vC = 14'b1111110010001101; // vC= -883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101110; // iC=-1618 
// vC = 14'b1111110110000011; // vC= -637 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100111; // iC=-1625 
// vC = 14'b1111110101001110; // vC= -690 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011001; // iC=-1767 
// vC = 14'b1111110110001101; // vC= -627 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001111; // iC=-1777 
// vC = 14'b1111110010001000; // vC= -888 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000101; // iC=-1595 
// vC = 14'b1111110011001001; // vC= -823 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010111; // iC=-1641 
// vC = 14'b1111110001101111; // vC= -913 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011110; // iC=-1698 
// vC = 14'b1111110001011100; // vC= -932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000111; // iC=-1465 
// vC = 14'b1111110001101001; // vC= -919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110101; // iC=-1483 
// vC = 14'b1111110001001011; // vC= -949 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011011; // iC=-1573 
// vC = 14'b1111110101011111; // vC= -673 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010001; // iC=-1519 
// vC = 14'b1111110011011001; // vC= -807 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100101; // iC=-1755 
// vC = 14'b1111110011000001; // vC= -831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001110; // iC=-1458 
// vC = 14'b1111110010001010; // vC= -886 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001110; // iC=-1714 
// vC = 14'b1111110101100001; // vC= -671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000101; // iC=-1723 
// vC = 14'b1111110100110100; // vC= -716 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000111; // iC=-1465 
// vC = 14'b1111110010110001; // vC= -847 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001010; // iC=-1590 
// vC = 14'b1111110100101010; // vC= -726 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111001; // iC=-1607 
// vC = 14'b1111110100010011; // vC= -749 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010000; // iC=-1520 
// vC = 14'b1111110001001001; // vC= -951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000111; // iC=-1465 
// vC = 14'b1111110000110110; // vC= -970 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111001; // iC=-1671 
// vC = 14'b1111110100000000; // vC= -768 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100001; // iC=-1503 
// vC = 14'b1111110010000001; // vC= -895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011111; // iC=-1569 
// vC = 14'b1111110011111100; // vC= -772 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010010; // iC=-1454 
// vC = 14'b1111110011101110; // vC= -786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011100; // iC=-1508 
// vC = 14'b1111110010110010; // vC= -846 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011000; // iC=-1384 
// vC = 14'b1111110000110010; // vC= -974 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111000; // iC=-1544 
// vC = 14'b1111110100000101; // vC= -763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100101; // iC=-1691 
// vC = 14'b1111110000010111; // vC=-1001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011010; // iC=-1574 
// vC = 14'b1111110001001010; // vC= -950 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000101; // iC=-1531 
// vC = 14'b1111110000011000; // vC=-1000 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011100; // iC=-1636 
// vC = 14'b1111110010101111; // vC= -849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011011; // iC=-1509 
// vC = 14'b1111101111011010; // vC=-1062 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010010; // iC=-1390 
// vC = 14'b1111110000011010; // vC= -998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101011; // iC=-1557 
// vC = 14'b1111110011011100; // vC= -804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001000; // iC=-1464 
// vC = 14'b1111110000110000; // vC= -976 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100110; // iC=-1498 
// vC = 14'b1111110000111011; // vC= -965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100011; // iC=-1629 
// vC = 14'b1111101111101010; // vC=-1046 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111010; // iC=-1414 
// vC = 14'b1111110001101101; // vC= -915 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011010; // iC=-1446 
// vC = 14'b1111110010111110; // vC= -834 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000000; // iC=-1536 
// vC = 14'b1111110000010010; // vC=-1006 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100000; // iC=-1632 
// vC = 14'b1111101111011000; // vC=-1064 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111111; // iC=-1601 
// vC = 14'b1111110000100100; // vC= -988 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111011; // iC=-1541 
// vC = 14'b1111110000011010; // vC= -998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111110; // iC=-1346 
// vC = 14'b1111110001100110; // vC= -922 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000001; // iC=-1471 
// vC = 14'b1111110000111110; // vC= -962 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100110; // iC=-1562 
// vC = 14'b1111110000011011; // vC= -997 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111110; // iC=-1602 
// vC = 14'b1111110001100001; // vC= -927 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100110; // iC=-1434 
// vC = 14'b1111101110000011; // vC=-1149 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010101; // iC=-1515 
// vC = 14'b1111110001000011; // vC= -957 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100111; // iC=-1369 
// vC = 14'b1111101111110011; // vC=-1037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001010; // iC=-1590 
// vC = 14'b1111110001001010; // vC= -950 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110001; // iC=-1423 
// vC = 14'b1111101110001100; // vC=-1140 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100100; // iC=-1564 
// vC = 14'b1111101111011100; // vC=-1060 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101110; // iC=-1490 
// vC = 14'b1111101111010011; // vC=-1069 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001011; // iC=-1461 
// vC = 14'b1111101111100000; // vC=-1056 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100011; // iC=-1373 
// vC = 14'b1111110000111001; // vC= -967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000000; // iC=-1408 
// vC = 14'b1111101111010000; // vC=-1072 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010101; // iC=-1515 
// vC = 14'b1111101100010011; // vC=-1261 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100001; // iC=-1247 
// vC = 14'b1111101101001010; // vC=-1206 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000100; // iC=-1340 
// vC = 14'b1111110000001111; // vC=-1009 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110110; // iC=-1482 
// vC = 14'b1111101110111000; // vC=-1096 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111101; // iC=-1347 
// vC = 14'b1111101100100100; // vC=-1244 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100001; // iC=-1375 
// vC = 14'b1111101101101110; // vC=-1170 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101110; // iC=-1426 
// vC = 14'b1111101101101100; // vC=-1172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110100; // iC=-1228 
// vC = 14'b1111101111101110; // vC=-1042 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001100; // iC=-1524 
// vC = 14'b1111101100000110; // vC=-1274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110101; // iC=-1355 
// vC = 14'b1111101111001101; // vC=-1075 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111001; // iC=-1351 
// vC = 14'b1111101100111000; // vC=-1224 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010000; // iC=-1392 
// vC = 14'b1111101111001111; // vC=-1073 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011111; // iC=-1505 
// vC = 14'b1111101110100101; // vC=-1115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100110; // iC=-1370 
// vC = 14'b1111101101001000; // vC=-1208 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100100; // iC=-1244 
// vC = 14'b1111101111000110; // vC=-1082 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011010; // iC=-1190 
// vC = 14'b1111101110000101; // vC=-1147 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010011; // iC=-1389 
// vC = 14'b1111101101101100; // vC=-1172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110100; // iC=-1228 
// vC = 14'b1111101101011010; // vC=-1190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011111; // iC=-1249 
// vC = 14'b1111101110001111; // vC=-1137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100101; // iC=-1435 
// vC = 14'b1111101110000000; // vC=-1152 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101110; // iC=-1170 
// vC = 14'b1111101011001100; // vC=-1332 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101011; // iC=-1365 
// vC = 14'b1111101111010010; // vC=-1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010011; // iC=-1453 
// vC = 14'b1111101110001110; // vC=-1138 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010100; // iC=-1324 
// vC = 14'b1111101100001011; // vC=-1269 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010110; // iC=-1258 
// vC = 14'b1111101101100111; // vC=-1177 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111001; // iC=-1223 
// vC = 14'b1111101100110010; // vC=-1230 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001110; // iC=-1330 
// vC = 14'b1111101100100111; // vC=-1241 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101010; // iC=-1430 
// vC = 14'b1111101100011011; // vC=-1253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110011; // iC=-1421 
// vC = 14'b1111101010011001; // vC=-1383 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010000; // iC=-1200 
// vC = 14'b1111101001111001; // vC=-1415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010101; // iC=-1387 
// vC = 14'b1111101011100110; // vC=-1306 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100000; // iC=-1312 
// vC = 14'b1111101011110010; // vC=-1294 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100100; // iC=-1244 
// vC = 14'b1111101110000100; // vC=-1148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111101; // iC=-1091 
// vC = 14'b1111101101111011; // vC=-1157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101100; // iC=-1364 
// vC = 14'b1111101010011110; // vC=-1378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010101; // iC=-1131 
// vC = 14'b1111101011011110; // vC=-1314 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000011; // iC=-1149 
// vC = 14'b1111101010111101; // vC=-1347 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011111; // iC=-1121 
// vC = 14'b1111101101000101; // vC=-1211 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000000; // iC=-1216 
// vC = 14'b1111101100000110; // vC=-1274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001111; // iC=-1265 
// vC = 14'b1111101010011011; // vC=-1381 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011111; // iC=-1377 
// vC = 14'b1111101011100010; // vC=-1310 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001101; // iC=-1331 
// vC = 14'b1111101100111000; // vC=-1224 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001110; // iC=-1138 
// vC = 14'b1111101100101111; // vC=-1233 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011001; // iC=-1063 
// vC = 14'b1111101010001101; // vC=-1395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111000; // iC=-1032 
// vC = 14'b1111101101000100; // vC=-1212 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000111; // iC=-1081 
// vC = 14'b1111101011100110; // vC=-1306 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100010; // iC=-1118 
// vC = 14'b1111101011111111; // vC=-1281 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011000; // iC=-1192 
// vC = 14'b1111101000111110; // vC=-1474 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101000; // iC=-1112 
// vC = 14'b1111101010010110; // vC=-1386 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011111; // iC=-1121 
// vC = 14'b1111101100100010; // vC=-1246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100010; // iC=-1182 
// vC = 14'b1111101011000101; // vC=-1339 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000101; // iC=-1275 
// vC = 14'b1111101001111000; // vC=-1416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011111; // iC=-1313 
// vC = 14'b1111101100001100; // vC=-1268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000100; // iC=-1276 
// vC = 14'b1111101000001011; // vC=-1525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001110; // iC=-1010 
// vC = 14'b1111101011011000; // vC=-1320 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100100; // iC= -988 
// vC = 14'b1111101011010010; // vC=-1326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001101; // iC=-1139 
// vC = 14'b1111101010001001; // vC=-1399 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001001; // iC=-1207 
// vC = 14'b1111101000001100; // vC=-1524 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100000; // iC=-1248 
// vC = 14'b1111101010110010; // vC=-1358 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010001; // iC=-1135 
// vC = 14'b1111101100000101; // vC=-1275 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101110; // iC=-1106 
// vC = 14'b1111101011010111; // vC=-1321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101000; // iC=-1240 
// vC = 14'b1111101000010001; // vC=-1519 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001010; // iC=-1078 
// vC = 14'b1111101001011010; // vC=-1446 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000110; // iC=-1210 
// vC = 14'b1111100111110010; // vC=-1550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011110; // iC=-1186 
// vC = 14'b1111101011011110; // vC=-1314 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110010; // iC= -974 
// vC = 14'b1111101001010101; // vC=-1451 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110001; // iC=-1167 
// vC = 14'b1111101010000010; // vC=-1406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010000; // iC=-1136 
// vC = 14'b1111101001110000; // vC=-1424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111010; // iC=-1222 
// vC = 14'b1111100111011111; // vC=-1569 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100111; // iC= -921 
// vC = 14'b1111100110101110; // vC=-1618 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011101; // iC=-1187 
// vC = 14'b1111100111101000; // vC=-1560 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000110; // iC=-1082 
// vC = 14'b1111101010101100; // vC=-1364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000100; // iC=-1020 
// vC = 14'b1111101001111101; // vC=-1411 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010000; // iC=-1136 
// vC = 14'b1111101011011000; // vC=-1320 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011101; // iC=-1187 
// vC = 14'b1111100111100000; // vC=-1568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b1111100110100100; // vC=-1628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000101; // iC= -955 
// vC = 14'b1111101001100011; // vC=-1437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001101; // iC= -947 
// vC = 14'b1111100110011000; // vC=-1640 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000110; // iC=-1082 
// vC = 14'b1111101001101010; // vC=-1430 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111000; // iC=-1160 
// vC = 14'b1111101001100000; // vC=-1440 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110110; // iC= -842 
// vC = 14'b1111101000010100; // vC=-1516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101010; // iC= -982 
// vC = 14'b1111100110110010; // vC=-1614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100010; // iC= -990 
// vC = 14'b1111101001110100; // vC=-1420 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111101; // iC= -963 
// vC = 14'b1111101001100110; // vC=-1434 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000110; // iC= -826 
// vC = 14'b1111101010000010; // vC=-1406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011000; // iC=-1064 
// vC = 14'b1111101000000001; // vC=-1535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010011; // iC=-1005 
// vC = 14'b1111100111100000; // vC=-1568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111010; // iC=-1030 
// vC = 14'b1111101000111011; // vC=-1477 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011111; // iC= -929 
// vC = 14'b1111100111101010; // vC=-1558 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110101; // iC= -843 
// vC = 14'b1111100101100100; // vC=-1692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000101; // iC=-1019 
// vC = 14'b1111100110111110; // vC=-1602 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001110; // iC=-1074 
// vC = 14'b1111101001101001; // vC=-1431 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100010; // iC= -862 
// vC = 14'b1111101001010011; // vC=-1453 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011111; // iC=-1057 
// vC = 14'b1111100111001101; // vC=-1587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111110; // iC= -962 
// vC = 14'b1111101000110110; // vC=-1482 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000111; // iC= -889 
// vC = 14'b1111100111000001; // vC=-1599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111011; // iC= -773 
// vC = 14'b1111100111010010; // vC=-1582 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111110; // iC= -770 
// vC = 14'b1111101000010111; // vC=-1513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110000; // iC= -784 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000101; // iC= -827 
// vC = 14'b1111100111000001; // vC=-1599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110110; // iC= -842 
// vC = 14'b1111100110010111; // vC=-1641 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110001; // iC= -847 
// vC = 14'b1111100111011011; // vC=-1573 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010001; // iC= -815 
// vC = 14'b1111100110110010; // vC=-1614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111100; // iC= -964 
// vC = 14'b1111100101011001; // vC=-1703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101111; // iC= -785 
// vC = 14'b1111100110101110; // vC=-1618 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100000; // iC= -736 
// vC = 14'b1111100111001101; // vC=-1587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011001; // iC= -871 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101000; // iC= -984 
// vC = 14'b1111100110110111; // vC=-1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110001; // iC= -719 
// vC = 14'b1111101000110010; // vC=-1486 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010110; // iC= -810 
// vC = 14'b1111101001001011; // vC=-1461 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011010; // iC= -934 
// vC = 14'b1111100110010111; // vC=-1641 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000001; // iC= -895 
// vC = 14'b1111101000111110; // vC=-1474 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101010; // iC= -854 
// vC = 14'b1111101000100101; // vC=-1499 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010111; // iC= -873 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110000; // iC= -720 
// vC = 14'b1111100111011100; // vC=-1572 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101110; // iC= -850 
// vC = 14'b1111100111011110; // vC=-1570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010010; // iC= -814 
// vC = 14'b1111100100110010; // vC=-1742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100110; // iC= -666 
// vC = 14'b1111100110011111; // vC=-1633 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101100; // iC= -852 
// vC = 14'b1111100100111011; // vC=-1733 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110111; // iC= -841 
// vC = 14'b1111100110011100; // vC=-1636 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010111; // iC= -745 
// vC = 14'b1111100101010001; // vC=-1711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110110; // iC= -842 
// vC = 14'b1111100110101101; // vC=-1619 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001101; // iC= -883 
// vC = 14'b1111100110100001; // vC=-1631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011110; // iC= -610 
// vC = 14'b1111100110001110; // vC=-1650 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110011; // iC= -653 
// vC = 14'b1111101000101100; // vC=-1492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101001; // iC= -855 
// vC = 14'b1111100110101111; // vC=-1617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101110; // iC= -850 
// vC = 14'b1111100111101000; // vC=-1560 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011010; // iC= -742 
// vC = 14'b1111100111101101; // vC=-1555 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100101; // iC= -795 
// vC = 14'b1111100011011111; // vC=-1825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000111; // iC= -633 
// vC = 14'b1111101000001011; // vC=-1525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101010; // iC= -854 
// vC = 14'b1111100111100110; // vC=-1562 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000110; // iC= -570 
// vC = 14'b1111100011010011; // vC=-1837 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100001; // iC= -799 
// vC = 14'b1111100011100000; // vC=-1824 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001011; // iC= -693 
// vC = 14'b1111100111111001; // vC=-1543 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100001; // iC= -735 
// vC = 14'b1111100100010000; // vC=-1776 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110010; // iC= -590 
// vC = 14'b1111100011011101; // vC=-1827 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110110; // iC= -650 
// vC = 14'b1111100111000010; // vC=-1598 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111101; // iC= -707 
// vC = 14'b1111100011000111; // vC=-1849 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111110110; // iC= -522 
// vC = 14'b1111100111000011; // vC=-1597 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101010; // iC= -790 
// vC = 14'b1111100110111010; // vC=-1606 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011000; // iC= -552 
// vC = 14'b1111100101111100; // vC=-1668 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010010; // iC= -558 
// vC = 14'b1111100110110110; // vC=-1610 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111110111; // iC= -521 
// vC = 14'b1111100111001001; // vC=-1591 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110110; // iC= -650 
// vC = 14'b1111100011110101; // vC=-1803 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110010; // iC= -718 
// vC = 14'b1111100110101000; // vC=-1624 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010101; // iC= -555 
// vC = 14'b1111100111001010; // vC=-1590 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100000; // iC= -544 
// vC = 14'b1111100110110110; // vC=-1610 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100100; // iC= -732 
// vC = 14'b1111100111010011; // vC=-1581 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000101; // iC= -763 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110010; // iC= -462 
// vC = 14'b1111100110010101; // vC=-1643 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110100; // iC= -460 
// vC = 14'b1111100110110011; // vC=-1613 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100010; // iC= -606 
// vC = 14'b1111100111011011; // vC=-1573 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011011; // iC= -485 
// vC = 14'b1111100101010000; // vC=-1712 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111001; // iC= -711 
// vC = 14'b1111100101111100; // vC=-1668 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111111; // iC= -577 
// vC = 14'b1111100011110000; // vC=-1808 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001101; // iC= -435 
// vC = 14'b1111100110000111; // vC=-1657 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100011; // iC= -605 
// vC = 14'b1111100100001101; // vC=-1779 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010010; // iC= -494 
// vC = 14'b1111100111010111; // vC=-1577 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100011; // iC= -477 
// vC = 14'b1111100100010001; // vC=-1775 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001100; // iC= -500 
// vC = 14'b1111100111010011; // vC=-1581 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010000; // iC= -368 
// vC = 14'b1111100110110011; // vC=-1613 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010101; // iC= -363 
// vC = 14'b1111100011100101; // vC=-1819 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100011; // iC= -349 
// vC = 14'b1111100110010001; // vC=-1647 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001000; // iC= -440 
// vC = 14'b1111100010001111; // vC=-1905 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101101; // iC= -275 
// vC = 14'b1111100111000101; // vC=-1595 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001110; // iC= -434 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111001; // iC= -391 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101010; // iC= -534 
// vC = 14'b1111100010111001; // vC=-1863 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010101001; // iC= -343 
// vC = 14'b1111100101001010; // vC=-1718 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010001; // iC= -303 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111000; // iC= -200 
// vC = 14'b1111100011010100; // vC=-1836 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111110; // iC= -450 
// vC = 14'b1111100100001010; // vC=-1782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111110; // iC= -322 
// vC = 14'b1111100100101001; // vC=-1751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000001; // iC= -191 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011110000; // iC= -272 
// vC = 14'b1111100101010010; // vC=-1710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101000; // iC= -216 
// vC = 14'b1111100110110011; // vC=-1613 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010000; // iC= -112 
// vC = 14'b1111100010011011; // vC=-1893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011101; // iC= -291 
// vC = 14'b1111100110001101; // vC=-1651 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010100; // iC= -300 
// vC = 14'b1111100010110011; // vC=-1869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010101010; // iC= -342 
// vC = 14'b1111100010000010; // vC=-1918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001000; // iC= -248 
// vC = 14'b1111100010110000; // vC=-1872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001110; // iC= -242 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111100; // iC=   -4 
// vC = 14'b1111100100010000; // vC=-1776 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101000; // iC= -152 
// vC = 14'b1111100011001001; // vC=-1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001010; // iC=  -54 
// vC = 14'b1111100011000100; // vC=-1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101110001; // iC= -143 
// vC = 14'b1111100110011111; // vC=-1633 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111011101; // iC=  -35 
// vC = 14'b1111100101011111; // vC=-1697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101001; // iC=   41 
// vC = 14'b1111100101101000; // vC=-1688 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100000; // iC=   96 
// vC = 14'b1111100100100100; // vC=-1756 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110011; // iC=  115 
// vC = 14'b1111100101100001; // vC=-1695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010001; // iC=  -47 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101000; // iC=  104 
// vC = 14'b1111100100010110; // vC=-1770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010010; // iC= -110 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000000; // iC=  128 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101110; // iC=  174 
// vC = 14'b1111100100001000; // vC=-1784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111000; // iC=  -72 
// vC = 14'b1111100111000010; // vC=-1598 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010100; // iC=   84 
// vC = 14'b1111100001111110; // vC=-1922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010000; // iC=  272 
// vC = 14'b1111100010111111; // vC=-1857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100011; // iC=   35 
// vC = 14'b1111100011001110; // vC=-1842 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100001; // iC=  225 
// vC = 14'b1111100101001101; // vC=-1715 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001010; // iC=  266 
// vC = 14'b1111100110110001; // vC=-1615 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111111; // iC=  255 
// vC = 14'b1111100110100011; // vC=-1629 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101011; // iC=  107 
// vC = 14'b1111100101110001; // vC=-1679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110000; // iC=  240 
// vC = 14'b1111100101001001; // vC=-1719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000001; // iC=  321 
// vC = 14'b1111100100001001; // vC=-1783 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010010; // iC=  466 
// vC = 14'b1111100101101010; // vC=-1686 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001110; // iC=  270 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110100; // iC=  372 
// vC = 14'b1111100011011010; // vC=-1830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110010; // iC=  370 
// vC = 14'b1111100011010101; // vC=-1835 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111100; // iC=  508 
// vC = 14'b1111100110101000; // vC=-1624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001011; // iC=  587 
// vC = 14'b1111100110001100; // vC=-1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010100; // iC=  532 
// vC = 14'b1111100011110100; // vC=-1804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010011; // iC=  339 
// vC = 14'b1111100010011100; // vC=-1892 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011110; // iC=  414 
// vC = 14'b1111100100000000; // vC=-1792 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010101; // iC=  597 
// vC = 14'b1111100110000011; // vC=-1661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001010; // iC=  650 
// vC = 14'b1111100100000011; // vC=-1789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110000; // iC=  560 
// vC = 14'b1111100110100011; // vC=-1629 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011001; // iC=  601 
// vC = 14'b1111100101111011; // vC=-1669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010101; // iC=  725 
// vC = 14'b1111100101010110; // vC=-1706 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101101; // iC=  493 
// vC = 14'b1111100101100101; // vC=-1691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101110; // iC=  622 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011011; // iC=  731 
// vC = 14'b1111100110000110; // vC=-1658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110000; // iC=  816 
// vC = 14'b1111100011100111; // vC=-1817 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000011; // iC=  707 
// vC = 14'b1111100011000110; // vC=-1850 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000101; // iC=  773 
// vC = 14'b1111100110110100; // vC=-1612 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000011; // iC=  707 
// vC = 14'b1111100111010101; // vC=-1579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001111; // iC=  719 
// vC = 14'b1111100101100000; // vC=-1696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001111; // iC=  655 
// vC = 14'b1111100110010111; // vC=-1641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101010; // iC=  874 
// vC = 14'b1111100100010011; // vC=-1773 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000111; // iC=  711 
// vC = 14'b1111100110010101; // vC=-1643 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011100; // iC=  924 
// vC = 14'b1111100101100101; // vC=-1691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100010; // iC=  994 
// vC = 14'b1111100110011010; // vC=-1638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111001; // iC=  761 
// vC = 14'b1111100110100001; // vC=-1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001000; // iC=  904 
// vC = 14'b1111100111111011; // vC=-1541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111000; // iC=  824 
// vC = 14'b1111100101000011; // vC=-1725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111111; // iC= 1087 
// vC = 14'b1111100111101011; // vC=-1557 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010001; // iC=  977 
// vC = 14'b1111100111001011; // vC=-1589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001101; // iC= 1037 
// vC = 14'b1111100110010000; // vC=-1648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100001; // iC=  993 
// vC = 14'b1111100110000110; // vC=-1658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101000; // iC= 1064 
// vC = 14'b1111100011111001; // vC=-1799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001101; // iC= 1101 
// vC = 14'b1111100100011100; // vC=-1764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111100; // iC=  956 
// vC = 14'b1111100110001010; // vC=-1654 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010101; // iC= 1237 
// vC = 14'b1111100101101011; // vC=-1685 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111000; // iC= 1272 
// vC = 14'b1111100100100011; // vC=-1757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011000; // iC= 1176 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110110; // iC= 1206 
// vC = 14'b1111100110001001; // vC=-1655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010011; // iC= 1299 
// vC = 14'b1111101000100010; // vC=-1502 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111010; // iC= 1338 
// vC = 14'b1111100110100111; // vC=-1625 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011101; // iC= 1309 
// vC = 14'b1111100111010010; // vC=-1582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001100; // iC= 1100 
// vC = 14'b1111100110010001; // vC=-1647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011001; // iC= 1113 
// vC = 14'b1111100110001011; // vC=-1653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110001; // iC= 1201 
// vC = 14'b1111100110001001; // vC=-1655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100001; // iC= 1377 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011101; // iC= 1181 
// vC = 14'b1111100110100111; // vC=-1625 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011111; // iC= 1247 
// vC = 14'b1111100111000111; // vC=-1593 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011010; // iC= 1498 
// vC = 14'b1111101000001101; // vC=-1523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100000; // iC= 1440 
// vC = 14'b1111100111101100; // vC=-1556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000011; // iC= 1475 
// vC = 14'b1111100101110110; // vC=-1674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101110; // iC= 1326 
// vC = 14'b1111101000011110; // vC=-1506 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101111; // iC= 1327 
// vC = 14'b1111101010100110; // vC=-1370 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000010; // iC= 1410 
// vC = 14'b1111100111101010; // vC=-1558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011100; // iC= 1372 
// vC = 14'b1111101001011101; // vC=-1443 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011001; // iC= 1497 
// vC = 14'b1111100111111010; // vC=-1542 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111001; // iC= 1401 
// vC = 14'b1111101001111100; // vC=-1412 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001100; // iC= 1356 
// vC = 14'b1111101010110001; // vC=-1359 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100100; // iC= 1444 
// vC = 14'b1111101000110011; // vC=-1485 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100101; // iC= 1445 
// vC = 14'b1111101001110001; // vC=-1423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011110; // iC= 1438 
// vC = 14'b1111100111011101; // vC=-1571 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111111; // iC= 1407 
// vC = 14'b1111101010000011; // vC=-1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101011; // iC= 1451 
// vC = 14'b1111101011001001; // vC=-1335 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010101; // iC= 1493 
// vC = 14'b1111101001111110; // vC=-1410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001111; // iC= 1615 
// vC = 14'b1111101000011110; // vC=-1506 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111011; // iC= 1467 
// vC = 14'b1111101010000110; // vC=-1402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011101; // iC= 1565 
// vC = 14'b1111101011011010; // vC=-1318 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100001; // iC= 1505 
// vC = 14'b1111101011011010; // vC=-1318 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100111; // iC= 1767 
// vC = 14'b1111101001000001; // vC=-1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001001; // iC= 1737 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001101; // iC= 1549 
// vC = 14'b1111101011111000; // vC=-1288 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011011; // iC= 1819 
// vC = 14'b1111101010101000; // vC=-1368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100101; // iC= 1637 
// vC = 14'b1111101001000001; // vC=-1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111011; // iC= 1531 
// vC = 14'b1111101001111101; // vC=-1411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110100; // iC= 1588 
// vC = 14'b1111101011110011; // vC=-1293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b1111101001110110; // vC=-1418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100001; // iC= 1697 
// vC = 14'b1111101000100001; // vC=-1503 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111111; // iC= 1727 
// vC = 14'b1111101001001000; // vC=-1464 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000110; // iC= 1606 
// vC = 14'b1111101011000110; // vC=-1338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100001; // iC= 1761 
// vC = 14'b1111101010101000; // vC=-1368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011111; // iC= 1759 
// vC = 14'b1111101010011100; // vC=-1380 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010101; // iC= 1685 
// vC = 14'b1111101001001101; // vC=-1459 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b1111101010000101; // vC=-1403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110001; // iC= 1777 
// vC = 14'b1111101010001100; // vC=-1396 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001011; // iC= 1675 
// vC = 14'b1111101011011111; // vC=-1313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101000; // iC= 1832 
// vC = 14'b1111101011111000; // vC=-1288 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110000; // iC= 1904 
// vC = 14'b1111101010001011; // vC=-1397 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100010; // iC= 1954 
// vC = 14'b1111101101111000; // vC=-1160 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111011; // iC= 1723 
// vC = 14'b1111101001110000; // vC=-1424 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010111; // iC= 1879 
// vC = 14'b1111101100000110; // vC=-1274 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b1111101101011111; // vC=-1185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101001; // iC= 1833 
// vC = 14'b1111101100011011; // vC=-1253 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101101; // iC= 1709 
// vC = 14'b1111101011101100; // vC=-1300 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b1111101011111000; // vC=-1288 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110100; // iC= 1716 
// vC = 14'b1111101101110100; // vC=-1164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111010; // iC= 1722 
// vC = 14'b1111101111010111; // vC=-1065 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111000; // iC= 1976 
// vC = 14'b1111101111000110; // vC=-1082 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b1111101011110001; // vC=-1295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100010; // iC= 1954 
// vC = 14'b1111101110001010; // vC=-1142 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b1111101011001111; // vC=-1329 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101110; // iC= 2030 
// vC = 14'b1111110000001010; // vC=-1014 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100101; // iC= 1765 
// vC = 14'b1111101011100001; // vC=-1311 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b1111110000010110; // vC=-1002 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b1111101011110100; // vC=-1292 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000001; // iC= 1921 
// vC = 14'b1111110000000000; // vC=-1024 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b1111101111100011; // vC=-1053 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101110; // iC= 2030 
// vC = 14'b1111101110101110; // vC=-1106 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111101110100001; // vC=-1119 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010100; // iC= 2068 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110000; // iC= 1840 
// vC = 14'b1111110000011100; // vC= -996 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b1111101111001010; // vC=-1078 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011110; // iC= 2078 
// vC = 14'b1111101111010000; // vC=-1072 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b1111101101110100; // vC=-1164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001001; // iC= 1993 
// vC = 14'b1111110000110000; // vC= -976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001000; // iC= 1992 
// vC = 14'b1111110000101001; // vC= -983 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001110; // iC= 1806 
// vC = 14'b1111101110011010; // vC=-1126 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101110; // iC= 1966 
// vC = 14'b1111110000011011; // vC= -997 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b1111110000010010; // vC=-1006 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100010; // iC= 2018 
// vC = 14'b1111110001100011; // vC= -925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000010; // iC= 2050 
// vC = 14'b1111110000000011; // vC=-1021 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b1111110000100110; // vC= -986 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110111; // iC= 1847 
// vC = 14'b1111110001100100; // vC= -924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b1111110010101101; // vC= -851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111101110111000; // vC=-1096 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000010; // iC= 1858 
// vC = 14'b1111110000110011; // vC= -973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b1111110010110000; // vC= -848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011111; // iC= 1887 
// vC = 14'b1111110011100011; // vC= -797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b1111110011001111; // vC= -817 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110100; // iC= 2100 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101110; // iC= 1902 
// vC = 14'b1111110011101111; // vC= -785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011111; // iC= 2079 
// vC = 14'b1111101111100011; // vC=-1053 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b1111110100000110; // vC= -762 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111110100001011; // vC= -757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100110; // iC= 1830 
// vC = 14'b1111110010000101; // vC= -891 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111110001110011; // vC= -909 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b1111101111111001; // vC=-1031 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b1111110010110111; // vC= -841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b1111110100101101; // vC= -723 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101010; // iC= 2090 
// vC = 14'b1111110100101010; // vC= -726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b1111110100101011; // vC= -725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010010; // iC= 1874 
// vC = 14'b1111110010000001; // vC= -895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011000; // iC= 1816 
// vC = 14'b1111110101001101; // vC= -691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b1111110010110010; // vC= -846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111111; // iC= 1983 
// vC = 14'b1111110100001111; // vC= -753 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111000; // iC= 1912 
// vC = 14'b1111110100011001; // vC= -743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b1111110101001101; // vC= -691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011110; // iC= 1822 
// vC = 14'b1111110001100011; // vC= -925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b1111110010001111; // vC= -881 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110000; // iC= 2032 
// vC = 14'b1111110100101100; // vC= -724 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010110; // iC= 2070 
// vC = 14'b1111110011100011; // vC= -797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001011; // iC= 1867 
// vC = 14'b1111110101111001; // vC= -647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111110011010101; // vC= -811 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111110011000000; // vC= -832 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000101; // iC= 1989 
// vC = 14'b1111110010101000; // vC= -856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b1111110110000111; // vC= -633 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b1111110011100011; // vC= -797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110101; // iC= 2037 
// vC = 14'b1111110110100110; // vC= -602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b1111110111100111; // vC= -537 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111100; // iC= 2108 
// vC = 14'b1111110100110000; // vC= -720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b1111110011100110; // vC= -794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110001; // iC= 1841 
// vC = 14'b1111110100101011; // vC= -725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b1111110110000111; // vC= -633 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010100; // iC= 1876 
// vC = 14'b1111111000000101; // vC= -507 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110110; // iC= 1910 
// vC = 14'b1111110100111011; // vC= -709 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001100; // iC= 2060 
// vC = 14'b1111110100010000; // vC= -752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110010; // iC= 2034 
// vC = 14'b1111110111000101; // vC= -571 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110100; // iC= 2100 
// vC = 14'b1111110101111001; // vC= -647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b1111110111110011; // vC= -525 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001000; // iC= 2120 
// vC = 14'b1111111001010111; // vC= -425 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010000; // iC= 2000 
// vC = 14'b1111111000010110; // vC= -490 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111110; // iC= 1982 
// vC = 14'b1111111000100000; // vC= -480 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b1111110101101011; // vC= -661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b1111111000101110; // vC= -466 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b1111110101000110; // vC= -698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b1111110111000011; // vC= -573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111111001111000; // vC= -392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110011; // iC= 2099 
// vC = 14'b1111111001011111; // vC= -417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011100; // iC= 2012 
// vC = 14'b1111110111001101; // vC= -563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b1111110111100101; // vC= -539 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101110; // iC= 2030 
// vC = 14'b1111111000101000; // vC= -472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111111010111101; // vC= -323 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b1111111010011111; // vC= -353 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001111; // iC= 2127 
// vC = 14'b1111111001111111; // vC= -385 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b1111110111010111; // vC= -553 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b1111111000100101; // vC= -475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010111; // iC= 1879 
// vC = 14'b1111110110101111; // vC= -593 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b1111111011100101; // vC= -283 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111000; // iC= 2104 
// vC = 14'b1111111010010111; // vC= -361 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111110111001100; // vC= -564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111101; // iC= 2045 
// vC = 14'b1111111011111000; // vC= -264 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b1111111100010001; // vC= -239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111000; // iC= 1912 
// vC = 14'b1111111010011110; // vC= -354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110101; // iC= 2037 
// vC = 14'b1111111100010011; // vC= -237 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011110; // iC= 2078 
// vC = 14'b1111111010111001; // vC= -327 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100001; // iC= 2017 
// vC = 14'b1111111000110101; // vC= -459 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111011; // iC= 1915 
// vC = 14'b1111111001001011; // vC= -437 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110111; // iC= 1847 
// vC = 14'b1111111010011001; // vC= -359 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b1111111011010010; // vC= -302 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100101; // iC= 1957 
// vC = 14'b1111111100100000; // vC= -224 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b1111111100010101; // vC= -235 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001000; // iC= 1864 
// vC = 14'b1111111100011010; // vC= -230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111000; // iC= 1976 
// vC = 14'b1111111001111010; // vC= -390 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111100; // iC= 2044 
// vC = 14'b1111111001111110; // vC= -386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b1111111101110111; // vC= -137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b1111111011011010; // vC= -294 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110010; // iC= 1842 
// vC = 14'b1111111010011000; // vC= -360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110011; // iC= 2099 
// vC = 14'b1111111001111110; // vC= -386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111010; // iC= 1850 
// vC = 14'b1111111011110101; // vC= -267 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001011; // iC= 1995 
// vC = 14'b1111111100000010; // vC= -254 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111000; // iC= 2104 
// vC = 14'b1111111011110101; // vC= -267 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b1111111001111100; // vC= -388 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111100; // iC= 2044 
// vC = 14'b1111111100010101; // vC= -235 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b1111111011010100; // vC= -300 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100000; // iC= 1824 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011110; // iC= 2078 
// vC = 14'b1111111101100100; // vC= -156 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101101; // iC= 2093 
// vC = 14'b1111111110101000; // vC=  -88 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110000; // iC= 1968 
// vC = 14'b1111111100011101; // vC= -227 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000011; // iC= 1923 
// vC = 14'b1111111111111011; // vC=   -5 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b1111111011111110; // vC= -258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011010; // iC= 1882 
// vC = 14'b1111111111101111; // vC=  -17 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b1111111111101011; // vC=  -21 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b1111111111000100; // vC=  -60 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b1111111110110111; // vC=  -73 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011011; // iC= 1947 
// vC = 14'b1111111101000011; // vC= -189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101001; // iC= 1833 
// vC = 14'b1111111110101001; // vC=  -87 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b1111111100101100; // vC= -212 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b1111111111100111; // vC=  -25 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b1111111110001010; // vC= -118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011000; // iC= 1816 
// vC = 14'b1111111110000111; // vC= -121 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001111; // iC= 1807 
// vC = 14'b0000000001000010; // vC=   66 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001101; // iC= 1869 
// vC = 14'b0000000001001100; // vC=   76 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011111; // iC= 2015 
// vC = 14'b1111111101011010; // vC= -166 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100000; // iC= 1824 
// vC = 14'b1111111101100111; // vC= -153 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001111; // iC= 1999 
// vC = 14'b0000000000010011; // vC=   19 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001101; // iC= 1869 
// vC = 14'b1111111111100100; // vC=  -28 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100011; // iC= 1955 
// vC = 14'b0000000000011011; // vC=   27 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b0000000001011100; // vC=   92 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110100; // iC= 1780 
// vC = 14'b0000000001101000; // vC=  104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b0000000000010100; // vC=   20 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101111; // iC= 1903 
// vC = 14'b0000000000110110; // vC=   54 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100110; // iC= 1766 
// vC = 14'b0000000010111000; // vC=  184 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101010; // iC= 1898 
// vC = 14'b0000000001011011; // vC=   91 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100110; // iC= 2022 
// vC = 14'b0000000001000111; // vC=   71 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b0000000001111011; // vC=  123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010101; // iC= 1749 
// vC = 14'b1111111111111110; // vC=   -2 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110101; // iC= 1845 
// vC = 14'b0000000010000100; // vC=  132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111001; // iC= 1849 
// vC = 14'b0000000011011100; // vC=  220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000000011101111; // vC=  239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100000; // iC= 1760 
// vC = 14'b0000000001001100; // vC=   76 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001101; // iC= 1741 
// vC = 14'b0000000010011010; // vC=  154 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011111; // iC= 2015 
// vC = 14'b0000000010101001; // vC=  169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b1111111111101101; // vC=  -19 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100000; // iC= 2016 
// vC = 14'b0000000001001010; // vC=   74 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111100; // iC= 2044 
// vC = 14'b0000000001011100; // vC=   92 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100110; // iC= 2022 
// vC = 14'b0000000011110011; // vC=  243 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100000; // iC= 2016 
// vC = 14'b0000000011000000; // vC=  192 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111000; // iC= 1784 
// vC = 14'b1111111111111101; // vC=   -3 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101001; // iC= 1897 
// vC = 14'b0000000101000101; // vC=  325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001110; // iC= 1934 
// vC = 14'b0000000011110100; // vC=  244 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111110; // iC= 1918 
// vC = 14'b0000000011111100; // vC=  252 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b0000000000110001; // vC=   49 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000100; // iC= 1924 
// vC = 14'b0000000010110100; // vC=  180 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b0000000001100000; // vC=   96 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000111; // iC= 1735 
// vC = 14'b0000000001101001; // vC=  105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110001; // iC= 1905 
// vC = 14'b0000000101010001; // vC=  337 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100111; // iC= 1831 
// vC = 14'b0000000101110111; // vC=  375 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110101; // iC= 1781 
// vC = 14'b0000000011110111; // vC=  247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100011; // iC= 1955 
// vC = 14'b0000000101110001; // vC=  369 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b0000000100110001; // vC=  305 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b0000000011000011; // vC=  195 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011101; // iC= 1821 
// vC = 14'b0000000001110000; // vC=  112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b0000000100111100; // vC=  316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111111; // iC= 1727 
// vC = 14'b0000000110001111; // vC=  399 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100011; // iC= 1891 
// vC = 14'b0000000110110000; // vC=  432 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010110; // iC= 1686 
// vC = 14'b0000000010110000; // vC=  176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b0000000110100010; // vC=  418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b0000000111010110; // vC=  470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101011; // iC= 1771 
// vC = 14'b0000000101011011; // vC=  347 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111100; // iC= 1852 
// vC = 14'b0000000101000100; // vC=  324 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111100; // iC= 1724 
// vC = 14'b0000000010110110; // vC=  182 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001000; // iC= 1736 
// vC = 14'b0000000101110110; // vC=  374 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b0000000101010011; // vC=  339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010001; // iC= 1681 
// vC = 14'b0000000011010110; // vC=  214 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000010; // iC= 1666 
// vC = 14'b0000000110000011; // vC=  387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b0000000100110000; // vC=  304 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001001; // iC= 1737 
// vC = 14'b0000000011101100; // vC=  236 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011000; // iC= 1752 
// vC = 14'b0000000100100111; // vC=  295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011101; // iC= 1821 
// vC = 14'b0000000011111001; // vC=  249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011010; // iC= 1690 
// vC = 14'b0000001000110101; // vC=  565 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b0000000101101010; // vC=  362 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001100; // iC= 1740 
// vC = 14'b0000000111111000; // vC=  504 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110011; // iC= 1779 
// vC = 14'b0000000110010000; // vC=  400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100000; // iC= 1888 
// vC = 14'b0000000101010010; // vC=  338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b0000000110111100; // vC=  444 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001111; // iC= 1807 
// vC = 14'b0000001001100100; // vC=  612 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000010; // iC= 1858 
// vC = 14'b0000000110100110; // vC=  422 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100010; // iC= 1890 
// vC = 14'b0000000110110010; // vC=  434 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b0000001001101001; // vC=  617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010110; // iC= 1878 
// vC = 14'b0000000101111000; // vC=  376 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111111; // iC= 1727 
// vC = 14'b0000001010001001; // vC=  649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101011; // iC= 1771 
// vC = 14'b0000000110100000; // vC=  416 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b0000001000001011; // vC=  523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011110; // iC= 1758 
// vC = 14'b0000000101110100; // vC=  372 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100000; // iC= 1824 
// vC = 14'b0000001000001100; // vC=  524 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110110; // iC= 1718 
// vC = 14'b0000001001011001; // vC=  601 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010111; // iC= 1623 
// vC = 14'b0000000111011011; // vC=  475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101011; // iC= 1707 
// vC = 14'b0000000110001100; // vC=  396 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101101; // iC= 1709 
// vC = 14'b0000001010110011; // vC=  691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011111; // iC= 1823 
// vC = 14'b0000001000110000; // vC=  560 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111100; // iC= 1724 
// vC = 14'b0000000111010100; // vC=  468 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010110; // iC= 1814 
// vC = 14'b0000001011100100; // vC=  740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011001; // iC= 1625 
// vC = 14'b0000001001011111; // vC=  607 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b0000001011011100; // vC=  732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010111; // iC= 1751 
// vC = 14'b0000001001110110; // vC=  630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111111; // iC= 1855 
// vC = 14'b0000000111000111; // vC=  455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001000; // iC= 1800 
// vC = 14'b0000001010110110; // vC=  694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111010; // iC= 1786 
// vC = 14'b0000001001110010; // vC=  626 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000000; // iC= 1600 
// vC = 14'b0000001011001110; // vC=  718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010001; // iC= 1681 
// vC = 14'b0000001011010101; // vC=  725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011111; // iC= 1695 
// vC = 14'b0000001011010111; // vC=  727 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101001; // iC= 1705 
// vC = 14'b0000001011011011; // vC=  731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110110; // iC= 1654 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111100; // iC= 1852 
// vC = 14'b0000001100001110; // vC=  782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001101; // iC= 1613 
// vC = 14'b0000001011110111; // vC=  759 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111100; // iC= 1596 
// vC = 14'b0000001001000101; // vC=  581 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001110; // iC= 1678 
// vC = 14'b0000001001000001; // vC=  577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101001; // iC= 1769 
// vC = 14'b0000001001111011; // vC=  635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110001; // iC= 1713 
// vC = 14'b0000001100100100; // vC=  804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011111; // iC= 1759 
// vC = 14'b0000001001010100; // vC=  596 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000110; // iC= 1670 
// vC = 14'b0000001001111100; // vC=  636 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111111; // iC= 1727 
// vC = 14'b0000001100110110; // vC=  822 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111110; // iC= 1662 
// vC = 14'b0000001011101110; // vC=  750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011111; // iC= 1823 
// vC = 14'b0000001010110011; // vC=  691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011101; // iC= 1693 
// vC = 14'b0000001010011010; // vC=  666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011100; // iC= 1820 
// vC = 14'b0000001100111001; // vC=  825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101111; // iC= 1775 
// vC = 14'b0000001100111100; // vC=  828 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001001; // iC= 1801 
// vC = 14'b0000001101101010; // vC=  874 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101001; // iC= 1513 
// vC = 14'b0000001010000101; // vC=  645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001000; // iC= 1736 
// vC = 14'b0000001010000110; // vC=  646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000100; // iC= 1604 
// vC = 14'b0000001101011011; // vC=  859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010001; // iC= 1809 
// vC = 14'b0000001011010000; // vC=  720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110100; // iC= 1524 
// vC = 14'b0000001101011100; // vC=  860 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011111; // iC= 1567 
// vC = 14'b0000001100011100; // vC=  796 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011001; // iC= 1689 
// vC = 14'b0000001111000101; // vC=  965 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010111; // iC= 1623 
// vC = 14'b0000001101011101; // vC=  861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000000; // iC= 1792 
// vC = 14'b0000001111010010; // vC=  978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101000; // iC= 1512 
// vC = 14'b0000001011111001; // vC=  761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101101; // iC= 1709 
// vC = 14'b0000001100000111; // vC=  775 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110111; // iC= 1591 
// vC = 14'b0000001111000111; // vC=  967 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001000; // iC= 1608 
// vC = 14'b0000001100001000; // vC=  776 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110111; // iC= 1719 
// vC = 14'b0000001011001011; // vC=  715 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100110; // iC= 1766 
// vC = 14'b0000001111110001; // vC= 1009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101011; // iC= 1451 
// vC = 14'b0000001111001010; // vC=  970 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010011; // iC= 1747 
// vC = 14'b0000001100101000; // vC=  808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000010; // iC= 1730 
// vC = 14'b0000001011011010; // vC=  730 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111001; // iC= 1529 
// vC = 14'b0000010000011111; // vC= 1055 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000101; // iC= 1605 
// vC = 14'b0000001101111010; // vC=  890 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110011; // iC= 1459 
// vC = 14'b0000001110001110; // vC=  910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010111; // iC= 1559 
// vC = 14'b0000001100010100; // vC=  788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000000; // iC= 1664 
// vC = 14'b0000001110011000; // vC=  920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010111; // iC= 1623 
// vC = 14'b0000010000110011; // vC= 1075 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111111; // iC= 1727 
// vC = 14'b0000010000000001; // vC= 1025 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000100; // iC= 1604 
// vC = 14'b0000001101011111; // vC=  863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001001; // iC= 1545 
// vC = 14'b0000010001000000; // vC= 1088 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010110; // iC= 1558 
// vC = 14'b0000001110110101; // vC=  949 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110110; // iC= 1462 
// vC = 14'b0000001111010111; // vC=  983 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000111; // iC= 1479 
// vC = 14'b0000001100110000; // vC=  816 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100100; // iC= 1508 
// vC = 14'b0000001111101100; // vC= 1004 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000100; // iC= 1412 
// vC = 14'b0000001111101001; // vC= 1001 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100010; // iC= 1506 
// vC = 14'b0000010001110100; // vC= 1140 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110101; // iC= 1525 
// vC = 14'b0000001101111011; // vC=  891 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100001; // iC= 1505 
// vC = 14'b0000010001011100; // vC= 1116 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000101; // iC= 1541 
// vC = 14'b0000001111001110; // vC=  974 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011001; // iC= 1369 
// vC = 14'b0000010000111010; // vC= 1082 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001001; // iC= 1417 
// vC = 14'b0000001111101010; // vC= 1002 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010000; // iC= 1360 
// vC = 14'b0000001101110111; // vC=  887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001010; // iC= 1674 
// vC = 14'b0000010010000100; // vC= 1156 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000101; // iC= 1477 
// vC = 14'b0000010000100011; // vC= 1059 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101100; // iC= 1644 
// vC = 14'b0000010010111000; // vC= 1208 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101110; // iC= 1646 
// vC = 14'b0000001111101111; // vC= 1007 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100011; // iC= 1635 
// vC = 14'b0000010010111001; // vC= 1209 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110111; // iC= 1463 
// vC = 14'b0000001110001010; // vC=  906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110000; // iC= 1328 
// vC = 14'b0000010000100100; // vC= 1060 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111111; // iC= 1535 
// vC = 14'b0000001111110001; // vC= 1009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110101; // iC= 1333 
// vC = 14'b0000010000011010; // vC= 1050 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001010; // iC= 1418 
// vC = 14'b0000001111011000; // vC=  984 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010111; // iC= 1367 
// vC = 14'b0000001110111100; // vC=  956 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001011; // iC= 1611 
// vC = 14'b0000001111000111; // vC=  967 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010010; // iC= 1618 
// vC = 14'b0000010001001110; // vC= 1102 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110000; // iC= 1456 
// vC = 14'b0000010011010110; // vC= 1238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100111; // iC= 1447 
// vC = 14'b0000010000101100; // vC= 1068 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011001; // iC= 1369 
// vC = 14'b0000010000010001; // vC= 1041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000100; // iC= 1540 
// vC = 14'b0000010010101010; // vC= 1194 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110110; // iC= 1462 
// vC = 14'b0000010011111000; // vC= 1272 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111100; // iC= 1404 
// vC = 14'b0000010100001011; // vC= 1291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010110; // iC= 1366 
// vC = 14'b0000010100001110; // vC= 1294 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000110; // iC= 1414 
// vC = 14'b0000010001101011; // vC= 1131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111011; // iC= 1403 
// vC = 14'b0000010011001101; // vC= 1229 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010101; // iC= 1493 
// vC = 14'b0000010000000010; // vC= 1026 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110001; // iC= 1265 
// vC = 14'b0000010001001111; // vC= 1103 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110110; // iC= 1270 
// vC = 14'b0000010100100101; // vC= 1317 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100011; // iC= 1443 
// vC = 14'b0000010100110000; // vC= 1328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010111; // iC= 1303 
// vC = 14'b0000010011001001; // vC= 1225 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011100; // iC= 1308 
// vC = 14'b0000010000011001; // vC= 1049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011110; // iC= 1438 
// vC = 14'b0000010000010101; // vC= 1045 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100100; // iC= 1508 
// vC = 14'b0000010011011111; // vC= 1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110101; // iC= 1525 
// vC = 14'b0000010011110001; // vC= 1265 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001000; // iC= 1416 
// vC = 14'b0000010101010100; // vC= 1364 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101111; // iC= 1263 
// vC = 14'b0000010001111111; // vC= 1151 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010000; // iC= 1360 
// vC = 14'b0000010011001110; // vC= 1230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011010; // iC= 1306 
// vC = 14'b0000010011101110; // vC= 1262 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000011; // iC= 1411 
// vC = 14'b0000010010100001; // vC= 1185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111010; // iC= 1338 
// vC = 14'b0000010101001100; // vC= 1356 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110010; // iC= 1394 
// vC = 14'b0000010100110011; // vC= 1331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011100; // iC= 1500 
// vC = 14'b0000010010101001; // vC= 1193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110101; // iC= 1461 
// vC = 14'b0000010101000010; // vC= 1346 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011000; // iC= 1304 
// vC = 14'b0000010001011111; // vC= 1119 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011001; // iC= 1305 
// vC = 14'b0000010101001000; // vC= 1352 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000011; // iC= 1283 
// vC = 14'b0000010010100100; // vC= 1188 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000111; // iC= 1159 
// vC = 14'b0000010101100100; // vC= 1380 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111010; // iC= 1210 
// vC = 14'b0000010101111100; // vC= 1404 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111101; // iC= 1149 
// vC = 14'b0000010011010101; // vC= 1237 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011001; // iC= 1177 
// vC = 14'b0000010110100010; // vC= 1442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100111; // iC= 1191 
// vC = 14'b0000010011010111; // vC= 1239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000000; // iC= 1216 
// vC = 14'b0000010110011011; // vC= 1435 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001010; // iC= 1418 
// vC = 14'b0000010100100100; // vC= 1316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111110; // iC= 1150 
// vC = 14'b0000010100011111; // vC= 1311 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110011; // iC= 1139 
// vC = 14'b0000010110110001; // vC= 1457 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110010; // iC= 1202 
// vC = 14'b0000010100011011; // vC= 1307 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001110; // iC= 1230 
// vC = 14'b0000010010011110; // vC= 1182 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010000; // iC= 1104 
// vC = 14'b0000010100000000; // vC= 1280 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111111; // iC= 1215 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000000; // iC= 1216 
// vC = 14'b0000010010110010; // vC= 1202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011101; // iC= 1117 
// vC = 14'b0000010101111110; // vC= 1406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111100; // iC= 1404 
// vC = 14'b0000010100000110; // vC= 1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010101; // iC= 1109 
// vC = 14'b0000010110011010; // vC= 1434 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101011; // iC= 1067 
// vC = 14'b0000010110011101; // vC= 1437 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001111; // iC= 1231 
// vC = 14'b0000010110001011; // vC= 1419 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001100; // iC= 1292 
// vC = 14'b0000010110100000; // vC= 1440 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001011; // iC= 1227 
// vC = 14'b0000010110111111; // vC= 1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000001; // iC= 1217 
// vC = 14'b0000010111010101; // vC= 1493 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101001; // iC= 1065 
// vC = 14'b0000010110001001; // vC= 1417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010101; // iC= 1237 
// vC = 14'b0000010100101101; // vC= 1325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110111; // iC= 1335 
// vC = 14'b0000010100000100; // vC= 1284 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001100; // iC= 1228 
// vC = 14'b0000010101010011; // vC= 1363 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001101; // iC= 1101 
// vC = 14'b0000010111010001; // vC= 1489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101001; // iC= 1193 
// vC = 14'b0000010100110010; // vC= 1330 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010100; // iC= 1044 
// vC = 14'b0000010011111111; // vC= 1279 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011011; // iC= 1115 
// vC = 14'b0000010011111010; // vC= 1274 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110010; // iC= 1010 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101001; // iC= 1065 
// vC = 14'b0000010100010110; // vC= 1302 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101001; // iC= 1065 
// vC = 14'b0000010100100111; // vC= 1319 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100010; // iC=  994 
// vC = 14'b0000011000010101; // vC= 1557 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110100; // iC= 1204 
// vC = 14'b0000010101001110; // vC= 1358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111100; // iC= 1020 
// vC = 14'b0000011000101010; // vC= 1578 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010000; // iC= 1040 
// vC = 14'b0000010110110100; // vC= 1460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001110; // iC= 1038 
// vC = 14'b0000011001010111; // vC= 1623 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000001; // iC= 1281 
// vC = 14'b0000010110101100; // vC= 1452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100000; // iC=  992 
// vC = 14'b0000011001100110; // vC= 1638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010010; // iC= 1106 
// vC = 14'b0000010110110100; // vC= 1460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101111; // iC= 1263 
// vC = 14'b0000010110001011; // vC= 1419 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010110; // iC= 1110 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111010; // iC= 1146 
// vC = 14'b0000010110101110; // vC= 1454 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001011; // iC= 1099 
// vC = 14'b0000011000010110; // vC= 1558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100110; // iC= 1062 
// vC = 14'b0000010101110010; // vC= 1394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001101; // iC= 1101 
// vC = 14'b0000010101110110; // vC= 1398 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001001; // iC= 1225 
// vC = 14'b0000011000100001; // vC= 1569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011101; // iC= 1053 
// vC = 14'b0000011001000110; // vC= 1606 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101000; // iC= 1000 
// vC = 14'b0000010101110000; // vC= 1392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101011; // iC=  939 
// vC = 14'b0000010111111111; // vC= 1535 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011100; // iC= 1052 
// vC = 14'b0000011000110011; // vC= 1587 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010101; // iC=  917 
// vC = 14'b0000011000001001; // vC= 1545 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011100; // iC= 1180 
// vC = 14'b0000011001101010; // vC= 1642 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100010; // iC=  994 
// vC = 14'b0000011000100111; // vC= 1575 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101111; // iC= 1071 
// vC = 14'b0000010111110010; // vC= 1522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110100; // iC= 1140 
// vC = 14'b0000011000101100; // vC= 1580 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000001; // iC= 1153 
// vC = 14'b0000011000011111; // vC= 1567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001000; // iC=  968 
// vC = 14'b0000011010001101; // vC= 1677 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111110; // iC= 1150 
// vC = 14'b0000010110000000; // vC= 1408 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101110; // iC= 1070 
// vC = 14'b0000010110010010; // vC= 1426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001000; // iC=  968 
// vC = 14'b0000010110000100; // vC= 1412 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000111; // iC= 1095 
// vC = 14'b0000011001101101; // vC= 1645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111111; // iC=  831 
// vC = 14'b0000011010010100; // vC= 1684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110011; // iC=  883 
// vC = 14'b0000011010000100; // vC= 1668 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110101; // iC=  949 
// vC = 14'b0000011011010101; // vC= 1749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000010; // iC= 1026 
// vC = 14'b0000010111111001; // vC= 1529 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001011; // iC=  971 
// vC = 14'b0000011000111110; // vC= 1598 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010010; // iC= 1106 
// vC = 14'b0000011001010110; // vC= 1622 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010100; // iC=  788 
// vC = 14'b0000011000110010; // vC= 1586 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110100; // iC= 1012 
// vC = 14'b0000011001010101; // vC= 1621 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000100; // iC= 1028 
// vC = 14'b0000011010101001; // vC= 1705 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101101; // iC=  877 
// vC = 14'b0000010110111101; // vC= 1469 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000111; // iC=  775 
// vC = 14'b0000011010011001; // vC= 1689 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100100; // iC=  932 
// vC = 14'b0000011001011010; // vC= 1626 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100000; // iC=  864 
// vC = 14'b0000011011101111; // vC= 1775 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011011; // iC=  859 
// vC = 14'b0000011010000010; // vC= 1666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100111; // iC=  999 
// vC = 14'b0000010111110111; // vC= 1527 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101000; // iC=  936 
// vC = 14'b0000010111011111; // vC= 1503 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110100; // iC=  948 
// vC = 14'b0000011010110011; // vC= 1715 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011001; // iC=  985 
// vC = 14'b0000011010010111; // vC= 1687 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100010; // iC=  802 
// vC = 14'b0000011011001110; // vC= 1742 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000000; // iC=  832 
// vC = 14'b0000011000101111; // vC= 1583 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111100; // iC=  764 
// vC = 14'b0000011100010101; // vC= 1813 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010000; // iC=  912 
// vC = 14'b0000011010111000; // vC= 1720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110101; // iC=  821 
// vC = 14'b0000011010000000; // vC= 1664 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011001; // iC=  921 
// vC = 14'b0000010111111100; // vC= 1532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111101; // iC=  893 
// vC = 14'b0000011000111111; // vC= 1599 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110010; // iC=  754 
// vC = 14'b0000011000100000; // vC= 1568 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011011; // iC=  987 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110110; // iC=  694 
// vC = 14'b0000011000110100; // vC= 1588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110011; // iC=  755 
// vC = 14'b0000011001101101; // vC= 1645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111001; // iC=  889 
// vC = 14'b0000011001011100; // vC= 1628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110011; // iC=  691 
// vC = 14'b0000011000010011; // vC= 1555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001111; // iC=  911 
// vC = 14'b0000011100110010; // vC= 1842 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001010; // iC=  650 
// vC = 14'b0000011001011111; // vC= 1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001111; // iC=  847 
// vC = 14'b0000011010101001; // vC= 1705 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110011; // iC=  627 
// vC = 14'b0000011100011001; // vC= 1817 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101111; // iC=  623 
// vC = 14'b0000011001010111; // vC= 1623 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011111; // iC=  799 
// vC = 14'b0000011010001010; // vC= 1674 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111110; // iC=  894 
// vC = 14'b0000011010001001; // vC= 1673 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111110; // iC=  702 
// vC = 14'b0000011000010001; // vC= 1553 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110000; // iC=  624 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110000; // iC=  752 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000001; // iC=  769 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110110; // iC=  886 
// vC = 14'b0000011000101100; // vC= 1580 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110000; // iC=  688 
// vC = 14'b0000011000101001; // vC= 1577 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111100; // iC=  764 
// vC = 14'b0000011010110101; // vC= 1717 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111110; // iC=  638 
// vC = 14'b0000011011110110; // vC= 1782 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100101; // iC=  741 
// vC = 14'b0000011100101101; // vC= 1837 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001100; // iC=  716 
// vC = 14'b0000011100011100; // vC= 1820 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110011; // iC=  627 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100001; // iC=  801 
// vC = 14'b0000011010000101; // vC= 1669 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110001; // iC=  817 
// vC = 14'b0000011101011101; // vC= 1885 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111001; // iC=  825 
// vC = 14'b0000011100100110; // vC= 1830 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101001; // iC=  681 
// vC = 14'b0000011011101111; // vC= 1775 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010111; // iC=  599 
// vC = 14'b0000011010001110; // vC= 1678 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110001; // iC=  753 
// vC = 14'b0000011010001110; // vC= 1678 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110101; // iC=  501 
// vC = 14'b0000011011010000; // vC= 1744 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110111; // iC=  567 
// vC = 14'b0000011010010010; // vC= 1682 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011101; // iC=  605 
// vC = 14'b0000011001000001; // vC= 1601 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111101; // iC=  445 
// vC = 14'b0000011001110010; // vC= 1650 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011000; // iC=  472 
// vC = 14'b0000011100110110; // vC= 1846 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010110; // iC=  534 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011110; // iC=  734 
// vC = 14'b0000011010001000; // vC= 1672 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111011; // iC=  507 
// vC = 14'b0000011110000101; // vC= 1925 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101000; // iC=  552 
// vC = 14'b0000011011100110; // vC= 1766 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101011; // iC=  491 
// vC = 14'b0000011001011010; // vC= 1626 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001011; // iC=  587 
// vC = 14'b0000011100010010; // vC= 1810 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001111; // iC=  655 
// vC = 14'b0000011100000110; // vC= 1798 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011111; // iC=  543 
// vC = 14'b0000011101100011; // vC= 1891 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000001; // iC=  321 
// vC = 14'b0000011100111000; // vC= 1848 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001100; // iC=  332 
// vC = 14'b0000011011011110; // vC= 1758 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010110; // iC=  598 
// vC = 14'b0000011110001001; // vC= 1929 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010111; // iC=  535 
// vC = 14'b0000011010011010; // vC= 1690 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111110; // iC=  382 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111000; // iC=  504 
// vC = 14'b0000011010000101; // vC= 1669 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110110; // iC=  374 
// vC = 14'b0000011001100100; // vC= 1636 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000001; // iC=  513 
// vC = 14'b0000011010011000; // vC= 1688 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111001; // iC=  249 
// vC = 14'b0000011100100101; // vC= 1829 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001011; // iC=  203 
// vC = 14'b0000011100111100; // vC= 1852 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100111; // iC=  295 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111111; // iC=  191 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111011; // iC=  315 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101010; // iC=  234 
// vC = 14'b0000011101111000; // vC= 1912 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100110; // iC=  294 
// vC = 14'b0000011100101000; // vC= 1832 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001110; // iC=  398 
// vC = 14'b0000011010001000; // vC= 1672 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110111; // iC=  311 
// vC = 14'b0000011010110111; // vC= 1719 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000100; // iC=  260 
// vC = 14'b0000011101001100; // vC= 1868 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100011; // iC=   99 
// vC = 14'b0000011100010010; // vC= 1810 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010101; // iC=  277 
// vC = 14'b0000011010100001; // vC= 1697 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101100; // iC=   44 
// vC = 14'b0000011100100010; // vC= 1826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100100; // iC=  164 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100100; // iC=   36 
// vC = 14'b0000011100001010; // vC= 1802 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001101; // iC=  141 
// vC = 14'b0000011101001111; // vC= 1871 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001110; // iC=   14 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111000; // iC=  184 
// vC = 14'b0000011110100011; // vC= 1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000001; // iC=    1 
// vC = 14'b0000011101001100; // vC= 1868 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000100; // iC=  196 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010111; // iC=   23 
// vC = 14'b0000011101101111; // vC= 1903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100010; // iC=  -30 
// vC = 14'b0000011101100011; // vC= 1891 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111111; // iC=  127 
// vC = 14'b0000011011000010; // vC= 1730 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100011; // iC= -157 
// vC = 14'b0000011011110101; // vC= 1781 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011000; // iC=   24 
// vC = 14'b0000011011100100; // vC= 1764 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100011; // iC=   35 
// vC = 14'b0000011010111000; // vC= 1720 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001100; // iC= -116 
// vC = 14'b0000011010010001; // vC= 1681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010110; // iC= -234 
// vC = 14'b0000011010110111; // vC= 1719 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111000; // iC=   -8 
// vC = 14'b0000011101010010; // vC= 1874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000110; // iC=    6 
// vC = 14'b0000011101010101; // vC= 1877 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011110; // iC= -226 
// vC = 14'b0000011010100001; // vC= 1697 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101000; // iC= -280 
// vC = 14'b0000011101000100; // vC= 1860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111010; // iC= -134 
// vC = 14'b0000011010101011; // vC= 1707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110111; // iC= -329 
// vC = 14'b0000011101101010; // vC= 1898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111010; // iC= -390 
// vC = 14'b0000011110010001; // vC= 1937 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100010; // iC= -222 
// vC = 14'b0000011001100111; // vC= 1639 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000010; // iC= -254 
// vC = 14'b0000011110011111; // vC= 1951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111001; // iC= -327 
// vC = 14'b0000011010111101; // vC= 1725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101110; // iC= -402 
// vC = 14'b0000011010010010; // vC= 1682 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010010; // iC= -430 
// vC = 14'b0000011110000101; // vC= 1925 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100111; // iC= -409 
// vC = 14'b0000011011101111; // vC= 1775 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011110; // iC= -354 
// vC = 14'b0000011101001001; // vC= 1865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011011; // iC= -485 
// vC = 14'b0000011010000100; // vC= 1668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010000; // iC= -304 
// vC = 14'b0000011101100111; // vC= 1895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010100; // iC= -364 
// vC = 14'b0000011100001010; // vC= 1802 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011011; // iC= -421 
// vC = 14'b0000011001010001; // vC= 1617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100001; // iC= -479 
// vC = 14'b0000011100001000; // vC= 1800 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000010; // iC= -638 
// vC = 14'b0000011101000010; // vC= 1858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010011; // iC= -557 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001101; // iC= -627 
// vC = 14'b0000011101110101; // vC= 1909 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010101; // iC= -619 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001011; // iC= -501 
// vC = 14'b0000011011011000; // vC= 1752 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101111; // iC= -785 
// vC = 14'b0000011101000100; // vC= 1860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000011; // iC= -637 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111110; // iC= -642 
// vC = 14'b0000011100001000; // vC= 1800 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000100; // iC= -828 
// vC = 14'b0000011010000100; // vC= 1668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111010; // iC= -838 
// vC = 14'b0000011011100111; // vC= 1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b0000011100111111; // vC= 1855 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000111; // iC= -825 
// vC = 14'b0000011011101001; // vC= 1769 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110000; // iC= -784 
// vC = 14'b0000011010110011; // vC= 1715 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010101; // iC= -939 
// vC = 14'b0000011011010010; // vC= 1746 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011001; // iC= -743 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101011; // iC= -725 
// vC = 14'b0000011101011001; // vC= 1881 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110000; // iC= -784 
// vC = 14'b0000011000111101; // vC= 1597 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001000; // iC= -824 
// vC = 14'b0000011011000001; // vC= 1729 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011100; // iC= -868 
// vC = 14'b0000011000111101; // vC= 1597 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111001; // iC= -967 
// vC = 14'b0000011101001101; // vC= 1869 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000111; // iC=-1145 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100000; // iC=-1056 
// vC = 14'b0000011100101110; // vC= 1838 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000100; // iC=-1084 
// vC = 14'b0000011001000110; // vC= 1606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100000; // iC=-1184 
// vC = 14'b0000011100110000; // vC= 1840 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001010; // iC=-1078 
// vC = 14'b0000011001101111; // vC= 1647 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101110; // iC=-1106 
// vC = 14'b0000011001000010; // vC= 1602 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010100; // iC=-1068 
// vC = 14'b0000010111111011; // vC= 1531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100011; // iC= -989 
// vC = 14'b0000011011110001; // vC= 1777 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100111; // iC=-1113 
// vC = 14'b0000011011001110; // vC= 1742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111000; // iC=-1032 
// vC = 14'b0000011000110011; // vC= 1587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110001; // iC=-1167 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001100; // iC=-1076 
// vC = 14'b0000011000101111; // vC= 1583 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001010; // iC=-1270 
// vC = 14'b0000011001100000; // vC= 1632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110100; // iC=-1292 
// vC = 14'b0000011000011111; // vC= 1567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000000; // iC=-1280 
// vC = 14'b0000011001001100; // vC= 1612 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010101; // iC=-1259 
// vC = 14'b0000010111000010; // vC= 1474 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111101; // iC=-1155 
// vC = 14'b0000010110111011; // vC= 1467 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100100; // iC=-1180 
// vC = 14'b0000011000110110; // vC= 1590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101000; // iC=-1368 
// vC = 14'b0000011001000101; // vC= 1605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000100; // iC=-1404 
// vC = 14'b0000011001111010; // vC= 1658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101011; // iC=-1493 
// vC = 14'b0000010111110010; // vC= 1522 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001011; // iC=-1269 
// vC = 14'b0000011010011110; // vC= 1694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110001; // iC=-1359 
// vC = 14'b0000010110101001; // vC= 1449 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000110; // iC=-1402 
// vC = 14'b0000011000110011; // vC= 1587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010101; // iC=-1387 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010010; // iC=-1390 
// vC = 14'b0000011010010001; // vC= 1681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000110; // iC=-1466 
// vC = 14'b0000011001000101; // vC= 1605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101001; // iC=-1303 
// vC = 14'b0000010111000101; // vC= 1477 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110010; // iC=-1358 
// vC = 14'b0000010101101100; // vC= 1388 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101010; // iC=-1366 
// vC = 14'b0000011000111110; // vC= 1598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000111; // iC=-1401 
// vC = 14'b0000011000110000; // vC= 1584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111010; // iC=-1606 
// vC = 14'b0000011010010011; // vC= 1683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101101; // iC=-1491 
// vC = 14'b0000010111000111; // vC= 1479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010100; // iC=-1452 
// vC = 14'b0000011001101101; // vC= 1645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100100; // iC=-1564 
// vC = 14'b0000010101111111; // vC= 1407 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001100; // iC=-1716 
// vC = 14'b0000011000011000; // vC= 1560 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101100; // iC=-1492 
// vC = 14'b0000011001010011; // vC= 1619 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010100; // iC=-1644 
// vC = 14'b0000010101011011; // vC= 1371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000001; // iC=-1535 
// vC = 14'b0000010110111101; // vC= 1469 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000111; // iC=-1657 
// vC = 14'b0000011000000010; // vC= 1538 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001010; // iC=-1718 
// vC = 14'b0000010110110011; // vC= 1459 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110100; // iC=-1804 
// vC = 14'b0000010111000010; // vC= 1474 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111000; // iC=-1608 
// vC = 14'b0000010101100010; // vC= 1378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010100; // iC=-1580 
// vC = 14'b0000010111011110; // vC= 1502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110111; // iC=-1609 
// vC = 14'b0000010110011010; // vC= 1434 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000001; // iC=-1791 
// vC = 14'b0000010011110111; // vC= 1271 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100001; // iC=-1567 
// vC = 14'b0000010110101010; // vC= 1450 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100010; // iC=-1566 
// vC = 14'b0000010101101100; // vC= 1388 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100101; // iC=-1819 
// vC = 14'b0000010100100001; // vC= 1313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011001; // iC=-1639 
// vC = 14'b0000010011111000; // vC= 1272 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b0000010100100001; // vC= 1313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110100; // iC=-1804 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010011; // iC=-1645 
// vC = 14'b0000010110100001; // vC= 1441 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b0000010111101100; // vC= 1516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011101; // iC=-1699 
// vC = 14'b0000010011100110; // vC= 1254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110001; // iC=-1807 
// vC = 14'b0000010100111011; // vC= 1339 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000010; // iC=-1726 
// vC = 14'b0000010100110111; // vC= 1335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110010; // iC=-1742 
// vC = 14'b0000010101101101; // vC= 1389 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b0000010110101100; // vC= 1452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111101; // iC=-1731 
// vC = 14'b0000010100100001; // vC= 1313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110011; // iC=-1869 
// vC = 14'b0000010011000000; // vC= 1216 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011111; // iC=-1697 
// vC = 14'b0000010100111111; // vC= 1343 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100000; // iC=-1824 
// vC = 14'b0000010011101100; // vC= 1260 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b0000010101010110; // vC= 1366 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001101; // iC=-1715 
// vC = 14'b0000010011110101; // vC= 1269 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010001; // iC=-1839 
// vC = 14'b0000010100001110; // vC= 1294 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111101; // iC=-1923 
// vC = 14'b0000010001001101; // vC= 1101 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b0000010010101111; // vC= 1199 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110101; // iC=-1803 
// vC = 14'b0000010001010000; // vC= 1104 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b0000010101011101; // vC= 1373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001111; // iC=-1841 
// vC = 14'b0000010011101111; // vC= 1263 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110000; // iC=-2000 
// vC = 14'b0000010100010011; // vC= 1299 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001111; // iC=-1777 
// vC = 14'b0000010010000101; // vC= 1157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b0000010001000010; // vC= 1090 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100011; // iC=-1757 
// vC = 14'b0000010100011011; // vC= 1307 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110010; // iC=-1806 
// vC = 14'b0000010000101011; // vC= 1067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010111; // iC=-1897 
// vC = 14'b0000010100100101; // vC= 1317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b0000010010000100; // vC= 1156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b0000010000010100; // vC= 1044 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b0000010001101001; // vC= 1129 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b0000010010011110; // vC= 1182 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111010; // iC=-1798 
// vC = 14'b0000010001100001; // vC= 1121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b0000010001000000; // vC= 1088 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010000; // iC=-2096 
// vC = 14'b0000010010101111; // vC= 1199 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b0000010010100001; // vC= 1185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100111; // iC=-1817 
// vC = 14'b0000001111000000; // vC=  960 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b0000001110011100; // vC=  924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010110; // iC=-2026 
// vC = 14'b0000001110101100; // vC=  940 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010110; // iC=-2090 
// vC = 14'b0000010001001111; // vC= 1103 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010100; // iC=-1900 
// vC = 14'b0000001111000111; // vC=  967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100010; // iC=-1886 
// vC = 14'b0000010001011001; // vC= 1113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101000; // iC=-1880 
// vC = 14'b0000001111000101; // vC=  965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101010; // iC=-1814 
// vC = 14'b0000001111111111; // vC= 1023 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b0000010000000011; // vC= 1027 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110110; // iC=-1994 
// vC = 14'b0000010001011110; // vC= 1118 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111111; // iC=-1985 
// vC = 14'b0000010001011011; // vC= 1115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b0000001111000101; // vC=  965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b0000001111011100; // vC=  988 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000010001110111; // vC= 1143 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b0000001110110001; // vC=  945 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b0000001111010110; // vC=  982 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001011; // iC=-1973 
// vC = 14'b0000010000010111; // vC= 1047 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b0000010000001101; // vC= 1037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111001; // iC=-1927 
// vC = 14'b0000001100111001; // vC=  825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010110; // iC=-1834 
// vC = 14'b0000010000110010; // vC= 1074 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b0000001101001011; // vC=  843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011010; // iC=-1830 
// vC = 14'b0000010000011001; // vC= 1049 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b0000010000001000; // vC= 1032 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011001; // iC=-1895 
// vC = 14'b0000001011111110; // vC=  766 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b0000001100011011; // vC=  795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010110; // iC=-2026 
// vC = 14'b0000001101101100; // vC=  876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000010; // iC=-1854 
// vC = 14'b0000001110101101; // vC=  941 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000100; // iC=-1980 
// vC = 14'b0000001110011010; // vC=  922 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b0000001010110010; // vC=  690 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b0000001111001011; // vC=  971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011000; // iC=-1896 
// vC = 14'b0000001101011100; // vC=  860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010100; // iC=-2092 
// vC = 14'b0000001110001100; // vC=  908 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010000; // iC=-1968 
// vC = 14'b0000001011011111; // vC=  735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b0000001110011011; // vC=  923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b0000001101001000; // vC=  840 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b0000001001110100; // vC=  628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111001; // iC=-1863 
// vC = 14'b0000001100001010; // vC=  778 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010010; // iC=-2094 
// vC = 14'b0000001010100110; // vC=  678 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b0000001011001011; // vC=  715 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010110; // iC=-1834 
// vC = 14'b0000001100111101; // vC=  829 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101110; // iC=-1874 
// vC = 14'b0000001011011010; // vC=  730 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b0000001001001001; // vC=  585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000001011001000; // vC=  712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100100; // iC=-2140 
// vC = 14'b0000001100011000; // vC=  792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000111; // iC=-1977 
// vC = 14'b0000001010011100; // vC=  668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b0000001000010011; // vC=  531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b0000001010111000; // vC=  696 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001111; // iC=-1905 
// vC = 14'b0000001000101110; // vC=  558 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110011; // iC=-1869 
// vC = 14'b0000001010101011; // vC=  683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010111; // iC=-1961 
// vC = 14'b0000001000110000; // vC=  560 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011011; // iC=-1829 
// vC = 14'b0000001011000100; // vC=  708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b0000001011011001; // vC=  729 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000110; // iC=-1914 
// vC = 14'b0000001001100110; // vC=  614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000001010101111; // vC=  687 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001111; // iC=-1841 
// vC = 14'b0000001001001000; // vC=  584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000000111011111; // vC=  479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111011; // iC=-2117 
// vC = 14'b0000001010011000; // vC=  664 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b0000000111001110; // vC=  462 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100100; // iC=-1820 
// vC = 14'b0000001000011100; // vC=  540 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011110; // iC=-2018 
// vC = 14'b0000001011001011; // vC=  715 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111110; // iC=-1922 
// vC = 14'b0000001000010011; // vC=  531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100011; // iC=-1821 
// vC = 14'b0000001000001111; // vC=  527 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010000; // iC=-1904 
// vC = 14'b0000001001111010; // vC=  634 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b0000000110000110; // vC=  390 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101111; // iC=-2001 
// vC = 14'b0000000110111110; // vC=  446 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000000101110000; // vC=  368 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b0000001001010011; // vC=  595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b0000000110100000; // vC=  416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b0000001001000110; // vC=  582 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100100; // iC=-1948 
// vC = 14'b0000000101100111; // vC=  359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001001; // iC=-2103 
// vC = 14'b0000000101111010; // vC=  378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b0000001000110000; // vC=  560 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110010; // iC=-1934 
// vC = 14'b0000001001010110; // vC=  598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b0000000100100000; // vC=  288 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010000; // iC=-2096 
// vC = 14'b0000000101000111; // vC=  327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b0000001000010001; // vC=  529 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001000; // iC=-2040 
// vC = 14'b0000000110100111; // vC=  423 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000000111110110; // vC=  502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110010; // iC=-1870 
// vC = 14'b0000001000011001; // vC=  537 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110001; // iC=-1871 
// vC = 14'b0000000111011110; // vC=  478 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000010; // iC=-1854 
// vC = 14'b0000000110110101; // vC=  437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b0000000111110010; // vC=  498 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b0000001000001111; // vC=  527 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b0000000110100011; // vC=  419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b0000000111110111; // vC=  503 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b0000000110110100; // vC=  436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b0000000100101101; // vC=  301 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111001; // iC=-2119 
// vC = 14'b0000000111010101; // vC=  469 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110011; // iC=-1997 
// vC = 14'b0000000011011011; // vC=  219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000000110000110; // vC=  390 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b0000000111001111; // vC=  463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b0000000011110010; // vC=  242 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000000101000101; // vC=  325 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000000011000010; // vC=  194 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001001; // iC=-1847 
// vC = 14'b0000000010111110; // vC=  190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b0000000011011011; // vC=  219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000000001011111; // vC=   95 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111001; // iC=-1863 
// vC = 14'b0000000101101101; // vC=  365 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001010; // iC=-1910 
// vC = 14'b0000000001001110; // vC=   78 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111000; // iC=-2120 
// vC = 14'b0000000100101000; // vC=  296 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000000011110110; // vC=  246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000000001011101; // vC=   93 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000000001010110; // vC=   86 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b0000000011101101; // vC=  237 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b0000000010001001; // vC=  137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100110; // iC=-1818 
// vC = 14'b0000000001001010; // vC=   74 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b0000000001110111; // vC=  119 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b0000000010101100; // vC=  172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010110; // iC=-1834 
// vC = 14'b1111111111110110; // vC=  -10 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b0000000010011101; // vC=  157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111001; // iC=-1991 
// vC = 14'b0000000100011000; // vC=  280 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110011; // iC=-1933 
// vC = 14'b0000000011001011; // vC=  203 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b0000000000101001; // vC=   41 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b0000000011011011; // vC=  219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b1111111111010010; // vC=  -46 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b0000000001000011; // vC=   67 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100100; // iC=-1948 
// vC = 14'b1111111111001100; // vC=  -52 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101111; // iC=-1809 
// vC = 14'b0000000000110010; // vC=   50 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b0000000011010111; // vC=  215 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001001; // iC=-1847 
// vC = 14'b0000000000011110; // vC=   30 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001110; // iC=-1842 
// vC = 14'b0000000001001000; // vC=   72 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b0000000001101111; // vC=  111 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b0000000001001001; // vC=   73 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b0000000001110010; // vC=  114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100101; // iC=-2075 
// vC = 14'b1111111111000111; // vC=  -57 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000011; // iC=-1853 
// vC = 14'b1111111111111000; // vC=   -8 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010000; // iC=-1904 
// vC = 14'b0000000010011011; // vC=  155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111110; // iC=-1794 
// vC = 14'b1111111101100100; // vC= -156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b1111111110111011; // vC=  -69 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b1111111111111010; // vC=   -6 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110010; // iC=-2062 
// vC = 14'b1111111110000001; // vC= -127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011110; // iC=-1826 
// vC = 14'b1111111100111110; // vC= -194 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100111; // iC=-1817 
// vC = 14'b1111111111001010; // vC=  -54 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010001; // iC=-1839 
// vC = 14'b1111111110011110; // vC=  -98 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100111; // iC=-1753 
// vC = 14'b1111111101010111; // vC= -169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b1111111101001011; // vC= -181 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b1111111111001001; // vC=  -55 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b1111111100000001; // vC= -255 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b1111111101111000; // vC= -136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011110; // iC=-2018 
// vC = 14'b1111111101100110; // vC= -154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101111; // iC=-2001 
// vC = 14'b1111111100000111; // vC= -249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011101; // iC=-1827 
// vC = 14'b0000000000010001; // vC=   17 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b1111111111110100; // vC=  -12 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111101; // iC=-1795 
// vC = 14'b1111111100000100; // vC= -252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b1111111111001001; // vC=  -55 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001010; // iC=-1846 
// vC = 14'b1111111100100110; // vC= -218 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010110; // iC=-1770 
// vC = 14'b1111111100011111; // vC= -225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b1111111111010001; // vC=  -47 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010001; // iC=-2031 
// vC = 14'b1111111111000110; // vC=  -58 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b1111111010100111; // vC= -345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001010; // iC=-1782 
// vC = 14'b1111111101111000; // vC= -136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b1111111100101010; // vC= -214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001100; // iC=-1780 
// vC = 14'b1111111110000000; // vC= -128 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000111; // iC=-1977 
// vC = 14'b1111111001111110; // vC= -386 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011000; // iC=-1896 
// vC = 14'b1111111011000000; // vC= -320 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b1111111010101011; // vC= -341 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b1111111100001010; // vC= -246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010111; // iC=-1897 
// vC = 14'b1111111001101110; // vC= -402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010111; // iC=-1833 
// vC = 14'b1111111001101100; // vC= -404 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b1111111010110111; // vC= -329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101010; // iC=-1814 
// vC = 14'b1111111110001100; // vC= -116 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b1111111001110111; // vC= -393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101111; // iC=-1809 
// vC = 14'b1111111001101010; // vC= -406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111010; // iC=-1798 
// vC = 14'b1111111011001101; // vC= -307 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111101; // iC=-1795 
// vC = 14'b1111111100001101; // vC= -243 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b1111111101010010; // vC= -174 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001010; // iC=-1718 
// vC = 14'b1111111001101101; // vC= -403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000101; // iC=-1915 
// vC = 14'b1111111010110001; // vC= -335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110100; // iC=-1932 
// vC = 14'b1111111010101100; // vC= -340 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110001; // iC=-1743 
// vC = 14'b1111111100100111; // vC= -217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b1111111000101011; // vC= -469 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111000; // iC=-1800 
// vC = 14'b1111111010111010; // vC= -326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b1111111011111000; // vC= -264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010001; // iC=-1775 
// vC = 14'b1111111001010100; // vC= -428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101011; // iC=-1749 
// vC = 14'b1111111100011111; // vC= -225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000100; // iC=-1788 
// vC = 14'b1111111000001111; // vC= -497 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101011; // iC=-1877 
// vC = 14'b1111111000000001; // vC= -511 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110010; // iC=-1806 
// vC = 14'b1111111100000111; // vC= -249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001011; // iC=-1653 
// vC = 14'b1111111010110000; // vC= -336 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000101; // iC=-1915 
// vC = 14'b1111111010100111; // vC= -345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011100; // iC=-1700 
// vC = 14'b1111111010010110; // vC= -362 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100110; // iC=-1690 
// vC = 14'b1111110111011100; // vC= -548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b1111111010000101; // vC= -379 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011000; // iC=-1704 
// vC = 14'b1111111010100111; // vC= -345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000101; // iC=-1659 
// vC = 14'b1111111010011100; // vC= -356 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110001; // iC=-1935 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000010; // iC=-1790 
// vC = 14'b1111111001010100; // vC= -428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011110; // iC=-1762 
// vC = 14'b1111110111101100; // vC= -532 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b1111110101110100; // vC= -652 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000001; // iC=-1663 
// vC = 14'b1111110111110000; // vC= -528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b1111111000001010; // vC= -502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110000; // iC=-1616 
// vC = 14'b1111111000001001; // vC= -503 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b1111110111001001; // vC= -567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b1111110101110100; // vC= -652 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b1111110101001010; // vC= -694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010001; // iC=-1647 
// vC = 14'b1111110111010011; // vC= -557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001001; // iC=-1655 
// vC = 14'b1111110101000010; // vC= -702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b1111111000111010; // vC= -454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110111; // iC=-1609 
// vC = 14'b1111111000011010; // vC= -486 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101101; // iC=-1619 
// vC = 14'b1111111000010011; // vC= -493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011100; // iC=-1636 
// vC = 14'b1111110111010110; // vC= -554 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101101; // iC=-1683 
// vC = 14'b1111111000101101; // vC= -467 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010110; // iC=-1706 
// vC = 14'b1111110110001100; // vC= -628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100010; // iC=-1822 
// vC = 14'b1111110101100000; // vC= -672 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100111; // iC=-1753 
// vC = 14'b1111110110111100; // vC= -580 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010001; // iC=-1775 
// vC = 14'b1111110110111100; // vC= -580 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001010; // iC=-1654 
// vC = 14'b1111110110001111; // vC= -625 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101000; // iC=-1688 
// vC = 14'b1111110011111110; // vC= -770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111000; // iC=-1800 
// vC = 14'b1111110100101001; // vC= -727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010001; // iC=-1583 
// vC = 14'b1111110101111000; // vC= -648 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011111; // iC=-1633 
// vC = 14'b1111110100001111; // vC= -753 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111111; // iC=-1601 
// vC = 14'b1111110111011100; // vC= -548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000000; // iC=-1792 
// vC = 14'b1111110111011100; // vC= -548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100010; // iC=-1694 
// vC = 14'b1111110010111010; // vC= -838 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111000; // iC=-1736 
// vC = 14'b1111110011001001; // vC= -823 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110001; // iC=-1551 
// vC = 14'b1111110101111100; // vC= -644 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111010; // iC=-1606 
// vC = 14'b1111110100111010; // vC= -710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100001; // iC=-1695 
// vC = 14'b1111110011101010; // vC= -790 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b1111110110101100; // vC= -596 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101110; // iC=-1746 
// vC = 14'b1111110100101001; // vC= -727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b1111110011000001; // vC= -831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b1111110011110000; // vC= -784 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011110; // iC=-1762 
// vC = 14'b1111110011001010; // vC= -822 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000100; // iC=-1660 
// vC = 14'b1111110011110111; // vC= -777 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001101; // iC=-1651 
// vC = 14'b1111110010111110; // vC= -834 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111101; // iC=-1795 
// vC = 14'b1111110010111011; // vC= -837 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110101; // iC=-1547 
// vC = 14'b1111110100101100; // vC= -724 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011000; // iC=-1512 
// vC = 14'b1111110101000101; // vC= -699 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110100; // iC=-1740 
// vC = 14'b1111110110001111; // vC= -625 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011000; // iC=-1640 
// vC = 14'b1111110100010100; // vC= -748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001001; // iC=-1783 
// vC = 14'b1111110010111000; // vC= -840 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100110; // iC=-1754 
// vC = 14'b1111110101000010; // vC= -702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100110; // iC=-1562 
// vC = 14'b1111110100100100; // vC= -732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100001; // iC=-1503 
// vC = 14'b1111110001001001; // vC= -951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011010; // iC=-1638 
// vC = 14'b1111110011100100; // vC= -796 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110011; // iC=-1741 
// vC = 14'b1111110010000001; // vC= -895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000011; // iC=-1533 
// vC = 14'b1111110100000101; // vC= -763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101111; // iC=-1553 
// vC = 14'b1111110010101101; // vC= -851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010111; // iC=-1705 
// vC = 14'b1111110010110010; // vC= -846 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001011; // iC=-1653 
// vC = 14'b1111110001011100; // vC= -932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010010; // iC=-1518 
// vC = 14'b1111110011101111; // vC= -785 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101000; // iC=-1560 
// vC = 14'b1111110100010001; // vC= -751 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100011; // iC=-1629 
// vC = 14'b1111110011001101; // vC= -819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b1111110100001111; // vC= -753 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111100; // iC=-1604 
// vC = 14'b1111101111011100; // vC=-1060 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111111; // iC=-1537 
// vC = 14'b1111110011101100; // vC= -788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010011; // iC=-1517 
// vC = 14'b1111110000011011; // vC= -997 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010000; // iC=-1712 
// vC = 14'b1111110000000110; // vC=-1018 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000010; // iC=-1470 
// vC = 14'b1111101111000001; // vC=-1087 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111010; // iC=-1734 
// vC = 14'b1111110001101000; // vC= -920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101110; // iC=-1426 
// vC = 14'b1111110011101011; // vC= -789 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110101; // iC=-1419 
// vC = 14'b1111110000100010; // vC= -990 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000111; // iC=-1529 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001100; // iC=-1652 
// vC = 14'b1111110000111100; // vC= -964 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101101; // iC=-1427 
// vC = 14'b1111101111110101; // vC=-1035 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101000; // iC=-1496 
// vC = 14'b1111101111111110; // vC=-1026 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011100; // iC=-1380 
// vC = 14'b1111110001011000; // vC= -936 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001010; // iC=-1462 
// vC = 14'b1111101111100101; // vC=-1051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011000; // iC=-1448 
// vC = 14'b1111110000010000; // vC=-1008 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010000; // iC=-1584 
// vC = 14'b1111110000011011; // vC= -997 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010110; // iC=-1386 
// vC = 14'b1111101111100111; // vC=-1049 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100011; // iC=-1437 
// vC = 14'b1111110000110101; // vC= -971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100111; // iC=-1561 
// vC = 14'b1111110001011111; // vC= -929 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001100; // iC=-1524 
// vC = 14'b1111110001111010; // vC= -902 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110111; // iC=-1673 
// vC = 14'b1111101111110010; // vC=-1038 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101101; // iC=-1363 
// vC = 14'b1111101101110101; // vC=-1163 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000011; // iC=-1405 
// vC = 14'b1111110000110010; // vC= -974 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000110; // iC=-1338 
// vC = 14'b1111101101101100; // vC=-1172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011010; // iC=-1574 
// vC = 14'b1111101101110110; // vC=-1162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011001; // iC=-1447 
// vC = 14'b1111101100111011; // vC=-1221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111111; // iC=-1473 
// vC = 14'b1111110000010111; // vC=-1001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011100; // iC=-1636 
// vC = 14'b1111101111101010; // vC=-1046 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011110; // iC=-1314 
// vC = 14'b1111101100111110; // vC=-1218 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000111; // iC=-1337 
// vC = 14'b1111110001100001; // vC= -927 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101001; // iC=-1431 
// vC = 14'b1111101110010000; // vC=-1136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001101; // iC=-1523 
// vC = 14'b1111110000010010; // vC=-1006 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010000; // iC=-1392 
// vC = 14'b1111101100110000; // vC=-1232 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001001; // iC=-1399 
// vC = 14'b1111101101111111; // vC=-1153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010100; // iC=-1324 
// vC = 14'b1111101101000111; // vC=-1209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010101; // iC=-1579 
// vC = 14'b1111101110111010; // vC=-1094 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010001; // iC=-1455 
// vC = 14'b1111101111000011; // vC=-1085 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000010; // iC=-1342 
// vC = 14'b1111101111100000; // vC=-1056 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001110; // iC=-1394 
// vC = 14'b1111101110110101; // vC=-1099 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010000; // iC=-1584 
// vC = 14'b1111101111000001; // vC=-1087 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101000; // iC=-1304 
// vC = 14'b1111101100001010; // vC=-1270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110101; // iC=-1483 
// vC = 14'b1111101110001111; // vC=-1137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000101; // iC=-1275 
// vC = 14'b1111110000001000; // vC=-1016 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110100; // iC=-1420 
// vC = 14'b1111101101101100; // vC=-1172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001010; // iC=-1270 
// vC = 14'b1111101110100100; // vC=-1116 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101110; // iC=-1362 
// vC = 14'b1111110000000000; // vC=-1024 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011010; // iC=-1446 
// vC = 14'b1111101011111111; // vC=-1281 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100011; // iC=-1501 
// vC = 14'b1111101101001011; // vC=-1205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001101; // iC=-1267 
// vC = 14'b1111101100100100; // vC=-1244 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100101; // iC=-1243 
// vC = 14'b1111101111000100; // vC=-1084 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111001; // iC=-1223 
// vC = 14'b1111101100011011; // vC=-1253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100101; // iC=-1243 
// vC = 14'b1111101111011001; // vC=-1063 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011100; // iC=-1380 
// vC = 14'b1111101101100011; // vC=-1181 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111101; // iC=-1475 
// vC = 14'b1111101110011001; // vC=-1127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101101; // iC=-1235 
// vC = 14'b1111101100001100; // vC=-1268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011110; // iC=-1250 
// vC = 14'b1111101110010111; // vC=-1129 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010110; // iC=-1258 
// vC = 14'b1111101010111111; // vC=-1345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010101; // iC=-1259 
// vC = 14'b1111101110011110; // vC=-1122 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011100; // iC=-1252 
// vC = 14'b1111101110010110; // vC=-1130 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000001; // iC=-1215 
// vC = 14'b1111101011101011; // vC=-1301 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001001; // iC=-1271 
// vC = 14'b1111101100110110; // vC=-1226 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111101; // iC=-1219 
// vC = 14'b1111101101101110; // vC=-1170 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001010; // iC=-1462 
// vC = 14'b1111101100111010; // vC=-1222 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100100; // iC=-1308 
// vC = 14'b1111101010000011; // vC=-1405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101101; // iC=-1363 
// vC = 14'b1111101101100101; // vC=-1179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101010; // iC=-1430 
// vC = 14'b1111101101100010; // vC=-1182 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011000; // iC=-1448 
// vC = 14'b1111101101110100; // vC=-1164 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111111; // iC=-1153 
// vC = 14'b1111101011111110; // vC=-1282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010110; // iC=-1258 
// vC = 14'b1111101101100011; // vC=-1181 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001000; // iC=-1400 
// vC = 14'b1111101100101010; // vC=-1238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000100; // iC=-1276 
// vC = 14'b1111101001111000; // vC=-1416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100110; // iC=-1178 
// vC = 14'b1111101001111110; // vC=-1410 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100100; // iC=-1372 
// vC = 14'b1111101101101111; // vC=-1169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100111; // iC=-1241 
// vC = 14'b1111101101101010; // vC=-1174 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110111; // iC=-1289 
// vC = 14'b1111101011010110; // vC=-1322 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010010; // iC=-1198 
// vC = 14'b1111101100001100; // vC=-1268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110100; // iC=-1164 
// vC = 14'b1111101010001111; // vC=-1393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001010; // iC=-1334 
// vC = 14'b1111101000010101; // vC=-1515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001001; // iC=-1143 
// vC = 14'b1111101010001000; // vC=-1400 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010000; // iC=-1200 
// vC = 14'b1111101001100101; // vC=-1435 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011110; // iC=-1122 
// vC = 14'b1111101100010001; // vC=-1263 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111011; // iC=-1221 
// vC = 14'b1111101000011110; // vC=-1506 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001100; // iC=-1076 
// vC = 14'b1111101001010100; // vC=-1452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011100; // iC=-1252 
// vC = 14'b1111101000000101; // vC=-1531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010001; // iC=-1199 
// vC = 14'b1111101010001000; // vC=-1400 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111111; // iC=-1345 
// vC = 14'b1111101100100011; // vC=-1245 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001010; // iC=-1078 
// vC = 14'b1111101100011010; // vC=-1254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101011; // iC=-1109 
// vC = 14'b1111101001101111; // vC=-1425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001111; // iC=-1073 
// vC = 14'b1111101100010110; // vC=-1258 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101010; // iC=-1174 
// vC = 14'b1111101000010100; // vC=-1516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100010; // iC=-1118 
// vC = 14'b1111101001110001; // vC=-1423 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011100; // iC=-1252 
// vC = 14'b1111101010110011; // vC=-1357 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000100; // iC=-1020 
// vC = 14'b1111101011000010; // vC=-1342 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011100; // iC=-1060 
// vC = 14'b1111101010100110; // vC=-1370 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010010; // iC=-1262 
// vC = 14'b1111101100000011; // vC=-1277 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011001; // iC=-1063 
// vC = 14'b1111101001110101; // vC=-1419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001011; // iC=-1269 
// vC = 14'b1111101011101111; // vC=-1297 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001100; // iC=-1076 
// vC = 14'b1111101011101001; // vC=-1303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011010; // iC= -998 
// vC = 14'b1111101000100101; // vC=-1499 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000010; // iC=-1214 
// vC = 14'b1111100111111111; // vC=-1537 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111000; // iC=-1160 
// vC = 14'b1111100111110001; // vC=-1551 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011101; // iC=-1123 
// vC = 14'b1111101010001000; // vC=-1400 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000001; // iC= -959 
// vC = 14'b1111101011001110; // vC=-1330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110011; // iC=-1229 
// vC = 14'b1111101000100111; // vC=-1497 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011100; // iC=-1252 
// vC = 14'b1111101000011111; // vC=-1505 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100001; // iC=-1119 
// vC = 14'b1111101010001010; // vC=-1398 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000001; // iC=-1151 
// vC = 14'b1111101001110001; // vC=-1423 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110100; // iC= -972 
// vC = 14'b1111100110010111; // vC=-1641 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010010; // iC=-1134 
// vC = 14'b1111101001100111; // vC=-1433 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011110; // iC= -994 
// vC = 14'b1111100111000010; // vC=-1598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111111; // iC=-1025 
// vC = 14'b1111100111010100; // vC=-1580 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001101; // iC=-1075 
// vC = 14'b1111100101110111; // vC=-1673 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000100; // iC= -892 
// vC = 14'b1111100111111110; // vC=-1538 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000101; // iC=-1083 
// vC = 14'b1111101010100110; // vC=-1370 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010001; // iC=-1071 
// vC = 14'b1111100111000010; // vC=-1598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100000; // iC=-1056 
// vC = 14'b1111100111110111; // vC=-1545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101100; // iC=-1044 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110110; // iC=-1034 
// vC = 14'b1111101001000110; // vC=-1466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010000; // iC=-1008 
// vC = 14'b1111100111111011; // vC=-1541 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100110; // iC=-1050 
// vC = 14'b1111100101101011; // vC=-1685 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011111; // iC=-1057 
// vC = 14'b1111101001010011; // vC=-1453 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000011; // iC=-1149 
// vC = 14'b1111100101101110; // vC=-1682 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010011; // iC= -941 
// vC = 14'b1111101000010100; // vC=-1516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011100; // iC= -996 
// vC = 14'b1111101010000101; // vC=-1403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110110; // iC= -970 
// vC = 14'b1111100111011001; // vC=-1575 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101110; // iC= -914 
// vC = 14'b1111100101111001; // vC=-1671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011000; // iC=-1000 
// vC = 14'b1111100111110000; // vC=-1552 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100001; // iC=-1119 
// vC = 14'b1111100101000100; // vC=-1724 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111010; // iC= -838 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000100; // iC= -892 
// vC = 14'b1111100111000110; // vC=-1594 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110001; // iC= -847 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101110; // iC=-1106 
// vC = 14'b1111101001100001; // vC=-1439 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001110; // iC=-1010 
// vC = 14'b1111101001100001; // vC=-1439 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010100; // iC= -812 
// vC = 14'b1111100100100101; // vC=-1755 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100101; // iC= -859 
// vC = 14'b1111100110011010; // vC=-1638 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101011; // iC= -853 
// vC = 14'b1111100111100010; // vC=-1566 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110101; // iC= -843 
// vC = 14'b1111101000000101; // vC=-1531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001001; // iC=-1015 
// vC = 14'b1111100101110001; // vC=-1679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111110; // iC= -770 
// vC = 14'b1111100101000011; // vC=-1725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111010; // iC= -838 
// vC = 14'b1111100101101010; // vC=-1686 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001100; // iC= -948 
// vC = 14'b1111100111010010; // vC=-1582 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111101; // iC= -835 
// vC = 14'b1111100100001010; // vC=-1782 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000001; // iC=-1023 
// vC = 14'b1111100110111101; // vC=-1603 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000111; // iC= -889 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110011; // iC= -973 
// vC = 14'b1111100110101110; // vC=-1618 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011111; // iC= -993 
// vC = 14'b1111100101110110; // vC=-1674 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111100; // iC= -708 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011011; // iC= -997 
// vC = 14'b1111100100001101; // vC=-1779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110101; // iC= -779 
// vC = 14'b1111100110110110; // vC=-1610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110100; // iC= -780 
// vC = 14'b1111100110110101; // vC=-1611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111100; // iC= -900 
// vC = 14'b1111100101010111; // vC=-1705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000101; // iC= -955 
// vC = 14'b1111100111001110; // vC=-1586 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101001; // iC= -791 
// vC = 14'b1111100111110110; // vC=-1546 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111001; // iC= -711 
// vC = 14'b1111100011011010; // vC=-1830 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110011; // iC= -717 
// vC = 14'b1111100111000010; // vC=-1598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011010; // iC= -806 
// vC = 14'b1111100100100100; // vC=-1756 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000011; // iC= -829 
// vC = 14'b1111100101000000; // vC=-1728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111011; // iC= -709 
// vC = 14'b1111100101001110; // vC=-1714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101110; // iC= -722 
// vC = 14'b1111100111001010; // vC=-1590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001001; // iC= -695 
// vC = 14'b1111100101001101; // vC=-1715 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011010; // iC= -806 
// vC = 14'b1111100100101100; // vC=-1748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011011; // iC= -805 
// vC = 14'b1111100110001001; // vC=-1655 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101111; // iC= -657 
// vC = 14'b1111100011110011; // vC=-1805 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011101; // iC= -803 
// vC = 14'b1111100011000100; // vC=-1852 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110000; // iC= -784 
// vC = 14'b1111100110111111; // vC=-1601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110001; // iC= -591 
// vC = 14'b1111100110000101; // vC=-1659 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111001; // iC= -711 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000110; // iC= -826 
// vC = 14'b1111100011101111; // vC=-1809 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101100; // iC= -724 
// vC = 14'b1111100100000110; // vC=-1786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111101; // iC= -643 
// vC = 14'b1111100100011111; // vC=-1761 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010001; // iC= -559 
// vC = 14'b1111100111000010; // vC=-1598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111000; // iC= -840 
// vC = 14'b1111100100111011; // vC=-1733 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011100; // iC= -676 
// vC = 14'b1111100100100001; // vC=-1759 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111000; // iC= -648 
// vC = 14'b1111100110010100; // vC=-1644 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110111; // iC= -713 
// vC = 14'b1111100010111101; // vC=-1859 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001000; // iC= -632 
// vC = 14'b1111100100001101; // vC=-1779 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110100; // iC= -652 
// vC = 14'b1111100101101100; // vC=-1684 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101001; // iC= -663 
// vC = 14'b1111100011110110; // vC=-1802 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001010; // iC= -822 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010111; // iC= -809 
// vC = 14'b1111100011111001; // vC=-1799 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100100; // iC= -796 
// vC = 14'b1111100011110101; // vC=-1803 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110010; // iC= -718 
// vC = 14'b1111100101010101; // vC=-1707 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110011; // iC= -653 
// vC = 14'b1111100101011100; // vC=-1700 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001001; // iC= -631 
// vC = 14'b1111100010000111; // vC=-1913 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110100; // iC= -716 
// vC = 14'b1111100101101000; // vC=-1688 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110111; // iC= -649 
// vC = 14'b1111100010011001; // vC=-1895 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000111; // iC= -569 
// vC = 14'b1111100110011100; // vC=-1636 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001000; // iC= -760 
// vC = 14'b1111100101011110; // vC=-1698 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101011; // iC= -597 
// vC = 14'b1111100011110000; // vC=-1808 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100101; // iC= -667 
// vC = 14'b1111100011100101; // vC=-1819 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011111; // iC= -737 
// vC = 14'b1111100101001000; // vC=-1720 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110110; // iC= -586 
// vC = 14'b1111100010011100; // vC=-1892 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000010; // iC= -702 
// vC = 14'b1111100010111011; // vC=-1861 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101000; // iC= -536 
// vC = 14'b1111100010011101; // vC=-1891 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110000; // iC= -464 
// vC = 14'b1111100010110100; // vC=-1868 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011110; // iC= -418 
// vC = 14'b1111100101011101; // vC=-1699 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000110; // iC= -442 
// vC = 14'b1111100100100001; // vC=-1759 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110101; // iC= -459 
// vC = 14'b1111100011110010; // vC=-1806 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011100; // iC= -548 
// vC = 14'b1111100010110011; // vC=-1869 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100011; // iC= -605 
// vC = 14'b1111100100000001; // vC=-1791 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000100; // iC= -316 
// vC = 14'b1111100110101001; // vC=-1623 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101111; // iC= -401 
// vC = 14'b1111100100011011; // vC=-1765 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010011; // iC= -493 
// vC = 14'b1111100101011100; // vC=-1700 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001110; // iC= -498 
// vC = 14'b1111100100100110; // vC=-1754 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101100; // iC= -468 
// vC = 14'b1111100100111111; // vC=-1729 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000100; // iC= -316 
// vC = 14'b1111100011001101; // vC=-1843 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010100; // iC= -492 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100101; // iC= -347 
// vC = 14'b1111100101111110; // vC=-1666 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011110101; // iC= -267 
// vC = 14'b1111100101010101; // vC=-1707 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011101; // iC= -291 
// vC = 14'b1111100010000101; // vC=-1915 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001101; // iC= -435 
// vC = 14'b1111100101001111; // vC=-1713 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001101; // iC= -371 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001000; // iC= -312 
// vC = 14'b1111100010011110; // vC=-1890 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010001; // iC= -431 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011100011; // iC= -285 
// vC = 14'b1111100100101001; // vC=-1751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010100; // iC= -172 
// vC = 14'b1111100100100110; // vC=-1754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101100; // iC= -212 
// vC = 14'b1111100101001110; // vC=-1714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001011; // iC= -181 
// vC = 14'b1111100011001000; // vC=-1848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101001; // iC= -279 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100101; // iC=  -91 
// vC = 14'b1111100100000110; // vC=-1786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111110010; // iC=  -14 
// vC = 14'b1111100001110010; // vC=-1934 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100001; // iC=  -95 
// vC = 14'b1111100001101011; // vC=-1941 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000001; // iC=  -63 
// vC = 14'b1111100110010010; // vC=-1646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001111; // iC=  -49 
// vC = 14'b1111100010100010; // vC=-1886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001011; // iC= -245 
// vC = 14'b1111100101101001; // vC=-1687 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010100; // iC=   20 
// vC = 14'b1111100011110000; // vC=-1808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001000; // iC=  -56 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010100; // iC=   20 
// vC = 14'b1111100011100000; // vC=-1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010101; // iC= -171 
// vC = 14'b1111100010000001; // vC=-1919 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101001; // iC=  -23 
// vC = 14'b1111100101010110; // vC=-1706 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110110011; // iC=  -77 
// vC = 14'b1111100011011011; // vC=-1829 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011100; // iC=   92 
// vC = 14'b1111100100100101; // vC=-1755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010001; // iC= -111 
// vC = 14'b1111100001010111; // vC=-1961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001111; // iC=   79 
// vC = 14'b1111100100110111; // vC=-1737 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000110010; // iC=   50 
// vC = 14'b1111100010101010; // vC=-1878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100010; // iC=   34 
// vC = 14'b1111100101000010; // vC=-1726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010011; // iC=  147 
// vC = 14'b1111100001010111; // vC=-1961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110110; // iC=  246 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011111; // iC=   31 
// vC = 14'b1111100011001111; // vC=-1841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011000; // iC=   88 
// vC = 14'b1111100100101111; // vC=-1745 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100101; // iC=  165 
// vC = 14'b1111100010000011; // vC=-1917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011110; // iC=  350 
// vC = 14'b1111100001100001; // vC=-1951 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110100; // iC=  180 
// vC = 14'b1111100100000111; // vC=-1785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110010; // iC=  178 
// vC = 14'b1111100011101101; // vC=-1811 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011000; // iC=  344 
// vC = 14'b1111100011110111; // vC=-1801 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111010; // iC=  250 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101001; // iC=  425 
// vC = 14'b1111100010111111; // vC=-1857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011010; // iC=  474 
// vC = 14'b1111100001101101; // vC=-1939 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010101; // iC=  533 
// vC = 14'b1111100010000011; // vC=-1917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001111; // iC=  399 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100100; // iC=  292 
// vC = 14'b1111100100000001; // vC=-1791 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100001; // iC=  545 
// vC = 14'b1111100011000111; // vC=-1849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101000; // iC=  360 
// vC = 14'b1111100011011010; // vC=-1830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100111; // iC=  551 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111110; // iC=  574 
// vC = 14'b1111100011101001; // vC=-1815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110011; // iC=  435 
// vC = 14'b1111100100011110; // vC=-1762 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100010; // iC=  610 
// vC = 14'b1111100011101011; // vC=-1813 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100001; // iC=  481 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101101; // iC=  749 
// vC = 14'b1111100010000110; // vC=-1914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101000; // iC=  680 
// vC = 14'b1111100101011100; // vC=-1700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101010; // iC=  746 
// vC = 14'b1111100101011111; // vC=-1697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100000; // iC=  800 
// vC = 14'b1111100101100001; // vC=-1695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011101; // iC=  669 
// vC = 14'b1111100011001001; // vC=-1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001000; // iC=  584 
// vC = 14'b1111100110000001; // vC=-1663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110111; // iC=  695 
// vC = 14'b1111100101100001; // vC=-1695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101001; // iC=  937 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110110; // iC=  886 
// vC = 14'b1111100101110001; // vC=-1679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101101; // iC=  685 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110001; // iC= 1009 
// vC = 14'b1111100010110100; // vC=-1868 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010111; // iC=  727 
// vC = 14'b1111100110001111; // vC=-1649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111000; // iC=  824 
// vC = 14'b1111100011010011; // vC=-1837 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000011; // iC=  899 
// vC = 14'b1111100011001001; // vC=-1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011001; // iC=  985 
// vC = 14'b1111100101101110; // vC=-1682 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101101; // iC= 1069 
// vC = 14'b1111100110010101; // vC=-1643 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110000; // iC= 1008 
// vC = 14'b1111100111100001; // vC=-1567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100001; // iC=  929 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011111; // iC=  927 
// vC = 14'b1111100100101001; // vC=-1751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001011; // iC= 1099 
// vC = 14'b1111100011011101; // vC=-1827 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110000; // iC= 1200 
// vC = 14'b1111100011100011; // vC=-1821 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001101; // iC= 1037 
// vC = 14'b1111100100000000; // vC=-1792 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111110; // iC=  958 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001111; // iC= 1231 
// vC = 14'b1111100110101110; // vC=-1618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000011; // iC= 1283 
// vC = 14'b1111100101101101; // vC=-1683 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001101; // iC= 1165 
// vC = 14'b1111100110111101; // vC=-1603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000110; // iC= 1158 
// vC = 14'b1111100100001001; // vC=-1783 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100100; // iC= 1188 
// vC = 14'b1111100110011011; // vC=-1637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001010; // iC= 1290 
// vC = 14'b1111100100001101; // vC=-1779 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111101; // iC= 1213 
// vC = 14'b1111100110100100; // vC=-1628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000001; // iC= 1089 
// vC = 14'b1111100101010001; // vC=-1711 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111101; // iC= 1277 
// vC = 14'b1111100111110111; // vC=-1545 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010101; // iC= 1173 
// vC = 14'b1111100100010111; // vC=-1769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000111; // iC= 1223 
// vC = 14'b1111100101110110; // vC=-1674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011100; // iC= 1308 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010011; // iC= 1363 
// vC = 14'b1111100101100000; // vC=-1696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100010; // iC= 1250 
// vC = 14'b1111101000100001; // vC=-1503 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100100; // iC= 1252 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001110; // iC= 1294 
// vC = 14'b1111101000000011; // vC=-1533 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001111; // iC= 1423 
// vC = 14'b1111100101110000; // vC=-1680 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111000; // iC= 1528 
// vC = 14'b1111101000111101; // vC=-1475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b1111100110000110; // vC=-1658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110100; // iC= 1524 
// vC = 14'b1111101000010101; // vC=-1515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001000; // iC= 1544 
// vC = 14'b1111101001000111; // vC=-1465 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101000; // iC= 1384 
// vC = 14'b1111100111000011; // vC=-1597 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110011; // iC= 1331 
// vC = 14'b1111101000110111; // vC=-1481 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101010; // iC= 1642 
// vC = 14'b1111100111001011; // vC=-1589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001110; // iC= 1550 
// vC = 14'b1111101001011111; // vC=-1441 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001101; // iC= 1421 
// vC = 14'b1111101000101111; // vC=-1489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010100; // iC= 1556 
// vC = 14'b1111100110010010; // vC=-1646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b1111101010011011; // vC=-1381 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101000; // iC= 1576 
// vC = 14'b1111100110100011; // vC=-1629 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010101; // iC= 1493 
// vC = 14'b1111101010110100; // vC=-1356 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100011; // iC= 1699 
// vC = 14'b1111100110111001; // vC=-1607 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111010; // iC= 1530 
// vC = 14'b1111101010111010; // vC=-1350 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010100; // iC= 1556 
// vC = 14'b1111101011000011; // vC=-1341 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011010; // iC= 1626 
// vC = 14'b1111101001001010; // vC=-1462 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001000; // iC= 1736 
// vC = 14'b1111101000011110; // vC=-1506 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010100; // iC= 1620 
// vC = 14'b1111101011011111; // vC=-1313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110001; // iC= 1649 
// vC = 14'b1111101000100110; // vC=-1498 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111100; // iC= 1660 
// vC = 14'b1111101001010011; // vC=-1453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010101; // iC= 1557 
// vC = 14'b1111101100000111; // vC=-1273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110111; // iC= 1655 
// vC = 14'b1111101010101011; // vC=-1365 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010110; // iC= 1622 
// vC = 14'b1111101010100000; // vC=-1376 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b1111101011111010; // vC=-1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111100; // iC= 1660 
// vC = 14'b1111101000001101; // vC=-1523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110101; // iC= 1781 
// vC = 14'b1111101010110110; // vC=-1354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111111; // iC= 1791 
// vC = 14'b1111101010100111; // vC=-1369 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000000; // iC= 1856 
// vC = 14'b1111101010101001; // vC=-1367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001110; // iC= 1806 
// vC = 14'b1111101010000101; // vC=-1403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001011; // iC= 1675 
// vC = 14'b1111101011001010; // vC=-1334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010101; // iC= 1685 
// vC = 14'b1111101101000110; // vC=-1210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000110; // iC= 1734 
// vC = 14'b1111101100001000; // vC=-1272 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000011; // iC= 1923 
// vC = 14'b1111101010101010; // vC=-1366 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111010; // iC= 1722 
// vC = 14'b1111101010011101; // vC=-1379 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110011; // iC= 1779 
// vC = 14'b1111101101100001; // vC=-1183 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000010; // iC= 1666 
// vC = 14'b1111101011000110; // vC=-1338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010001; // iC= 1681 
// vC = 14'b1111101010101010; // vC=-1366 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000001; // iC= 1729 
// vC = 14'b1111101011011011; // vC=-1317 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b1111101110010000; // vC=-1136 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100011; // iC= 1763 
// vC = 14'b1111101011101101; // vC=-1299 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111111; // iC= 1791 
// vC = 14'b1111101101000000; // vC=-1216 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100110; // iC= 1766 
// vC = 14'b1111101011110101; // vC=-1291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010001; // iC= 2001 
// vC = 14'b1111101100110100; // vC=-1228 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100010; // iC= 1762 
// vC = 14'b1111101010011100; // vC=-1380 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b1111101110111100; // vC=-1092 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100001; // iC= 2017 
// vC = 14'b1111101010100010; // vC=-1374 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110101; // iC= 1781 
// vC = 14'b1111101100110000; // vC=-1232 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111101010111100; // vC=-1348 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110111; // iC= 1911 
// vC = 14'b1111101111001111; // vC=-1073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011010; // iC= 1882 
// vC = 14'b1111101101110100; // vC=-1164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111010; // iC= 1914 
// vC = 14'b1111101101101100; // vC=-1172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b1111101110101101; // vC=-1107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011010; // iC= 2074 
// vC = 14'b1111101101001110; // vC=-1202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b1111101111000111; // vC=-1081 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111101011110110; // vC=-1290 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000010; // iC= 1922 
// vC = 14'b1111101100101100; // vC=-1236 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011000; // iC= 2072 
// vC = 14'b1111101111110010; // vC=-1038 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b1111110000001111; // vC=-1009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b1111101101110100; // vC=-1164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111011; // iC= 1915 
// vC = 14'b1111101100110110; // vC=-1226 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010001; // iC= 1809 
// vC = 14'b1111101110111101; // vC=-1091 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011110; // iC= 2078 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010100; // iC= 1876 
// vC = 14'b1111101101111110; // vC=-1154 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011111; // iC= 1823 
// vC = 14'b1111101111000110; // vC=-1082 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b1111110000101001; // vC= -983 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111110010000011; // vC= -893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111110000101100; // vC= -980 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b1111110010011101; // vC= -867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b1111101101111011; // vC=-1157 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100010; // iC= 2082 
// vC = 14'b1111110000101100; // vC= -980 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110001; // iC= 2097 
// vC = 14'b1111101111111101; // vC=-1027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000001; // iC= 1921 
// vC = 14'b1111101111100011; // vC=-1053 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001101; // iC= 1869 
// vC = 14'b1111110010000000; // vC= -896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b1111110000001110; // vC=-1010 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100101; // iC= 1893 
// vC = 14'b1111110001111101; // vC= -899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111101111011000; // vC=-1064 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b1111110011010100; // vC= -812 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100010; // iC= 2082 
// vC = 14'b1111110011110101; // vC= -779 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b1111101110111111; // vC=-1089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b1111101111110110; // vC=-1034 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110100; // iC= 2036 
// vC = 14'b1111101111100111; // vC=-1049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b1111110001011100; // vC= -932 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b1111101111101110; // vC=-1042 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111100; // iC= 1980 
// vC = 14'b1111110010100111; // vC= -857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101111; // iC= 1839 
// vC = 14'b1111110011100111; // vC= -793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b1111110001100110; // vC= -922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b1111110011110000; // vC= -784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111010; // iC= 2106 
// vC = 14'b1111110100001111; // vC= -753 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111110010000010; // vC= -894 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111110101010010; // vC= -686 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110110; // iC= 2038 
// vC = 14'b1111110000111011; // vC= -965 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001111; // iC= 1871 
// vC = 14'b1111110100100000; // vC= -736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101100; // iC= 2092 
// vC = 14'b1111110001101001; // vC= -919 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b1111110011011001; // vC= -807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000110; // iC= 2118 
// vC = 14'b1111110101111001; // vC= -647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111110; // iC= 1854 
// vC = 14'b1111110100111100; // vC= -708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b1111110010010100; // vC= -876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111110100101001; // vC= -727 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101110; // iC= 1838 
// vC = 14'b1111110101101101; // vC= -659 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b1111110011111010; // vC= -774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b1111110010100110; // vC= -858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111000; // iC= 1848 
// vC = 14'b1111110101101110; // vC= -658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011100; // iC= 1948 
// vC = 14'b1111110110110011; // vC= -589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111011; // iC= 1915 
// vC = 14'b1111110101001001; // vC= -695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000110; // iC= 2118 
// vC = 14'b1111110011101110; // vC= -786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b1111110011001101; // vC= -819 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101010; // iC= 2090 
// vC = 14'b1111110100011001; // vC= -743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b1111110101111111; // vC= -641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b1111110110011101; // vC= -611 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b1111110111100111; // vC= -537 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010011; // iC= 1875 
// vC = 14'b1111110111001100; // vC= -564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110110; // iC= 1910 
// vC = 14'b1111110111010001; // vC= -559 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100011; // iC= 2083 
// vC = 14'b1111110111101000; // vC= -536 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011100; // iC= 2076 
// vC = 14'b1111110111111110; // vC= -514 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111110111011101; // vC= -547 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010110; // iC= 2070 
// vC = 14'b1111110101101100; // vC= -660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111110; // iC= 2046 
// vC = 14'b1111110101111011; // vC= -645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101110; // iC= 1902 
// vC = 14'b1111111001001100; // vC= -436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101100; // iC= 2092 
// vC = 14'b1111111000010001; // vC= -495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b1111110110010100; // vC= -620 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101101; // iC= 2093 
// vC = 14'b1111110100111100; // vC= -708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101110; // iC= 2158 
// vC = 14'b1111110110101011; // vC= -597 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b1111110111011110; // vC= -546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b1111111000110000; // vC= -464 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b1111111010000100; // vC= -380 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011010; // iC= 1882 
// vC = 14'b1111111000111110; // vC= -450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000110; // iC= 2118 
// vC = 14'b1111111010010001; // vC= -367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000000; // iC= 2112 
// vC = 14'b1111111001010100; // vC= -428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100010; // iC= 2146 
// vC = 14'b1111110111010011; // vC= -557 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110101; // iC= 1845 
// vC = 14'b1111111010100111; // vC= -345 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111010; // iC= 1850 
// vC = 14'b1111111001000100; // vC= -444 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101100; // iC= 2092 
// vC = 14'b1111110110101000; // vC= -600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b1111111010011110; // vC= -354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100000; // iC= 2080 
// vC = 14'b1111111001110110; // vC= -394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b1111111011000110; // vC= -314 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101001; // iC= 2153 
// vC = 14'b1111111011011100; // vC= -292 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101011; // iC= 2155 
// vC = 14'b1111110111110100; // vC= -524 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010101; // iC= 2133 
// vC = 14'b1111111011100101; // vC= -283 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b1111111010001111; // vC= -369 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b1111111001001100; // vC= -436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b1111111011110011; // vC= -269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b1111111010010000; // vC= -368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b1111111010111111; // vC= -321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111111010100011; // vC= -349 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b1111111100101010; // vC= -214 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011111; // iC= 2143 
// vC = 14'b1111111101000010; // vC= -190 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100101; // iC= 1957 
// vC = 14'b1111111011110011; // vC= -269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b1111111011011011; // vC= -293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001101; // iC= 1997 
// vC = 14'b1111111011010110; // vC= -298 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b1111111001001101; // vC= -435 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b1111111100101110; // vC= -210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000001; // iC= 2049 
// vC = 14'b1111111001011010; // vC= -422 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b1111111010000010; // vC= -382 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100001; // iC= 2145 
// vC = 14'b1111111100110010; // vC= -206 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100111; // iC= 1831 
// vC = 14'b1111111101111101; // vC= -131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111111101101000; // vC= -152 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101010; // iC= 1898 
// vC = 14'b1111111011010110; // vC= -298 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101100; // iC= 2092 
// vC = 14'b1111111100000011; // vC= -253 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b1111111001110110; // vC= -394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b1111111011010110; // vC= -298 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b1111111100100000; // vC= -224 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100101; // iC= 1829 
// vC = 14'b1111111010101110; // vC= -338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b1111111011101101; // vC= -275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111101; // iC= 2045 
// vC = 14'b1111111101111010; // vC= -134 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001111; // iC= 1871 
// vC = 14'b1111111011100100; // vC= -284 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000101; // iC= 2117 
// vC = 14'b1111111011100111; // vC= -281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010101; // iC= 2133 
// vC = 14'b1111111101001101; // vC= -179 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b1111111011101101; // vC= -275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001110; // iC= 1870 
// vC = 14'b1111111101001101; // vC= -179 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010000; // iC= 2000 
// vC = 14'b1111111100101110; // vC= -210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b1111111111110011; // vC=  -13 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101101; // iC= 2093 
// vC = 14'b1111111111001000; // vC=  -56 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001000; // iC= 1992 
// vC = 14'b1111111100100111; // vC= -217 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110011; // iC= 2099 
// vC = 14'b1111111101011111; // vC= -161 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100110; // iC= 2022 
// vC = 14'b0000000000010111; // vC=   23 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100010; // iC= 2018 
// vC = 14'b1111111100100101; // vC= -219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011101; // iC= 1885 
// vC = 14'b1111111100100001; // vC= -223 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010101; // iC= 1813 
// vC = 14'b1111111110101010; // vC=  -86 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110001; // iC= 2097 
// vC = 14'b1111111110101001; // vC=  -87 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111111111000101; // vC=  -59 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001000; // iC= 2120 
// vC = 14'b1111111111111111; // vC=   -1 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111010; // iC= 1978 
// vC = 14'b0000000000011110; // vC=   30 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010010; // iC= 2066 
// vC = 14'b0000000001010100; // vC=   84 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111011; // iC= 1851 
// vC = 14'b0000000000100000; // vC=   32 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110111; // iC= 1911 
// vC = 14'b1111111111101010; // vC=  -22 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b0000000000101101; // vC=   45 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000101; // iC= 1861 
// vC = 14'b0000000001101011; // vC=  107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111011; // iC= 1851 
// vC = 14'b0000000001100100; // vC=  100 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b0000000001011111; // vC=   95 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011000; // iC= 1880 
// vC = 14'b0000000000100100; // vC=   36 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001110; // iC= 1934 
// vC = 14'b0000000000101110; // vC=   46 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100011; // iC= 1827 
// vC = 14'b0000000000000011; // vC=    3 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110101; // iC= 1909 
// vC = 14'b0000000001111011; // vC=  123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110000; // iC= 1840 
// vC = 14'b1111111111011101; // vC=  -35 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b0000000010111001; // vC=  185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b0000000010000011; // vC=  131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100101; // iC= 1957 
// vC = 14'b0000000010011000; // vC=  152 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110001; // iC= 2097 
// vC = 14'b0000000011010101; // vC=  213 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b1111111111100010; // vC=  -30 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001000; // iC= 1864 
// vC = 14'b0000000001110011; // vC=  115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b0000000001101010; // vC=  106 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010001; // iC= 2065 
// vC = 14'b0000000010110000; // vC=  176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b0000000001110010; // vC=  114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100100; // iC= 1828 
// vC = 14'b0000000100100011; // vC=  291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101001; // iC= 1769 
// vC = 14'b0000000000101111; // vC=   47 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110110; // iC= 1782 
// vC = 14'b0000000011011110; // vC=  222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b0000000011111000; // vC=  248 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110001; // iC= 1969 
// vC = 14'b0000000000100110; // vC=   38 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b0000000101001110; // vC=  334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110001; // iC= 1841 
// vC = 14'b0000000011001101; // vC=  205 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000010; // iC= 1858 
// vC = 14'b0000000101000100; // vC=  324 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100010; // iC= 1890 
// vC = 14'b0000000001110001; // vC=  113 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110110; // iC= 1782 
// vC = 14'b0000000100101100; // vC=  300 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b0000000101000010; // vC=  322 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100100; // iC= 1828 
// vC = 14'b0000000101011110; // vC=  350 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100111; // iC= 2023 
// vC = 14'b0000000001100100; // vC=  100 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b0000000100111100; // vC=  316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b0000000101101011; // vC=  363 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100101; // iC= 1765 
// vC = 14'b0000000100001111; // vC=  271 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011110; // iC= 1758 
// vC = 14'b0000000100101010; // vC=  298 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010011; // iC= 1747 
// vC = 14'b0000000101111110; // vC=  382 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b0000000011010110; // vC=  214 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100001; // iC= 1761 
// vC = 14'b0000000011010111; // vC=  215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b0000000101010111; // vC=  343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b0000000111001100; // vC=  460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101110; // iC= 1966 
// vC = 14'b0000000111000101; // vC=  453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b0000000100001000; // vC=  264 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001111; // iC= 1871 
// vC = 14'b0000000011111110; // vC=  254 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001011; // iC= 1995 
// vC = 14'b0000000110011111; // vC=  415 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b0000000101010011; // vC=  339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010010; // iC= 2002 
// vC = 14'b0000000100000000; // vC=  256 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100000; // iC= 1824 
// vC = 14'b0000001000001101; // vC=  525 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b0000000100000111; // vC=  263 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001001; // iC= 1993 
// vC = 14'b0000000100111100; // vC=  316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000000; // iC= 1856 
// vC = 14'b0000000110101111; // vC=  431 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b0000001000000110; // vC=  518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101001; // iC= 1705 
// vC = 14'b0000001000111110; // vC=  574 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000010; // iC= 1986 
// vC = 14'b0000001000110111; // vC=  567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110100; // iC= 1844 
// vC = 14'b0000000101001111; // vC=  335 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b0000000101100010; // vC=  354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001010; // iC= 1994 
// vC = 14'b0000000110011111; // vC=  415 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111010; // iC= 1722 
// vC = 14'b0000000100110100; // vC=  308 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000000; // iC= 1856 
// vC = 14'b0000000111111100; // vC=  508 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101001; // iC= 1833 
// vC = 14'b0000000101000011; // vC=  323 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100000; // iC= 1888 
// vC = 14'b0000000110110100; // vC=  436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101100; // iC= 1772 
// vC = 14'b0000000101001101; // vC=  333 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000001000001101; // vC=  525 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000000111011011; // vC=  475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110011; // iC= 1971 
// vC = 14'b0000001000010000; // vC=  528 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011011; // iC= 1755 
// vC = 14'b0000000111100001; // vC=  481 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000110; // iC= 1734 
// vC = 14'b0000001001010001; // vC=  593 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000011; // iC= 1859 
// vC = 14'b0000000110100101; // vC=  421 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110101; // iC= 1909 
// vC = 14'b0000001001010111; // vC=  599 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100100; // iC= 1764 
// vC = 14'b0000001001100001; // vC=  609 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100101; // iC= 1701 
// vC = 14'b0000000111100111; // vC=  487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101011; // iC= 1707 
// vC = 14'b0000000111010011; // vC=  467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b0000001011001010; // vC=  714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110000; // iC= 1840 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101110; // iC= 1902 
// vC = 14'b0000001000101000; // vC=  552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110101; // iC= 1845 
// vC = 14'b0000000111011010; // vC=  474 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100100; // iC= 1892 
// vC = 14'b0000001011010110; // vC=  726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011110; // iC= 1822 
// vC = 14'b0000000111000111; // vC=  455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010011; // iC= 1875 
// vC = 14'b0000001010010001; // vC=  657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001010; // iC= 1866 
// vC = 14'b0000001011011011; // vC=  731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111101; // iC= 1789 
// vC = 14'b0000001011011001; // vC=  729 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b0000001001001001; // vC=  585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101100; // iC= 1708 
// vC = 14'b0000001001000000; // vC=  576 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010001; // iC= 1617 
// vC = 14'b0000001011101001; // vC=  745 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b0000001100100111; // vC=  807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b0000001011110111; // vC=  759 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000111; // iC= 1799 
// vC = 14'b0000001100011011; // vC=  795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b0000001000010111; // vC=  535 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001010; // iC= 1738 
// vC = 14'b0000001001001001; // vC=  585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110111; // iC= 1655 
// vC = 14'b0000001001110011; // vC=  627 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101010; // iC= 1770 
// vC = 14'b0000001101100010; // vC=  866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001010; // iC= 1866 
// vC = 14'b0000001010000100; // vC=  644 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111000; // iC= 1656 
// vC = 14'b0000001101100000; // vC=  864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000010; // iC= 1602 
// vC = 14'b0000001001111101; // vC=  637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010111; // iC= 1623 
// vC = 14'b0000001000111011; // vC=  571 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110001; // iC= 1777 
// vC = 14'b0000001100110100; // vC=  820 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100001; // iC= 1697 
// vC = 14'b0000001100010000; // vC=  784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101101; // iC= 1837 
// vC = 14'b0000001101000101; // vC=  837 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100000; // iC= 1760 
// vC = 14'b0000001100000101; // vC=  773 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101110; // iC= 1582 
// vC = 14'b0000001010001000; // vC=  648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011000; // iC= 1624 
// vC = 14'b0000001010010010; // vC=  658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000000; // iC= 1600 
// vC = 14'b0000001010110010; // vC=  690 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101110; // iC= 1774 
// vC = 14'b0000001010111110; // vC=  702 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101111; // iC= 1711 
// vC = 14'b0000001011010001; // vC=  721 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100000; // iC= 1824 
// vC = 14'b0000001010101110; // vC=  686 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111101; // iC= 1725 
// vC = 14'b0000001101110101; // vC=  885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000101; // iC= 1797 
// vC = 14'b0000001110100101; // vC=  933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011110; // iC= 1566 
// vC = 14'b0000001011101111; // vC=  751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111110; // iC= 1662 
// vC = 14'b0000001010111011; // vC=  699 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010110; // iC= 1622 
// vC = 14'b0000001011001111; // vC=  719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111001; // iC= 1529 
// vC = 14'b0000001111001001; // vC=  969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000010; // iC= 1730 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001010; // iC= 1738 
// vC = 14'b0000001101011001; // vC=  857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010111; // iC= 1559 
// vC = 14'b0000001110001000; // vC=  904 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111101; // iC= 1597 
// vC = 14'b0000001111001001; // vC=  969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100101; // iC= 1509 
// vC = 14'b0000001111000010; // vC=  962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101100; // iC= 1772 
// vC = 14'b0000010000010110; // vC= 1046 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101100; // iC= 1772 
// vC = 14'b0000001101000101; // vC=  837 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101001; // iC= 1641 
// vC = 14'b0000001110111010; // vC=  954 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001011; // iC= 1803 
// vC = 14'b0000001111100001; // vC=  993 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b0000010000001110; // vC= 1038 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000000; // iC= 1792 
// vC = 14'b0000001111000101; // vC=  965 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110010; // iC= 1714 
// vC = 14'b0000001101100000; // vC=  864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110010; // iC= 1714 
// vC = 14'b0000001101001111; // vC=  847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000000; // iC= 1664 
// vC = 14'b0000001111110010; // vC= 1010 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000000; // iC= 1728 
// vC = 14'b0000010000011011; // vC= 1051 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000101; // iC= 1605 
// vC = 14'b0000010000111001; // vC= 1081 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100010; // iC= 1570 
// vC = 14'b0000001111111100; // vC= 1020 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101001; // iC= 1577 
// vC = 14'b0000001100111101; // vC=  829 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100001; // iC= 1761 
// vC = 14'b0000001111110011; // vC= 1011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010100; // iC= 1556 
// vC = 14'b0000010001011110; // vC= 1118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010000; // iC= 1616 
// vC = 14'b0000010001011000; // vC= 1112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011001; // iC= 1625 
// vC = 14'b0000001110011001; // vC=  921 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000101; // iC= 1477 
// vC = 14'b0000010000001110; // vC= 1038 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111001; // iC= 1721 
// vC = 14'b0000010000100010; // vC= 1058 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001111; // iC= 1679 
// vC = 14'b0000001110110101; // vC=  949 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001111; // iC= 1743 
// vC = 14'b0000001110111100; // vC=  956 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110000; // iC= 1584 
// vC = 14'b0000010000100101; // vC= 1061 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000110; // iC= 1734 
// vC = 14'b0000001110101010; // vC=  938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000001; // iC= 1729 
// vC = 14'b0000001110101111; // vC=  943 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011101; // iC= 1693 
// vC = 14'b0000010000100001; // vC= 1057 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101011; // iC= 1451 
// vC = 14'b0000010000111101; // vC= 1085 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001011; // iC= 1419 
// vC = 14'b0000010001000110; // vC= 1094 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011001; // iC= 1433 
// vC = 14'b0000001110001100; // vC=  908 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011000; // iC= 1688 
// vC = 14'b0000001111110000; // vC= 1008 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100101; // iC= 1637 
// vC = 14'b0000001111100000; // vC=  992 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100101; // iC= 1701 
// vC = 14'b0000001111100011; // vC=  995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110001; // iC= 1585 
// vC = 14'b0000001111000001; // vC=  961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010110; // iC= 1558 
// vC = 14'b0000010001110101; // vC= 1141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011000; // iC= 1624 
// vC = 14'b0000001111110101; // vC= 1013 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101011; // iC= 1579 
// vC = 14'b0000001111100100; // vC=  996 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111101; // iC= 1533 
// vC = 14'b0000010001101001; // vC= 1129 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010010; // iC= 1490 
// vC = 14'b0000010011101100; // vC= 1260 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101001; // iC= 1577 
// vC = 14'b0000010001111011; // vC= 1147 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010011; // iC= 1619 
// vC = 14'b0000010010000100; // vC= 1156 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010001; // iC= 1553 
// vC = 14'b0000001111101111; // vC= 1007 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100101; // iC= 1381 
// vC = 14'b0000010011101001; // vC= 1257 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100110; // iC= 1446 
// vC = 14'b0000001111110100; // vC= 1012 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101110; // iC= 1518 
// vC = 14'b0000010000001011; // vC= 1035 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101000; // iC= 1320 
// vC = 14'b0000010011011010; // vC= 1242 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010000; // iC= 1360 
// vC = 14'b0000010001000000; // vC= 1088 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100101; // iC= 1381 
// vC = 14'b0000010010100101; // vC= 1189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101011; // iC= 1515 
// vC = 14'b0000010010011000; // vC= 1176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101011; // iC= 1387 
// vC = 14'b0000010011101101; // vC= 1261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010110; // iC= 1366 
// vC = 14'b0000010000011001; // vC= 1049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110000; // iC= 1328 
// vC = 14'b0000010001100001; // vC= 1121 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001111; // iC= 1487 
// vC = 14'b0000010001111010; // vC= 1146 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000010; // iC= 1346 
// vC = 14'b0000010011011111; // vC= 1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111111; // iC= 1343 
// vC = 14'b0000010100101111; // vC= 1327 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100001; // iC= 1505 
// vC = 14'b0000010011101001; // vC= 1257 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000010; // iC= 1282 
// vC = 14'b0000010101001111; // vC= 1359 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001000; // iC= 1416 
// vC = 14'b0000010010001100; // vC= 1164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101110; // iC= 1518 
// vC = 14'b0000010010001011; // vC= 1163 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000011; // iC= 1475 
// vC = 14'b0000010010111000; // vC= 1208 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011000; // iC= 1496 
// vC = 14'b0000010011010001; // vC= 1233 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100110; // iC= 1446 
// vC = 14'b0000010100000111; // vC= 1287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111010; // iC= 1274 
// vC = 14'b0000010011110010; // vC= 1266 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101101; // iC= 1325 
// vC = 14'b0000010011111011; // vC= 1275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001011; // iC= 1419 
// vC = 14'b0000010101111010; // vC= 1402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101101; // iC= 1261 
// vC = 14'b0000010100100001; // vC= 1313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101000; // iC= 1448 
// vC = 14'b0000010100100101; // vC= 1317 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111011; // iC= 1403 
// vC = 14'b0000010101111010; // vC= 1402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111111; // iC= 1215 
// vC = 14'b0000010011001101; // vC= 1229 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100100; // iC= 1316 
// vC = 14'b0000010010110011; // vC= 1203 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111001; // iC= 1465 
// vC = 14'b0000010010111101; // vC= 1213 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111100; // iC= 1340 
// vC = 14'b0000010110101111; // vC= 1455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110110; // iC= 1270 
// vC = 14'b0000010100000101; // vC= 1285 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101100; // iC= 1260 
// vC = 14'b0000010111000011; // vC= 1475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111001; // iC= 1209 
// vC = 14'b0000010110011011; // vC= 1435 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111101; // iC= 1213 
// vC = 14'b0000010111000010; // vC= 1474 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111010; // iC= 1274 
// vC = 14'b0000010110010110; // vC= 1430 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010010; // iC= 1234 
// vC = 14'b0000010101000101; // vC= 1349 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101111; // iC= 1327 
// vC = 14'b0000010110110000; // vC= 1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110111; // iC= 1335 
// vC = 14'b0000010100000000; // vC= 1280 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010100; // iC= 1428 
// vC = 14'b0000010100110011; // vC= 1331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101001; // iC= 1257 
// vC = 14'b0000010011001011; // vC= 1227 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111100; // iC= 1404 
// vC = 14'b0000010100110001; // vC= 1329 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010110; // iC= 1366 
// vC = 14'b0000010101000010; // vC= 1346 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110001; // iC= 1393 
// vC = 14'b0000010011101111; // vC= 1263 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101111; // iC= 1327 
// vC = 14'b0000010100000011; // vC= 1283 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101101; // iC= 1389 
// vC = 14'b0000010011011100; // vC= 1244 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010001; // iC= 1297 
// vC = 14'b0000011000011100; // vC= 1564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011100; // iC= 1372 
// vC = 14'b0000010101110111; // vC= 1399 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110111; // iC= 1143 
// vC = 14'b0000010111011100; // vC= 1500 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101111; // iC= 1199 
// vC = 14'b0000010100111010; // vC= 1338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000000; // iC= 1408 
// vC = 14'b0000010100001111; // vC= 1295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000010; // iC= 1154 
// vC = 14'b0000010100001000; // vC= 1288 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100110; // iC= 1382 
// vC = 14'b0000011000000110; // vC= 1542 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000011; // iC= 1091 
// vC = 14'b0000010100111011; // vC= 1339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101000; // iC= 1320 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101100; // iC= 1260 
// vC = 14'b0000010111011101; // vC= 1501 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010100; // iC= 1364 
// vC = 14'b0000011000010100; // vC= 1556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101010; // iC= 1258 
// vC = 14'b0000011000100110; // vC= 1574 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011001; // iC= 1305 
// vC = 14'b0000010110000100; // vC= 1412 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111111; // iC= 1087 
// vC = 14'b0000010111100111; // vC= 1511 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101111; // iC= 1327 
// vC = 14'b0000010111011110; // vC= 1502 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011011; // iC= 1307 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001111; // iC= 1103 
// vC = 14'b0000011000011101; // vC= 1565 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101001; // iC= 1257 
// vC = 14'b0000011001110111; // vC= 1655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001011; // iC= 1163 
// vC = 14'b0000010111010101; // vC= 1493 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111111; // iC= 1023 
// vC = 14'b0000010110001111; // vC= 1423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010010; // iC= 1234 
// vC = 14'b0000010111000001; // vC= 1473 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001011; // iC= 1163 
// vC = 14'b0000010110001110; // vC= 1422 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101000; // iC= 1064 
// vC = 14'b0000011010010011; // vC= 1683 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111110; // iC= 1150 
// vC = 14'b0000010101011110; // vC= 1374 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001001; // iC= 1225 
// vC = 14'b0000010101110010; // vC= 1394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001011; // iC= 1035 
// vC = 14'b0000011000000000; // vC= 1536 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100001; // iC= 1057 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010001; // iC= 1041 
// vC = 14'b0000010110001111; // vC= 1423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010101; // iC= 1045 
// vC = 14'b0000010111100110; // vC= 1510 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011111; // iC= 1055 
// vC = 14'b0000010101111011; // vC= 1403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110100; // iC= 1204 
// vC = 14'b0000011000101110; // vC= 1582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111101; // iC=  957 
// vC = 14'b0000011001101110; // vC= 1646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011011; // iC= 1051 
// vC = 14'b0000010110111110; // vC= 1470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011110; // iC= 1246 
// vC = 14'b0000011000111111; // vC= 1599 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010001; // iC=  977 
// vC = 14'b0000010110011001; // vC= 1433 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110100; // iC= 1076 
// vC = 14'b0000011001000001; // vC= 1601 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110101; // iC= 1013 
// vC = 14'b0000011000101101; // vC= 1581 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000000; // iC= 1152 
// vC = 14'b0000010110110100; // vC= 1460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100010; // iC= 1058 
// vC = 14'b0000011001110010; // vC= 1650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000101; // iC= 1029 
// vC = 14'b0000011001100101; // vC= 1637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111101; // iC= 1213 
// vC = 14'b0000010111100001; // vC= 1505 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001110; // iC= 1102 
// vC = 14'b0000011000000001; // vC= 1537 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100010; // iC= 1058 
// vC = 14'b0000011001001000; // vC= 1608 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001001; // iC=  905 
// vC = 14'b0000011011000110; // vC= 1734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110110; // iC= 1078 
// vC = 14'b0000011001100011; // vC= 1635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100101; // iC= 1125 
// vC = 14'b0000010111011000; // vC= 1496 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110101; // iC=  885 
// vC = 14'b0000011001011111; // vC= 1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100111; // iC= 1063 
// vC = 14'b0000010111101000; // vC= 1512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111100; // iC= 1020 
// vC = 14'b0000011010010000; // vC= 1680 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111111; // iC=  959 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010000; // iC=  912 
// vC = 14'b0000011000110101; // vC= 1589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100110; // iC=  998 
// vC = 14'b0000011100010000; // vC= 1808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000111; // iC= 1159 
// vC = 14'b0000011010101100; // vC= 1708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001011; // iC= 1099 
// vC = 14'b0000011011011011; // vC= 1755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101111; // iC=  943 
// vC = 14'b0000011010101000; // vC= 1704 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011011; // iC=  859 
// vC = 14'b0000011000100010; // vC= 1570 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111101; // iC=  957 
// vC = 14'b0000011011101001; // vC= 1769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001000; // iC= 1032 
// vC = 14'b0000011011101100; // vC= 1772 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110000; // iC= 1072 
// vC = 14'b0000011011111110; // vC= 1790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000100; // iC=  836 
// vC = 14'b0000011010011111; // vC= 1695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010100; // iC=  980 
// vC = 14'b0000011011111101; // vC= 1789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000001; // iC= 1025 
// vC = 14'b0000011010011001; // vC= 1689 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000110; // iC=  838 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101000; // iC= 1064 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100000; // iC= 1056 
// vC = 14'b0000011001101110; // vC= 1646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011101; // iC=  925 
// vC = 14'b0000011100011010; // vC= 1818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001101; // iC=  781 
// vC = 14'b0000011010101010; // vC= 1706 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101000; // iC=  808 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010001; // iC=  913 
// vC = 14'b0000011011101011; // vC= 1771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110110; // iC=  886 
// vC = 14'b0000011100100011; // vC= 1827 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100111; // iC=  743 
// vC = 14'b0000011000011011; // vC= 1563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000111; // iC=  775 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110110; // iC=  950 
// vC = 14'b0000011011010111; // vC= 1751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010011; // iC=  723 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001011; // iC=  843 
// vC = 14'b0000011000110100; // vC= 1588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101010; // iC=  938 
// vC = 14'b0000011010111100; // vC= 1724 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011000; // iC=  920 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000001; // iC=  961 
// vC = 14'b0000011001010101; // vC= 1621 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110011; // iC=  819 
// vC = 14'b0000011001110000; // vC= 1648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001001; // iC=  905 
// vC = 14'b0000011010110001; // vC= 1713 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010101; // iC=  789 
// vC = 14'b0000011001011111; // vC= 1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001100; // iC=  716 
// vC = 14'b0000011100110100; // vC= 1844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000101; // iC=  837 
// vC = 14'b0000011011001011; // vC= 1739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101000; // iC=  680 
// vC = 14'b0000011100010110; // vC= 1814 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111101; // iC=  765 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100110; // iC=  870 
// vC = 14'b0000011010000001; // vC= 1665 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111001; // iC=  697 
// vC = 14'b0000011101110011; // vC= 1907 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011100; // iC=  860 
// vC = 14'b0000011101100011; // vC= 1891 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010110; // iC=  790 
// vC = 14'b0000011110001111; // vC= 1935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110100; // iC=  756 
// vC = 14'b0000011011001100; // vC= 1740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101000; // iC=  808 
// vC = 14'b0000011001101010; // vC= 1642 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110101; // iC=  821 
// vC = 14'b0000011100001101; // vC= 1805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111110; // iC=  702 
// vC = 14'b0000011011000101; // vC= 1733 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110010; // iC=  690 
// vC = 14'b0000011101011111; // vC= 1887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011011; // iC=  795 
// vC = 14'b0000011100011100; // vC= 1820 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000111; // iC=  711 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011110; // iC=  670 
// vC = 14'b0000011100100111; // vC= 1831 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111100; // iC=  636 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100111; // iC=  871 
// vC = 14'b0000011010100101; // vC= 1701 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100000; // iC=  736 
// vC = 14'b0000011110101010; // vC= 1962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110110; // iC=  694 
// vC = 14'b0000011110011001; // vC= 1945 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111001; // iC=  633 
// vC = 14'b0000011011100001; // vC= 1761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000101; // iC=  581 
// vC = 14'b0000011001111110; // vC= 1662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011110; // iC=  798 
// vC = 14'b0000011110110010; // vC= 1970 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110000; // iC=  624 
// vC = 14'b0000011110111100; // vC= 1980 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000100; // iC=  580 
// vC = 14'b0000011011100100; // vC= 1764 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011001; // iC=  537 
// vC = 14'b0000011100011001; // vC= 1817 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011111; // iC=  543 
// vC = 14'b0000011011101001; // vC= 1769 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000000; // iC=  576 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001100; // iC=  524 
// vC = 14'b0000011110011000; // vC= 1944 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001000; // iC=  776 
// vC = 14'b0000011101100010; // vC= 1890 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110110; // iC=  630 
// vC = 14'b0000011010010101; // vC= 1685 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100000; // iC=  736 
// vC = 14'b0000011110011101; // vC= 1949 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000000; // iC=  640 
// vC = 14'b0000011101000111; // vC= 1863 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100001; // iC=  737 
// vC = 14'b0000011101100011; // vC= 1891 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011000; // iC=  472 
// vC = 14'b0000011100111100; // vC= 1852 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110000; // iC=  688 
// vC = 14'b0000011110001110; // vC= 1934 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110011; // iC=  563 
// vC = 14'b0000011011010000; // vC= 1744 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001010; // iC=  458 
// vC = 14'b0000011111010101; // vC= 2005 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111010; // iC=  698 
// vC = 14'b0000011100100110; // vC= 1830 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000001; // iC=  449 
// vC = 14'b0000011100001100; // vC= 1804 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010000; // iC=  720 
// vC = 14'b0000011111010001; // vC= 2001 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100100; // iC=  612 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100000; // iC=  480 
// vC = 14'b0000011110110000; // vC= 1968 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001110; // iC=  654 
// vC = 14'b0000011111001100; // vC= 1996 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111110; // iC=  574 
// vC = 14'b0000011101001110; // vC= 1870 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100101; // iC=  677 
// vC = 14'b0000011111101101; // vC= 2029 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110110; // iC=  374 
// vC = 14'b0000011100111010; // vC= 1850 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000011; // iC=  643 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011101; // iC=  605 
// vC = 14'b0000011101000000; // vC= 1856 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010000; // iC=  400 
// vC = 14'b0000011011011110; // vC= 1758 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111011; // iC=  379 
// vC = 14'b0000011100011100; // vC= 1820 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000100; // iC=  580 
// vC = 14'b0000011110101010; // vC= 1962 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111101; // iC=  445 
// vC = 14'b0000011011001101; // vC= 1741 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111010; // iC=  506 
// vC = 14'b0000100000000010; // vC= 2050 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101110; // iC=  366 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111110; // iC=  254 
// vC = 14'b0000011111000011; // vC= 1987 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101110; // iC=  494 
// vC = 14'b0000011100101101; // vC= 1837 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000110; // iC=  198 
// vC = 14'b0000011111010111; // vC= 2007 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010111; // iC=  471 
// vC = 14'b0000011111111011; // vC= 2043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101011; // iC=  363 
// vC = 14'b0000011111010011; // vC= 2003 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010000; // iC=  464 
// vC = 14'b0000011111000110; // vC= 1990 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010110; // iC=  278 
// vC = 14'b0000011111000000; // vC= 1984 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000111; // iC=  327 
// vC = 14'b0000011101100010; // vC= 1890 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001110; // iC=  142 
// vC = 14'b0000100000000101; // vC= 2053 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101100; // iC=  236 
// vC = 14'b0000011011110101; // vC= 1781 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100111; // iC=  103 
// vC = 14'b0000011101000101; // vC= 1861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110010; // iC=  306 
// vC = 14'b0000011111111101; // vC= 2045 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011100; // iC=  348 
// vC = 14'b0000011101110001; // vC= 1905 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100000; // iC=  160 
// vC = 14'b0000011111100110; // vC= 2022 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100111; // iC=  167 
// vC = 14'b0000011011010101; // vC= 1749 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110100; // iC=  308 
// vC = 14'b0000011100001000; // vC= 1800 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010000; // iC=  144 
// vC = 14'b0000011100001001; // vC= 1801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011111; // iC=  287 
// vC = 14'b0000011100101110; // vC= 1838 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010000; // iC=   16 
// vC = 14'b0000011111000011; // vC= 1987 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011001; // iC=   25 
// vC = 14'b0000011101110000; // vC= 1904 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111011110; // iC=  -34 
// vC = 14'b0000011110100111; // vC= 1959 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001011; // iC=   75 
// vC = 14'b0000011011111110; // vC= 1790 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001011; // iC=   75 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001001; // iC=   73 
// vC = 14'b0000011111010101; // vC= 2005 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010110; // iC=   22 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000101; // iC=  -59 
// vC = 14'b0000100000000100; // vC= 2052 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000001; // iC= -191 
// vC = 14'b0000100000010010; // vC= 2066 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001010; // iC= -118 
// vC = 14'b0000011100110100; // vC= 1844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010100; // iC= -108 
// vC = 14'b0000011100001011; // vC= 1803 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101011001; // iC= -167 
// vC = 14'b0000011110011010; // vC= 1946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000011; // iC=    3 
// vC = 14'b0000011110011010; // vC= 1946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110110111; // iC=  -73 
// vC = 14'b0000011110111101; // vC= 1981 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000100; // iC= -252 
// vC = 14'b0000011101111101; // vC= 1917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010001; // iC= -367 
// vC = 14'b0000011111011100; // vC= 2012 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000010; // iC= -254 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001100; // iC= -308 
// vC = 14'b0000011101111000; // vC= 1912 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001111; // iC= -433 
// vC = 14'b0000011011001101; // vC= 1741 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001100; // iC= -244 
// vC = 14'b0000011110101011; // vC= 1963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000111; // iC= -313 
// vC = 14'b0000011111010111; // vC= 2007 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101000; // iC= -216 
// vC = 14'b0000011011100000; // vC= 1760 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011100100; // iC= -284 
// vC = 14'b0000011011111101; // vC= 1789 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001110; // iC= -370 
// vC = 14'b0000011100110001; // vC= 1841 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000000001; // iC= -511 
// vC = 14'b0000011110101111; // vC= 1967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011111; // iC= -289 
// vC = 14'b0000011011111011; // vC= 1787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100111; // iC= -409 
// vC = 14'b0000011100000110; // vC= 1798 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001100; // iC= -628 
// vC = 14'b0000011111010000; // vC= 2000 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010100; // iC= -492 
// vC = 14'b0000011101010101; // vC= 1877 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101011; // iC= -469 
// vC = 14'b0000011101111010; // vC= 1914 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001110; // iC= -498 
// vC = 14'b0000011101010100; // vC= 1876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000110; // iC= -698 
// vC = 14'b0000011110001010; // vC= 1930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000111; // iC= -633 
// vC = 14'b0000011011100011; // vC= 1763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101110; // iC= -722 
// vC = 14'b0000011101001100; // vC= 1868 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111011; // iC= -645 
// vC = 14'b0000011111000111; // vC= 1991 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010110; // iC= -554 
// vC = 14'b0000011011000110; // vC= 1734 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110010; // iC= -782 
// vC = 14'b0000011010101101; // vC= 1709 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010001; // iC= -559 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000000; // iC= -768 
// vC = 14'b0000011100010011; // vC= 1811 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101111; // iC= -785 
// vC = 14'b0000011010100111; // vC= 1703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000000; // iC= -832 
// vC = 14'b0000011011101110; // vC= 1774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000001; // iC= -959 
// vC = 14'b0000011011001100; // vC= 1740 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100000; // iC= -928 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010011; // iC= -813 
// vC = 14'b0000011100110000; // vC= 1840 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011011; // iC= -741 
// vC = 14'b0000011100100001; // vC= 1825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010010; // iC= -878 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000111; // iC= -889 
// vC = 14'b0000011010110000; // vC= 1712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101011; // iC=-1045 
// vC = 14'b0000011100011101; // vC= 1821 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111101; // iC=-1091 
// vC = 14'b0000011100100010; // vC= 1826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111111; // iC=-1025 
// vC = 14'b0000011011101110; // vC= 1774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100100; // iC=-1052 
// vC = 14'b0000011101010010; // vC= 1874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110100; // iC= -972 
// vC = 14'b0000011010011011; // vC= 1691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111111; // iC= -897 
// vC = 14'b0000011101100001; // vC= 1889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011000; // iC=-1064 
// vC = 14'b0000011101110111; // vC= 1911 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011100; // iC=-1124 
// vC = 14'b0000011101001010; // vC= 1866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010010; // iC=-1134 
// vC = 14'b0000011001001101; // vC= 1613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000101; // iC=-1211 
// vC = 14'b0000011010010001; // vC= 1681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000111; // iC=-1209 
// vC = 14'b0000011100110011; // vC= 1843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000010; // iC=-1086 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100011; // iC=-1181 
// vC = 14'b0000011010100010; // vC= 1698 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110110; // iC=-1098 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001011; // iC=-1205 
// vC = 14'b0000011000111101; // vC= 1597 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010001; // iC=-1263 
// vC = 14'b0000011100000100; // vC= 1796 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101111; // iC=-1297 
// vC = 14'b0000011101011101; // vC= 1885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111110; // iC=-1282 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111000; // iC=-1352 
// vC = 14'b0000011100101001; // vC= 1833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001111; // iC=-1265 
// vC = 14'b0000011100001011; // vC= 1803 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101110; // iC=-1234 
// vC = 14'b0000011001001010; // vC= 1610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011010; // iC=-1190 
// vC = 14'b0000011100010010; // vC= 1810 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011111; // iC=-1377 
// vC = 14'b0000011010010000; // vC= 1680 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010011; // iC=-1325 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111010; // iC=-1286 
// vC = 14'b0000011011101010; // vC= 1770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100001; // iC=-1375 
// vC = 14'b0000011010000011; // vC= 1667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011110; // iC=-1570 
// vC = 14'b0000011011110010; // vC= 1778 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101001; // iC=-1559 
// vC = 14'b0000010111101001; // vC= 1513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110100; // iC=-1420 
// vC = 14'b0000011010100110; // vC= 1702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110100; // iC=-1612 
// vC = 14'b0000010111101000; // vC= 1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111101; // iC=-1539 
// vC = 14'b0000011000100011; // vC= 1571 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110001; // iC=-1551 
// vC = 14'b0000011010100101; // vC= 1701 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011111; // iC=-1377 
// vC = 14'b0000010111101001; // vC= 1513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011011; // iC=-1637 
// vC = 14'b0000010110111010; // vC= 1466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100000; // iC=-1568 
// vC = 14'b0000011001001011; // vC= 1611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011000; // iC=-1640 
// vC = 14'b0000011001010000; // vC= 1616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000011; // iC=-1533 
// vC = 14'b0000011000100001; // vC= 1569 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100001; // iC=-1503 
// vC = 14'b0000010111011100; // vC= 1500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110010; // iC=-1678 
// vC = 14'b0000011000011110; // vC= 1566 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001011; // iC=-1589 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111001; // iC=-1543 
// vC = 14'b0000011001100110; // vC= 1638 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011000; // iC=-1576 
// vC = 14'b0000011010100000; // vC= 1696 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001000; // iC=-1592 
// vC = 14'b0000011001110101; // vC= 1653 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111100; // iC=-1732 
// vC = 14'b0000010111011000; // vC= 1496 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010001; // iC=-1647 
// vC = 14'b0000011001110001; // vC= 1649 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111110; // iC=-1666 
// vC = 14'b0000010111001110; // vC= 1486 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b0000011010000101; // vC= 1669 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000000; // iC=-1600 
// vC = 14'b0000010110000101; // vC= 1413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101010; // iC=-1814 
// vC = 14'b0000011001011011; // vC= 1627 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101111; // iC=-1745 
// vC = 14'b0000010101011001; // vC= 1369 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001101; // iC=-1715 
// vC = 14'b0000010111111010; // vC= 1530 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110000; // iC=-1872 
// vC = 14'b0000010111010101; // vC= 1493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b0000010111001111; // vC= 1487 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010110; // iC=-1642 
// vC = 14'b0000010110101011; // vC= 1451 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101111; // iC=-1745 
// vC = 14'b0000010111110100; // vC= 1524 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011000; // iC=-1896 
// vC = 14'b0000010100100001; // vC= 1313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100110; // iC=-1754 
// vC = 14'b0000011000010111; // vC= 1559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011111; // iC=-1697 
// vC = 14'b0000010100000010; // vC= 1282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001000; // iC=-1784 
// vC = 14'b0000011000001011; // vC= 1547 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010110; // iC=-1706 
// vC = 14'b0000010101000010; // vC= 1346 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010101; // iC=-1835 
// vC = 14'b0000010100011010; // vC= 1306 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110110; // iC=-1994 
// vC = 14'b0000011000000110; // vC= 1542 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000010101100000; // vC= 1376 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111001; // iC=-1927 
// vC = 14'b0000010111001000; // vC= 1480 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100111; // iC=-1753 
// vC = 14'b0000010011101011; // vC= 1259 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b0000010111101110; // vC= 1518 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100001; // iC=-1887 
// vC = 14'b0000010100010101; // vC= 1301 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001110; // iC=-1842 
// vC = 14'b0000010110111001; // vC= 1465 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b0000010110000000; // vC= 1408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000010111001001; // vC= 1481 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b0000010111000101; // vC= 1477 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111100; // iC=-1988 
// vC = 14'b0000010100110110; // vC= 1334 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010110; // iC=-1770 
// vC = 14'b0000010100001010; // vC= 1290 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b0000010010111011; // vC= 1211 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010100; // iC=-1900 
// vC = 14'b0000010101100110; // vC= 1382 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000101; // iC=-1851 
// vC = 14'b0000010010001100; // vC= 1164 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b0000010011110110; // vC= 1270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000100; // iC=-1980 
// vC = 14'b0000010011001000; // vC= 1224 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111001; // iC=-1863 
// vC = 14'b0000010101001100; // vC= 1356 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100001; // iC=-2079 
// vC = 14'b0000010001001010; // vC= 1098 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010100; // iC=-2028 
// vC = 14'b0000010011000100; // vC= 1220 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b0000010010001101; // vC= 1165 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011001; // iC=-1831 
// vC = 14'b0000010011010010; // vC= 1234 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011010; // iC=-1830 
// vC = 14'b0000010000101110; // vC= 1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b0000010000101011; // vC= 1067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000010010101000; // vC= 1192 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b0000010001011101; // vC= 1117 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010001; // iC=-2031 
// vC = 14'b0000010000010110; // vC= 1046 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b0000010100100101; // vC= 1317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000101; // iC=-2107 
// vC = 14'b0000010011110100; // vC= 1268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000010010110011; // vC= 1203 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000010010000111; // vC= 1159 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b0000010000010101; // vC= 1045 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000100; // iC=-1980 
// vC = 14'b0000010010101100; // vC= 1196 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100100; // iC=-1884 
// vC = 14'b0000010010001000; // vC= 1160 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b0000001111110000; // vC= 1008 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111011; // iC=-2117 
// vC = 14'b0000010000111111; // vC= 1087 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000000; // iC=-1856 
// vC = 14'b0000010010011100; // vC= 1180 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000010010011110; // vC= 1182 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b0000010010001101; // vC= 1165 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101001; // iC=-2135 
// vC = 14'b0000010011001011; // vC= 1227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011000; // iC=-1832 
// vC = 14'b0000010001111100; // vC= 1148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000010000100111; // vC= 1063 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101010; // iC=-1878 
// vC = 14'b0000010000110110; // vC= 1078 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b0000010001101100; // vC= 1132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b0000010010101001; // vC= 1193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b0000010001111100; // vC= 1148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b0000010000010010; // vC= 1042 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010111; // iC=-2153 
// vC = 14'b0000001101011110; // vC=  862 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000010001000100; // vC= 1092 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000010001000010; // vC= 1090 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101111; // iC=-2001 
// vC = 14'b0000001111001011; // vC=  971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010010; // iC=-2094 
// vC = 14'b0000001111101101; // vC= 1005 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b0000001111101101; // vC= 1005 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b0000001111110110; // vC= 1014 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b0000001111001011; // vC=  971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000101; // iC=-1915 
// vC = 14'b0000001111101110; // vC= 1006 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b0000001100101001; // vC=  809 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101001; // iC=-2071 
// vC = 14'b0000001100110011; // vC=  819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110001; // iC=-2127 
// vC = 14'b0000001110001011; // vC=  907 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b0000001110100101; // vC=  933 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b0000001110100111; // vC=  935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b0000001011100110; // vC=  742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000110; // iC=-2106 
// vC = 14'b0000001110100111; // vC=  935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111100; // iC=-1988 
// vC = 14'b0000001100000001; // vC=  769 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b0000001111101111; // vC= 1007 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b0000001110001101; // vC=  909 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010010; // iC=-1966 
// vC = 14'b0000001010101100; // vC=  684 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111000; // iC=-2120 
// vC = 14'b0000001101000110; // vC=  838 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b0000001100000010; // vC=  770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b0000001011010010; // vC=  722 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011011; // iC=-2085 
// vC = 14'b0000001110111010; // vC=  954 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b0000001110000111; // vC=  903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000010; // iC=-1918 
// vC = 14'b0000001110001010; // vC=  906 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000001; // iC=-1919 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111001; // iC=-2119 
// vC = 14'b0000001110011011; // vC=  923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110011; // iC=-1997 
// vC = 14'b0000001001011010; // vC=  602 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101000; // iC=-1880 
// vC = 14'b0000001110001000; // vC=  904 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b0000001100000010; // vC=  770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110110; // iC=-2122 
// vC = 14'b0000001010010001; // vC=  657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101101; // iC=-2067 
// vC = 14'b0000001011111111; // vC=  767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b0000001010001111; // vC=  655 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b0000001001000010; // vC=  578 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b0000001010111000; // vC=  696 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111111; // iC=-1985 
// vC = 14'b0000001101000011; // vC=  835 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100011; // iC=-2141 
// vC = 14'b0000001100011011; // vC=  795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010101; // iC=-2027 
// vC = 14'b0000001010100111; // vC=  679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b0000001010010000; // vC=  656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000001001001010; // vC=  586 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010010; // iC=-2158 
// vC = 14'b0000001001101011; // vC=  619 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000001000011111; // vC=  543 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b0000000111011101; // vC=  477 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b0000001010010010; // vC=  658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011110; // iC=-2018 
// vC = 14'b0000001000100010; // vC=  546 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111001; // iC=-2119 
// vC = 14'b0000001000000011; // vC=  515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101110; // iC=-2194 
// vC = 14'b0000001001100110; // vC=  614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b0000000111100001; // vC=  481 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b0000001011001011; // vC=  715 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000001010110010; // vC=  690 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100111; // iC=-2009 
// vC = 14'b0000000111111110; // vC=  510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000001001100111; // vC=  615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010111; // iC=-2153 
// vC = 14'b0000000101111110; // vC=  382 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111000; // iC=-2056 
// vC = 14'b0000001001110011; // vC=  627 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000110; // iC=-1914 
// vC = 14'b0000000111110110; // vC=  502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101111; // iC=-1873 
// vC = 14'b0000001000000111; // vC=  519 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110101; // iC=-2187 
// vC = 14'b0000000101111000; // vC=  376 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110001; // iC=-1935 
// vC = 14'b0000000110101001; // vC=  425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000000111100101; // vC=  485 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b0000000101110101; // vC=  373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b0000000110011110; // vC=  414 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000001; // iC=-1919 
// vC = 14'b0000000110010110; // vC=  406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b0000000110100111; // vC=  423 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000000111010111; // vC=  471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000000100011010; // vC=  282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111001; // iC=-1927 
// vC = 14'b0000000111100111; // vC=  487 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b0000001000010100; // vC=  532 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111101; // iC=-2179 
// vC = 14'b0000000100111000; // vC=  312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110011; // iC=-1869 
// vC = 14'b0000000100100011; // vC=  291 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001010; // iC=-1910 
// vC = 14'b0000000111000101; // vC=  453 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b0000000101000000; // vC=  320 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000000011000101; // vC=  197 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b0000000100010010; // vC=  274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b0000000111100001; // vC=  481 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000000100101000; // vC=  296 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001111; // iC=-2097 
// vC = 14'b0000000011001010; // vC=  202 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000000100000100; // vC=  260 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000101; // iC=-1915 
// vC = 14'b0000000101010011; // vC=  339 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b0000000010100000; // vC=  160 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110011; // iC=-2125 
// vC = 14'b0000000010000011; // vC=  131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111011; // iC=-2181 
// vC = 14'b0000000011010110; // vC=  214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b0000000110101001; // vC=  425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111010; // iC=-1862 
// vC = 14'b0000000011111101; // vC=  253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000000; // iC=-2176 
// vC = 14'b0000000100000110; // vC=  262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000100; // iC=-1980 
// vC = 14'b0000000001110100; // vC=  116 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b0000000101000111; // vC=  327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111000; // iC=-1928 
// vC = 14'b0000000110000101; // vC=  389 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000010; // iC=-1854 
// vC = 14'b0000000101111011; // vC=  379 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101111; // iC=-1937 
// vC = 14'b0000000101110101; // vC=  373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000000001001010; // vC=   74 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000000010000010; // vC=  130 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b0000000001010100; // vC=   84 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000000010001101; // vC=  141 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b0000000011011100; // vC=  220 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101010; // iC=-1878 
// vC = 14'b0000000100110000; // vC=  304 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011000; // iC=-2152 
// vC = 14'b0000000001001010; // vC=   74 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111010; // iC=-1862 
// vC = 14'b0000000011101101; // vC=  237 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b0000000011011011; // vC=  219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010000; // iC=-1904 
// vC = 14'b0000000000011011; // vC=   27 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b0000000011100011; // vC=  227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000000010101100; // vC=  172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111000; // iC=-1928 
// vC = 14'b0000000001001010; // vC=   74 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011001; // iC=-2087 
// vC = 14'b1111111110101111; // vC=  -81 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000001; // iC=-1855 
// vC = 14'b0000000001011111; // vC=   95 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b1111111111011001; // vC=  -39 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b0000000001111111; // vC=  127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000100; // iC=-1852 
// vC = 14'b0000000001110001; // vC=  113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011000; // iC=-2152 
// vC = 14'b0000000001010101; // vC=   85 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b1111111110101010; // vC=  -86 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b0000000000010000; // vC=   16 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000010; // iC=-1854 
// vC = 14'b1111111101110110; // vC= -138 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b1111111111101000; // vC=  -24 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b0000000010001111; // vC=  143 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b1111111111110100; // vC=  -12 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010110; // iC=-2090 
// vC = 14'b1111111111010111; // vC=  -41 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b0000000010000100; // vC=  132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111001; // iC=-1991 
// vC = 14'b1111111110110001; // vC=  -79 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100001; // iC=-2079 
// vC = 14'b0000000000110000; // vC=   48 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b1111111110110001; // vC=  -79 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b1111111100110000; // vC= -208 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b0000000000000010; // vC=    2 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000100; // iC=-2044 
// vC = 14'b0000000001000101; // vC=   69 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b1111111111110110; // vC=  -10 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b1111111111011010; // vC=  -38 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000011; // iC=-1853 
// vC = 14'b0000000000000010; // vC=    2 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110110; // iC=-2122 
// vC = 14'b1111111011111100; // vC= -260 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001111; // iC=-1841 
// vC = 14'b1111111100011011; // vC= -229 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b1111111100100011; // vC= -221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010010; // iC=-1966 
// vC = 14'b1111111011111101; // vC= -259 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000000; // iC=-1856 
// vC = 14'b1111111110101110; // vC=  -82 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111101; // iC=-1859 
// vC = 14'b1111111111011100; // vC=  -36 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b1111111101011111; // vC= -161 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101001; // iC=-2007 
// vC = 14'b1111111100010110; // vC= -234 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b1111111101001001; // vC= -183 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b1111111101010111; // vC= -169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001010; // iC=-1782 
// vC = 14'b1111111011000101; // vC= -315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b1111111010101101; // vC= -339 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110011; // iC=-1933 
// vC = 14'b1111111110100110; // vC=  -90 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b1111111101010011; // vC= -173 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b1111111101100010; // vC= -158 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111010; // iC=-1862 
// vC = 14'b1111111101110011; // vC= -141 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b1111111011000111; // vC= -313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b1111111101110010; // vC= -142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100010; // iC=-1822 
// vC = 14'b1111111110010001; // vC= -111 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b1111111100000001; // vC= -255 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110100; // iC=-1932 
// vC = 14'b1111111001111010; // vC= -390 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b1111111101010110; // vC= -170 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b1111111011110000; // vC= -272 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b1111111011110011; // vC= -269 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100011; // iC=-1757 
// vC = 14'b1111111101100100; // vC= -156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001100; // iC=-1908 
// vC = 14'b1111111000101110; // vC= -466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b1111111001111101; // vC= -387 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101110; // iC=-1810 
// vC = 14'b1111111011100101; // vC= -283 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000110; // iC=-1786 
// vC = 14'b1111111010100001; // vC= -351 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b1111111001101000; // vC= -408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b1111111001100010; // vC= -414 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110010; // iC=-2062 
// vC = 14'b1111111010111110; // vC= -322 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b1111110111100000; // vC= -544 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110011; // iC=-1805 
// vC = 14'b1111111001011111; // vC= -417 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001111; // iC=-1777 
// vC = 14'b1111111001011000; // vC= -424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111100; // iC=-1732 
// vC = 14'b1111111000011110; // vC= -482 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b1111111000000000; // vC= -512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b1111111011110010; // vC= -270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111111011010001; // vC= -303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b1111111011001111; // vC= -305 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b1111111010001001; // vC= -375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111111001000010; // vC= -446 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001111; // iC=-1777 
// vC = 14'b1111111000010100; // vC= -492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b1111111010100010; // vC= -350 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b1111110111100100; // vC= -540 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010111; // iC=-2025 
// vC = 14'b1111111001001100; // vC= -436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b1111110110101101; // vC= -595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b1111110111000101; // vC= -571 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011000; // iC=-1896 
// vC = 14'b1111110110010010; // vC= -622 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011001; // iC=-1895 
// vC = 14'b1111110110001011; // vC= -629 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001100; // iC=-1908 
// vC = 14'b1111110111101000; // vC= -536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110100; // iC=-1932 
// vC = 14'b1111110111111111; // vC= -513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b1111111010000101; // vC= -379 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011101; // iC=-1763 
// vC = 14'b1111110111101101; // vC= -531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010010; // iC=-1710 
// vC = 14'b1111110110000011; // vC= -637 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100111; // iC=-1881 
// vC = 14'b1111110110001010; // vC= -630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101000; // iC=-1688 
// vC = 14'b1111111000011000; // vC= -488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010010; // iC=-1838 
// vC = 14'b1111111001001010; // vC= -438 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100000; // iC=-1952 
// vC = 14'b1111111000100111; // vC= -473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111111; // iC=-1793 
// vC = 14'b1111110111000011; // vC= -573 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101110; // iC=-1810 
// vC = 14'b1111110110101101; // vC= -595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011000; // iC=-1768 
// vC = 14'b1111110101011010; // vC= -678 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000101; // iC=-1915 
// vC = 14'b1111111000101001; // vC= -471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111011; // iC=-1733 
// vC = 14'b1111110101011001; // vC= -679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010000; // iC=-1776 
// vC = 14'b1111110110001011; // vC= -629 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b1111110011100001; // vC= -799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101010; // iC=-1686 
// vC = 14'b1111110100111010; // vC= -710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b1111110101100100; // vC= -668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100000; // iC=-1824 
// vC = 14'b1111110110111001; // vC= -583 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000111; // iC=-1785 
// vC = 14'b1111110110011011; // vC= -613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b1111110101101111; // vC= -657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001010; // iC=-1654 
// vC = 14'b1111110101001100; // vC= -692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001110; // iC=-1778 
// vC = 14'b1111110011110101; // vC= -779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101000; // iC=-1816 
// vC = 14'b1111110101101100; // vC= -660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111010; // iC=-1734 
// vC = 14'b1111110110111011; // vC= -581 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100110; // iC=-1818 
// vC = 14'b1111110110001100; // vC= -628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100011; // iC=-1821 
// vC = 14'b1111110101000000; // vC= -704 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100101; // iC=-1691 
// vC = 14'b1111110010111010; // vC= -838 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001100; // iC=-1716 
// vC = 14'b1111110101011110; // vC= -674 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100110; // iC=-1690 
// vC = 14'b1111110100001001; // vC= -759 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000001; // iC=-1727 
// vC = 14'b1111110100010001; // vC= -751 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111001; // iC=-1799 
// vC = 14'b1111110001101111; // vC= -913 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011001; // iC=-1767 
// vC = 14'b1111110101010110; // vC= -682 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001100; // iC=-1588 
// vC = 14'b1111110011000001; // vC= -831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010001; // iC=-1839 
// vC = 14'b1111110101101001; // vC= -663 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000011; // iC=-1789 
// vC = 14'b1111110010110001; // vC= -847 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111011; // iC=-1669 
// vC = 14'b1111110010100110; // vC= -858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011010; // iC=-1638 
// vC = 14'b1111110100000101; // vC= -763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001001; // iC=-1591 
// vC = 14'b1111110100001011; // vC= -757 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100000; // iC=-1760 
// vC = 14'b1111110100000011; // vC= -765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000001; // iC=-1663 
// vC = 14'b1111110001001100; // vC= -948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000000; // iC=-1792 
// vC = 14'b1111110010100101; // vC= -859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010101; // iC=-1707 
// vC = 14'b1111110001101111; // vC= -913 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011111; // iC=-1697 
// vC = 14'b1111110000100000; // vC= -992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100001; // iC=-1759 
// vC = 14'b1111110001110110; // vC= -906 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101011; // iC=-1749 
// vC = 14'b1111110100011011; // vC= -741 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010011; // iC=-1645 
// vC = 14'b1111110011111001; // vC= -775 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100111; // iC=-1817 
// vC = 14'b1111110100101011; // vC= -725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100011; // iC=-1821 
// vC = 14'b1111110000110000; // vC= -976 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010000; // iC=-1520 
// vC = 14'b1111110011011110; // vC= -802 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100011; // iC=-1693 
// vC = 14'b1111110001101100; // vC= -916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011101; // iC=-1571 
// vC = 14'b1111110001000101; // vC= -955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000101; // iC=-1787 
// vC = 14'b1111101111011110; // vC=-1058 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111000; // iC=-1608 
// vC = 14'b1111110010100110; // vC= -858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100001; // iC=-1503 
// vC = 14'b1111110011010000; // vC= -816 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001010; // iC=-1782 
// vC = 14'b1111110010100110; // vC= -858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111000; // iC=-1672 
// vC = 14'b1111101111111100; // vC=-1028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110110; // iC=-1674 
// vC = 14'b1111101110110010; // vC=-1102 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010010; // iC=-1646 
// vC = 14'b1111110000000101; // vC=-1019 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000011; // iC=-1725 
// vC = 14'b1111110011000001; // vC= -831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101000; // iC=-1752 
// vC = 14'b1111110001100010; // vC= -926 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010110; // iC=-1514 
// vC = 14'b1111101110011100; // vC=-1124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110000; // iC=-1680 
// vC = 14'b1111101111001111; // vC=-1073 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000101; // iC=-1531 
// vC = 14'b1111110001011000; // vC= -936 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111110; // iC=-1666 
// vC = 14'b1111101111110011; // vC=-1037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101100; // iC=-1620 
// vC = 14'b1111101110101101; // vC=-1107 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111100; // iC=-1540 
// vC = 14'b1111110000011111; // vC= -993 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000111; // iC=-1465 
// vC = 14'b1111110000000001; // vC=-1023 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110101; // iC=-1547 
// vC = 14'b1111110010010001; // vC= -879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000000; // iC=-1472 
// vC = 14'b1111101110010100; // vC=-1132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100111; // iC=-1689 
// vC = 14'b1111101111100011; // vC=-1053 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100011; // iC=-1629 
// vC = 14'b1111110001011110; // vC= -930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100000; // iC=-1696 
// vC = 14'b1111110010001011; // vC= -885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110111; // iC=-1737 
// vC = 14'b1111101110101101; // vC=-1107 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010010; // iC=-1518 
// vC = 14'b1111110001100011; // vC= -925 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000000; // iC=-1600 
// vC = 14'b1111101110000110; // vC=-1146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010100; // iC=-1452 
// vC = 14'b1111101111100101; // vC=-1051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101100; // iC=-1556 
// vC = 14'b1111101110111111; // vC=-1089 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110010; // iC=-1678 
// vC = 14'b1111101101000010; // vC=-1214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011011; // iC=-1509 
// vC = 14'b1111101101001000; // vC=-1208 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100100; // iC=-1500 
// vC = 14'b1111110000011101; // vC= -995 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101000; // iC=-1560 
// vC = 14'b1111101110011100; // vC=-1124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011000; // iC=-1384 
// vC = 14'b1111101101010000; // vC=-1200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100011; // iC=-1693 
// vC = 14'b1111101101111000; // vC=-1160 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000000; // iC=-1600 
// vC = 14'b1111101111011110; // vC=-1058 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000011; // iC=-1405 
// vC = 14'b1111101111111101; // vC=-1027 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100110; // iC=-1690 
// vC = 14'b1111101101110010; // vC=-1166 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100111; // iC=-1561 
// vC = 14'b1111101100111110; // vC=-1218 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100101; // iC=-1563 
// vC = 14'b1111110000100000; // vC= -992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011100; // iC=-1380 
// vC = 14'b1111101110110111; // vC=-1097 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100101; // iC=-1627 
// vC = 14'b1111101111101101; // vC=-1043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100100; // iC=-1436 
// vC = 14'b1111101111100000; // vC=-1056 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011110; // iC=-1442 
// vC = 14'b1111101111100110; // vC=-1050 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001010; // iC=-1398 
// vC = 14'b1111101110011101; // vC=-1123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110100; // iC=-1356 
// vC = 14'b1111101110110010; // vC=-1102 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111000; // iC=-1480 
// vC = 14'b1111101011010111; // vC=-1321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000111; // iC=-1593 
// vC = 14'b1111101110010001; // vC=-1135 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010011; // iC=-1581 
// vC = 14'b1111101011111001; // vC=-1287 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101110; // iC=-1426 
// vC = 14'b1111101100111011; // vC=-1221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111011; // iC=-1605 
// vC = 14'b1111101110101010; // vC=-1110 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000011; // iC=-1533 
// vC = 14'b1111101011010001; // vC=-1327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111010; // iC=-1414 
// vC = 14'b1111101100010000; // vC=-1264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101101; // iC=-1299 
// vC = 14'b1111101110101000; // vC=-1112 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110000; // iC=-1424 
// vC = 14'b1111101010100011; // vC=-1373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010000; // iC=-1328 
// vC = 14'b1111101100000111; // vC=-1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000111; // iC=-1529 
// vC = 14'b1111101011100010; // vC=-1310 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101100; // iC=-1492 
// vC = 14'b1111101110010011; // vC=-1133 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101011; // iC=-1557 
// vC = 14'b1111101001111011; // vC=-1413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001001; // iC=-1527 
// vC = 14'b1111101001101110; // vC=-1426 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001111; // iC=-1457 
// vC = 14'b1111101100111011; // vC=-1221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010010; // iC=-1262 
// vC = 14'b1111101110000100; // vC=-1148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011110; // iC=-1378 
// vC = 14'b1111101101101100; // vC=-1172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001111; // iC=-1457 
// vC = 14'b1111101110001000; // vC=-1144 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000100; // iC=-1276 
// vC = 14'b1111101010101011; // vC=-1365 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100000; // iC=-1312 
// vC = 14'b1111101010001001; // vC=-1399 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001110; // iC=-1266 
// vC = 14'b1111101011110010; // vC=-1294 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010011; // iC=-1389 
// vC = 14'b1111101100111010; // vC=-1222 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011101; // iC=-1443 
// vC = 14'b1111101100100011; // vC=-1245 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111001; // iC=-1415 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100000; // iC=-1248 
// vC = 14'b1111101101000101; // vC=-1211 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000111; // iC=-1273 
// vC = 14'b1111101010000111; // vC=-1401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011011; // iC=-1253 
// vC = 14'b1111101010100100; // vC=-1372 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000011; // iC=-1213 
// vC = 14'b1111101101000011; // vC=-1213 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000010; // iC=-1342 
// vC = 14'b1111101100111100; // vC=-1220 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101000; // iC=-1432 
// vC = 14'b1111101100011101; // vC=-1251 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101011; // iC=-1429 
// vC = 14'b1111101010111010; // vC=-1350 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101100; // iC=-1236 
// vC = 14'b1111101011110111; // vC=-1289 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101010; // iC=-1430 
// vC = 14'b1111101001101000; // vC=-1432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001001; // iC=-1335 
// vC = 14'b1111101011011101; // vC=-1315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011001; // iC=-1383 
// vC = 14'b1111101001011010; // vC=-1446 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110011; // iC=-1293 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001001; // iC=-1335 
// vC = 14'b1111101000010101; // vC=-1515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001100; // iC=-1460 
// vC = 14'b1111101000101011; // vC=-1493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101111; // iC=-1169 
// vC = 14'b1111101001011011; // vC=-1445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000100; // iC=-1148 
// vC = 14'b1111101100000110; // vC=-1274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000011; // iC=-1277 
// vC = 14'b1111101001101111; // vC=-1425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100000; // iC=-1248 
// vC = 14'b1111101011001001; // vC=-1335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110000; // iC=-1424 
// vC = 14'b1111100111001111; // vC=-1585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110110; // iC=-1418 
// vC = 14'b1111101010000010; // vC=-1406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101001; // iC=-1367 
// vC = 14'b1111101011000111; // vC=-1337 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001001; // iC=-1335 
// vC = 14'b1111100111111010; // vC=-1542 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000111; // iC=-1401 
// vC = 14'b1111100111100001; // vC=-1567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001001; // iC=-1143 
// vC = 14'b1111101001000110; // vC=-1466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011000; // iC=-1320 
// vC = 14'b1111101010000101; // vC=-1403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001111; // iC=-1265 
// vC = 14'b1111101001011010; // vC=-1446 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001100; // iC=-1268 
// vC = 14'b1111100110110100; // vC=-1612 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000011; // iC=-1213 
// vC = 14'b1111101010110100; // vC=-1356 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010100; // iC=-1068 
// vC = 14'b1111101001011000; // vC=-1448 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100110; // iC=-1178 
// vC = 14'b1111100110110111; // vC=-1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010001; // iC=-1263 
// vC = 14'b1111101000011111; // vC=-1505 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011001; // iC=-1191 
// vC = 14'b1111100110100101; // vC=-1627 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011100; // iC=-1060 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100111; // iC=-1177 
// vC = 14'b1111100111001001; // vC=-1591 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010100; // iC=-1260 
// vC = 14'b1111100110000111; // vC=-1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100010; // iC=-1118 
// vC = 14'b1111100111001011; // vC=-1589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010110; // iC=-1258 
// vC = 14'b1111101000110101; // vC=-1483 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000100; // iC=-1084 
// vC = 14'b1111100110100000; // vC=-1632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010110; // iC=-1066 
// vC = 14'b1111100101111010; // vC=-1670 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000011; // iC=-1021 
// vC = 14'b1111101010001001; // vC=-1399 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010110; // iC=-1194 
// vC = 14'b1111101000101110; // vC=-1490 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000111; // iC=-1209 
// vC = 14'b1111100110110010; // vC=-1614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000010; // iC=-1086 
// vC = 14'b1111100110110111; // vC=-1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100010; // iC=-1118 
// vC = 14'b1111100110010110; // vC=-1642 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110001; // iC=-1295 
// vC = 14'b1111101000000000; // vC=-1536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110100; // iC=-1036 
// vC = 14'b1111100111000010; // vC=-1598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110111; // iC=-1097 
// vC = 14'b1111101001010000; // vC=-1456 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111010; // iC=-1030 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111100; // iC=-1092 
// vC = 14'b1111100101101111; // vC=-1681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000110; // iC=-1210 
// vC = 14'b1111100110000110; // vC=-1658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000010; // iC=-1150 
// vC = 14'b1111101001011011; // vC=-1445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011000; // iC=-1064 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100000; // iC=-1184 
// vC = 14'b1111100101111001; // vC=-1671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000111; // iC=-1081 
// vC = 14'b1111100101111111; // vC=-1665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011100; // iC=-1188 
// vC = 14'b1111100101011100; // vC=-1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110101; // iC=-1035 
// vC = 14'b1111100110101100; // vC=-1620 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111000; // iC=-1160 
// vC = 14'b1111100111101011; // vC=-1557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b1111100111110010; // vC=-1550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111001; // iC=-1031 
// vC = 14'b1111101000100100; // vC=-1500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011001; // iC= -999 
// vC = 14'b1111100111111101; // vC=-1539 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010110; // iC=-1194 
// vC = 14'b1111100101100111; // vC=-1689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111011; // iC=-1093 
// vC = 14'b1111100011111010; // vC=-1798 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011101; // iC=-1187 
// vC = 14'b1111100100100110; // vC=-1754 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111110; // iC=-1154 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111010; // iC=-1094 
// vC = 14'b1111100100001010; // vC=-1782 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001000; // iC=-1144 
// vC = 14'b1111101000011110; // vC=-1506 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001100; // iC=-1140 
// vC = 14'b1111100011110100; // vC=-1804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101010; // iC=-1046 
// vC = 14'b1111101000000110; // vC=-1530 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001110; // iC= -946 
// vC = 14'b1111100101011000; // vC=-1704 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101011; // iC=-1045 
// vC = 14'b1111100101111111; // vC=-1665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100010; // iC=-1054 
// vC = 14'b1111100100010111; // vC=-1769 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011110; // iC= -866 
// vC = 14'b1111100111101110; // vC=-1554 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001110; // iC= -882 
// vC = 14'b1111100111001011; // vC=-1589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001011; // iC=-1077 
// vC = 14'b1111100101100100; // vC=-1692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110000; // iC=-1104 
// vC = 14'b1111100111000100; // vC=-1596 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111111; // iC=-1025 
// vC = 14'b1111100101100101; // vC=-1691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100001; // iC= -863 
// vC = 14'b1111100101101111; // vC=-1681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000101; // iC= -827 
// vC = 14'b1111100011001110; // vC=-1842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100010; // iC=-1054 
// vC = 14'b1111100100100001; // vC=-1759 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000101; // iC=-1019 
// vC = 14'b1111100111001101; // vC=-1587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111011; // iC= -901 
// vC = 14'b1111100101000100; // vC=-1724 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110010; // iC= -846 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001010; // iC= -886 
// vC = 14'b1111100101111110; // vC=-1666 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000110; // iC= -954 
// vC = 14'b1111100101100100; // vC=-1692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001011; // iC= -885 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111110; // iC= -770 
// vC = 14'b1111100101010001; // vC=-1711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000011; // iC=-1021 
// vC = 14'b1111100111011100; // vC=-1572 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010011; // iC= -877 
// vC = 14'b1111100111000111; // vC=-1593 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011001; // iC= -871 
// vC = 14'b1111100011001111; // vC=-1841 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001111; // iC= -817 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111001; // iC= -839 
// vC = 14'b1111100110101101; // vC=-1619 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101000; // iC= -984 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111010; // iC= -710 
// vC = 14'b1111100010100101; // vC=-1883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000100; // iC= -828 
// vC = 14'b1111100101110110; // vC=-1674 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110101; // iC= -907 
// vC = 14'b1111100110000101; // vC=-1659 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111110; // iC= -834 
// vC = 14'b1111100110110001; // vC=-1615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100100; // iC= -988 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010000; // iC= -816 
// vC = 14'b1111100010110010; // vC=-1870 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011001; // iC= -935 
// vC = 14'b1111100010110011; // vC=-1869 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011111; // iC= -801 
// vC = 14'b1111100001111011; // vC=-1925 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101101; // iC= -723 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011110; // iC= -930 
// vC = 14'b1111100010111100; // vC=-1860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000011; // iC= -701 
// vC = 14'b1111100001101110; // vC=-1938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010110; // iC= -874 
// vC = 14'b1111100001111001; // vC=-1927 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001010; // iC= -886 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011101; // iC= -931 
// vC = 14'b1111100011010001; // vC=-1839 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011100; // iC= -740 
// vC = 14'b1111100001101110; // vC=-1938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111000; // iC= -840 
// vC = 14'b1111100100100010; // vC=-1758 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011010; // iC= -678 
// vC = 14'b1111100101000001; // vC=-1727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010100; // iC= -620 
// vC = 14'b1111100010110011; // vC=-1869 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111111; // iC= -769 
// vC = 14'b1111100101010100; // vC=-1708 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111001; // iC= -583 
// vC = 14'b1111100011101000; // vC=-1816 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101111; // iC= -785 
// vC = 14'b1111100011100100; // vC=-1820 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111101; // iC= -643 
// vC = 14'b1111100001111100; // vC=-1924 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010000; // iC= -688 
// vC = 14'b1111100011010100; // vC=-1836 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101011; // iC= -853 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100000; // iC= -800 
// vC = 14'b1111100010110010; // vC=-1870 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100010; // iC= -862 
// vC = 14'b1111100011111011; // vC=-1797 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000101; // iC= -699 
// vC = 14'b1111100010011100; // vC=-1892 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101101; // iC= -787 
// vC = 14'b1111100011100010; // vC=-1822 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110100; // iC= -780 
// vC = 14'b1111100101101110; // vC=-1682 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100100; // iC= -540 
// vC = 14'b1111100011010000; // vC=-1840 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110010; // iC= -590 
// vC = 14'b1111100001110101; // vC=-1931 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011001; // iC= -679 
// vC = 14'b1111100010010100; // vC=-1900 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111110; // iC= -770 
// vC = 14'b1111100000110100; // vC=-1996 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010100; // iC= -684 
// vC = 14'b1111100001000111; // vC=-1977 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100101; // iC= -667 
// vC = 14'b1111100100101100; // vC=-1748 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001110; // iC= -690 
// vC = 14'b1111100000100100; // vC=-2012 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001011; // iC= -501 
// vC = 14'b1111100010011000; // vC=-1896 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111001; // iC= -455 
// vC = 14'b1111100010011001; // vC=-1895 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000111; // iC= -697 
// vC = 14'b1111100010100100; // vC=-1884 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101110; // iC= -722 
// vC = 14'b1111100011110011; // vC=-1805 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110000; // iC= -656 
// vC = 14'b1111100001010111; // vC=-1961 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101000; // iC= -600 
// vC = 14'b1111100000011111; // vC=-2017 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011011; // iC= -613 
// vC = 14'b1111100011010000; // vC=-1840 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001011; // iC= -501 
// vC = 14'b1111100001000010; // vC=-1982 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001011; // iC= -437 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001101; // iC= -499 
// vC = 14'b1111100010011110; // vC=-1890 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100101; // iC= -347 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010010; // iC= -366 
// vC = 14'b1111100011001011; // vC=-1845 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000010; // iC= -446 
// vC = 14'b1111100011000100; // vC=-1852 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100010; // iC= -414 
// vC = 14'b1111100000010101; // vC=-2027 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001110; // iC= -562 
// vC = 14'b1111100000100001; // vC=-2015 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111110011; // iC= -525 
// vC = 14'b1111100010101101; // vC=-1875 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100010; // iC= -414 
// vC = 14'b1111100001011101; // vC=-1955 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010011; // iC= -365 
// vC = 14'b1111100000101110; // vC=-2002 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101001; // iC= -535 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001110; // iC= -498 
// vC = 14'b1111100000000101; // vC=-2043 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100100; // iC= -412 
// vC = 14'b1111100001100000; // vC=-1952 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010001; // iC= -303 
// vC = 14'b1111100010001101; // vC=-1907 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011110110; // iC= -266 
// vC = 14'b1111100000010111; // vC=-2025 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010111; // iC= -361 
// vC = 14'b1111100001011110; // vC=-1954 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001010; // iC= -182 
// vC = 14'b1111100011010010; // vC=-1838 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011111; // iC= -289 
// vC = 14'b1111100000011101; // vC=-2019 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010010; // iC= -366 
// vC = 14'b1111100100001000; // vC=-1784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011110001; // iC= -271 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011011; // iC= -229 
// vC = 14'b1111100011110010; // vC=-1806 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011011; // iC= -293 
// vC = 14'b1111100001111100; // vC=-1924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111111; // iC= -193 
// vC = 14'b1111100100101001; // vC=-1751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010100; // iC= -108 
// vC = 14'b1111100000111101; // vC=-1987 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101100; // iC= -212 
// vC = 14'b1111100011010111; // vC=-1833 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101001; // iC= -215 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010001; // iC= -175 
// vC = 14'b1111100001010011; // vC=-1965 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000100; // iC= -252 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101101; // iC= -275 
// vC = 14'b1111100000110001; // vC=-1999 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011100; // iC=   28 
// vC = 14'b1111100010011011; // vC=-1893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100011; // iC= -157 
// vC = 14'b1111100001111011; // vC=-1925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000110; // iC=    6 
// vC = 14'b1111100011111100; // vC=-1796 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000011; // iC=    3 
// vC = 14'b1111100001110001; // vC=-1935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001000; // iC=   72 
// vC = 14'b1111100001101111; // vC=-1937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011101; // iC=   29 
// vC = 14'b1111100010000100; // vC=-1916 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111111; // iC=   -1 
// vC = 14'b1111100000001101; // vC=-2035 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001100; // iC=   76 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010011; // iC=  147 
// vC = 14'b1111100000001101; // vC=-2035 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011011111; // iC=  223 
// vC = 14'b1111100000101001; // vC=-2007 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101111; // iC=  239 
// vC = 14'b1111100010101001; // vC=-1879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110101; // iC=  245 
// vC = 14'b1111100010011111; // vC=-1889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000101; // iC=  261 
// vC = 14'b1111100000100111; // vC=-2009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001101; // iC=  269 
// vC = 14'b1111100010111110; // vC=-1858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011101; // iC=   29 
// vC = 14'b1111100000001111; // vC=-2033 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010111; // iC=  279 
// vC = 14'b1111011111111111; // vC=-2049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111100; // iC=  188 
// vC = 14'b1111100011110110; // vC=-1802 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010001; // iC=  209 
// vC = 14'b1111100011001100; // vC=-1844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011100; // iC=  156 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000001; // iC=  385 
// vC = 14'b1111100000001110; // vC=-2034 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101111; // iC=  367 
// vC = 14'b1111100000001011; // vC=-2037 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101000; // iC=  360 
// vC = 14'b1111100001101011; // vC=-1941 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101001; // iC=  489 
// vC = 14'b1111100100001001; // vC=-1783 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100000; // iC=  416 
// vC = 14'b1111100100100110; // vC=-1754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101110; // iC=  366 
// vC = 14'b1111100001001011; // vC=-1973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111111; // iC=  511 
// vC = 14'b1111100000100100; // vC=-2012 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000000; // iC=  512 
// vC = 14'b1111100010000110; // vC=-1914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101010; // iC=  426 
// vC = 14'b1111100100011010; // vC=-1766 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100111; // iC=  423 
// vC = 14'b1111100010011111; // vC=-1889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110001; // iC=  625 
// vC = 14'b1111100010111101; // vC=-1859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100000; // iC=  416 
// vC = 14'b1111100010110000; // vC=-1872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000110; // iC=  646 
// vC = 14'b1111100010000111; // vC=-1913 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011011; // iC=  475 
// vC = 14'b1111100011001111; // vC=-1841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110000; // iC=  496 
// vC = 14'b1111100100101011; // vC=-1749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100011; // iC=  739 
// vC = 14'b1111100101010001; // vC=-1711 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110101; // iC=  565 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000111; // iC=  583 
// vC = 14'b1111100100000110; // vC=-1786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110100; // iC=  692 
// vC = 14'b1111100011000101; // vC=-1851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110100; // iC=  692 
// vC = 14'b1111100011111001; // vC=-1799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000001; // iC=  833 
// vC = 14'b1111100101011011; // vC=-1701 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011111; // iC=  799 
// vC = 14'b1111100001010110; // vC=-1962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111111; // iC=  639 
// vC = 14'b1111100001010000; // vC=-1968 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111111; // iC=  767 
// vC = 14'b1111100011101100; // vC=-1812 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010111; // iC=  791 
// vC = 14'b1111100100111100; // vC=-1732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010000; // iC=  976 
// vC = 14'b1111100101001001; // vC=-1719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000010; // iC=  834 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110011; // iC=  947 
// vC = 14'b1111100100110010; // vC=-1742 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110000; // iC= 1072 
// vC = 14'b1111100011000011; // vC=-1853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010110; // iC=  854 
// vC = 14'b1111100101011110; // vC=-1698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111000; // iC= 1016 
// vC = 14'b1111100001110110; // vC=-1930 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001000; // iC=  904 
// vC = 14'b1111100011111001; // vC=-1799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101010; // iC=  938 
// vC = 14'b1111100011111100; // vC=-1796 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100101; // iC=  933 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100100; // iC= 1188 
// vC = 14'b1111100110011111; // vC=-1633 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011100; // iC=  924 
// vC = 14'b1111100101001111; // vC=-1713 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010111; // iC= 1047 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001111; // iC= 1039 
// vC = 14'b1111100100111100; // vC=-1732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101010; // iC= 1258 
// vC = 14'b1111100100101010; // vC=-1750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100000; // iC= 1056 
// vC = 14'b1111100110010000; // vC=-1648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100101; // iC= 1253 
// vC = 14'b1111100101110111; // vC=-1673 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110111; // iC= 1207 
// vC = 14'b1111100101111010; // vC=-1670 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010111; // iC= 1367 
// vC = 14'b1111100011000000; // vC=-1856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101011; // iC= 1067 
// vC = 14'b1111100110111100; // vC=-1604 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000010; // iC= 1218 
// vC = 14'b1111100111000100; // vC=-1596 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101100; // iC= 1196 
// vC = 14'b1111100011001000; // vC=-1848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001011; // iC= 1291 
// vC = 14'b1111100011001111; // vC=-1841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110101; // iC= 1141 
// vC = 14'b1111100110011101; // vC=-1635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001111; // iC= 1231 
// vC = 14'b1111100110011101; // vC=-1635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000001; // iC= 1409 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101110; // iC= 1390 
// vC = 14'b1111100100010100; // vC=-1772 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111110; // iC= 1342 
// vC = 14'b1111100011101010; // vC=-1814 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111010; // iC= 1466 
// vC = 14'b1111100101110110; // vC=-1674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111101; // iC= 1533 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100001; // iC= 1313 
// vC = 14'b1111100110001110; // vC=-1650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011001; // iC= 1369 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010000; // iC= 1424 
// vC = 14'b1111101000010000; // vC=-1520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101001; // iC= 1577 
// vC = 14'b1111100101001010; // vC=-1718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101101; // iC= 1389 
// vC = 14'b1111101000110001; // vC=-1487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110001; // iC= 1393 
// vC = 14'b1111100100101001; // vC=-1751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111000; // iC= 1528 
// vC = 14'b1111100101001010; // vC=-1718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000000; // iC= 1536 
// vC = 14'b1111100111111110; // vC=-1538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100111; // iC= 1575 
// vC = 14'b1111100100011111; // vC=-1761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100011; // iC= 1571 
// vC = 14'b1111100111010001; // vC=-1583 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100001; // iC= 1697 
// vC = 14'b1111101001011110; // vC=-1442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010010; // iC= 1554 
// vC = 14'b1111101001011001; // vC=-1447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101010; // iC= 1642 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100101; // iC= 1509 
// vC = 14'b1111100101111100; // vC=-1668 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110001; // iC= 1585 
// vC = 14'b1111100111111000; // vC=-1544 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101111; // iC= 1775 
// vC = 14'b1111100111101111; // vC=-1553 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111000; // iC= 1656 
// vC = 14'b1111100110111101; // vC=-1603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101100; // iC= 1580 
// vC = 14'b1111100101101101; // vC=-1683 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110110; // iC= 1718 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000110; // iC= 1670 
// vC = 14'b1111101001110111; // vC=-1417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010100; // iC= 1620 
// vC = 14'b1111100111011000; // vC=-1576 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000011; // iC= 1667 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101010; // iC= 1834 
// vC = 14'b1111101010110110; // vC=-1354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100011; // iC= 1635 
// vC = 14'b1111101000011100; // vC=-1508 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111001; // iC= 1657 
// vC = 14'b1111100111101010; // vC=-1558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011001; // iC= 1817 
// vC = 14'b1111100110011110; // vC=-1634 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010011; // iC= 1747 
// vC = 14'b1111101000010101; // vC=-1515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101011; // iC= 1899 
// vC = 14'b1111101011001001; // vC=-1335 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110101; // iC= 1653 
// vC = 14'b1111100110100110; // vC=-1626 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010001; // iC= 1873 
// vC = 14'b1111101010111001; // vC=-1351 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011110; // iC= 1822 
// vC = 14'b1111101000000110; // vC=-1530 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000101; // iC= 1669 
// vC = 14'b1111101011011011; // vC=-1317 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111011; // iC= 1723 
// vC = 14'b1111101010010101; // vC=-1387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010010; // iC= 1682 
// vC = 14'b1111101001110011; // vC=-1421 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011011; // iC= 1755 
// vC = 14'b1111101100010110; // vC=-1258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010011; // iC= 1811 
// vC = 14'b1111101011011011; // vC=-1317 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b1111101010011101; // vC=-1379 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b1111101010010000; // vC=-1392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010110; // iC= 1814 
// vC = 14'b1111101100001110; // vC=-1266 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b1111101100100110; // vC=-1242 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001111; // iC= 1807 
// vC = 14'b1111101010110010; // vC=-1358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110110; // iC= 1974 
// vC = 14'b1111101101000101; // vC=-1211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101010; // iC= 1770 
// vC = 14'b1111101101001010; // vC=-1206 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b1111101101011001; // vC=-1191 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011000; // iC= 1880 
// vC = 14'b1111101001011010; // vC=-1446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101010; // iC= 1834 
// vC = 14'b1111101101100000; // vC=-1184 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b1111101001110000; // vC=-1424 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b1111101101101100; // vC=-1172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100011; // iC= 2083 
// vC = 14'b1111101010111100; // vC=-1348 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b1111101100100001; // vC=-1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110011; // iC= 1779 
// vC = 14'b1111101100110000; // vC=-1232 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111001; // iC= 1785 
// vC = 14'b1111101011111101; // vC=-1283 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b1111101110011111; // vC=-1121 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111101; // iC= 2045 
// vC = 14'b1111101011111111; // vC=-1281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000011; // iC= 1795 
// vC = 14'b1111101101011111; // vC=-1185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b1111101111010000; // vC=-1072 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b1111101011001001; // vC=-1335 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111110; // iC= 1854 
// vC = 14'b1111101111011001; // vC=-1063 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b1111101110100011; // vC=-1117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001111; // iC= 2063 
// vC = 14'b1111101100111110; // vC=-1218 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110011; // iC= 2099 
// vC = 14'b1111101111100000; // vC=-1056 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011100; // iC= 1884 
// vC = 14'b1111101100010111; // vC=-1257 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001011; // iC= 2123 
// vC = 14'b1111101111100110; // vC=-1050 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b1111101011101100; // vC=-1300 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b1111101100100100; // vC=-1244 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b1111101100011010; // vC=-1254 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010100; // iC= 2068 
// vC = 14'b1111101011111001; // vC=-1287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b1111101110010011; // vC=-1133 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b1111101101110011; // vC=-1165 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b1111101101110111; // vC=-1161 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011100; // iC= 2140 
// vC = 14'b1111101111110110; // vC=-1034 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011111; // iC= 2079 
// vC = 14'b1111101111101111; // vC=-1041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111110000001000; // vC=-1016 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b1111101100111100; // vC=-1220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011100; // iC= 2012 
// vC = 14'b1111110000010101; // vC=-1003 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101100; // iC= 1900 
// vC = 14'b1111101101101101; // vC=-1171 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011100; // iC= 2140 
// vC = 14'b1111101110011011; // vC=-1125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b1111101110101101; // vC=-1107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b1111101110001101; // vC=-1139 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000011; // iC= 2115 
// vC = 14'b1111110010011110; // vC= -866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111100; // iC= 1916 
// vC = 14'b1111110001011111; // vC= -929 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111101111111001; // vC=-1031 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011000; // iC= 2072 
// vC = 14'b1111110000000110; // vC=-1018 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110010; // iC= 2034 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100000; // iC= 2080 
// vC = 14'b1111110010000010; // vC= -894 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111101110100011; // vC=-1117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b1111110000111011; // vC= -965 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110100; // iC= 2164 
// vC = 14'b1111110000100110; // vC= -986 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b1111110000100011; // vC= -989 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101011; // iC= 1963 
// vC = 14'b1111110010001010; // vC= -886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b1111110010101100; // vC= -852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101111; // iC= 2159 
// vC = 14'b1111110001110110; // vC= -906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010011; // iC= 1875 
// vC = 14'b1111110011101111; // vC= -785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b1111110010001000; // vC= -888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100010; // iC= 2146 
// vC = 14'b1111101111100111; // vC=-1049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101110; // iC= 1966 
// vC = 14'b1111110100010111; // vC= -745 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010010; // iC= 2130 
// vC = 14'b1111110000110110; // vC= -970 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b1111110011110000; // vC= -784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111110011011011; // vC= -805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b1111110000010100; // vC=-1004 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b1111110101011010; // vC= -678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b1111110001001111; // vC= -945 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101010; // iC= 2090 
// vC = 14'b1111110011110100; // vC= -780 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b1111110010001111; // vC= -881 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000010; // iC= 1986 
// vC = 14'b1111110010000111; // vC= -889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000101; // iC= 2117 
// vC = 14'b1111110001010000; // vC= -944 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b1111110100111100; // vC= -708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b1111110100010000; // vC= -752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101011; // iC= 1899 
// vC = 14'b1111110101101001; // vC= -663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100101; // iC= 2149 
// vC = 14'b1111110011111111; // vC= -769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b1111110101011111; // vC= -673 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001100; // iC= 2188 
// vC = 14'b1111110010110001; // vC= -847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111110011100000; // vC= -800 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b1111110110110100; // vC= -588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b1111110110100011; // vC= -605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b1111110111011101; // vC= -547 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b1111110100011100; // vC= -740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011111; // iC= 1887 
// vC = 14'b1111110100111010; // vC= -710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100000; // iC= 2144 
// vC = 14'b1111110110000010; // vC= -638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b1111110110010011; // vC= -621 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111110101010110; // vC= -682 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110101; // iC= 2037 
// vC = 14'b1111110100100001; // vC= -735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000010; // iC= 1922 
// vC = 14'b1111110110110001; // vC= -591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011010; // iC= 2074 
// vC = 14'b1111110111011011; // vC= -549 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b1111110101110000; // vC= -656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010101; // iC= 2197 
// vC = 14'b1111110110000010; // vC= -638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000110; // iC= 2182 
// vC = 14'b1111110110000001; // vC= -639 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011111; // iC= 2207 
// vC = 14'b1111110101111010; // vC= -646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b1111110111111111; // vC= -513 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b1111111000110100; // vC= -460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011011; // iC= 2203 
// vC = 14'b1111110101101111; // vC= -657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b1111110101011001; // vC= -679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011110; // iC= 2206 
// vC = 14'b1111110110111110; // vC= -578 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b1111110110101100; // vC= -596 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b1111111000111100; // vC= -452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010101; // iC= 2005 
// vC = 14'b1111111001011110; // vC= -418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100010; // iC= 2146 
// vC = 14'b1111111001001010; // vC= -438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111010; // iC= 1978 
// vC = 14'b1111111000101001; // vC= -471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001001; // iC= 2185 
// vC = 14'b1111111000100010; // vC= -478 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110101; // iC= 2101 
// vC = 14'b1111110110000110; // vC= -634 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101110; // iC= 2158 
// vC = 14'b1111110111111110; // vC= -514 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110011; // iC= 2099 
// vC = 14'b1111110111000101; // vC= -571 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101100; // iC= 2092 
// vC = 14'b1111111010001110; // vC= -370 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000110; // iC= 2118 
// vC = 14'b1111110110110010; // vC= -590 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111100; // iC= 2044 
// vC = 14'b1111111001111111; // vC= -385 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b1111111010000100; // vC= -380 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b1111111001000001; // vC= -447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100011; // iC= 2083 
// vC = 14'b1111110111100111; // vC= -537 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b1111111011101110; // vC= -274 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b1111111100000101; // vC= -251 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b1111111010101101; // vC= -339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110000; // iC= 1904 
// vC = 14'b1111111001101111; // vC= -401 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010011; // iC= 2067 
// vC = 14'b1111111011001001; // vC= -311 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101101; // iC= 1901 
// vC = 14'b1111111011001100; // vC= -308 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011001; // iC= 2137 
// vC = 14'b1111111100000111; // vC= -249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111111001101101; // vC= -403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110000; // iC= 1968 
// vC = 14'b1111111101010100; // vC= -172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010010; // iC= 2194 
// vC = 14'b1111111001001000; // vC= -440 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000011; // iC= 2179 
// vC = 14'b1111111101010000; // vC= -176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b1111111100010011; // vC= -237 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001111; // iC= 2127 
// vC = 14'b1111111100100101; // vC= -219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100111; // iC= 2087 
// vC = 14'b1111111010100010; // vC= -350 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111111010111011; // vC= -325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011100; // iC= 2012 
// vC = 14'b1111111010000010; // vC= -382 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001101; // iC= 2125 
// vC = 14'b1111111001011111; // vC= -417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001110; // iC= 2126 
// vC = 14'b1111111101010110; // vC= -170 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b1111111100100011; // vC= -221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110101; // iC= 2101 
// vC = 14'b1111111011111001; // vC= -263 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100001; // iC= 2081 
// vC = 14'b1111111100011010; // vC= -230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011101; // iC= 1885 
// vC = 14'b1111111010101001; // vC= -343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b1111111100001100; // vC= -244 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b1111111101001111; // vC= -177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000010; // iC= 2050 
// vC = 14'b1111111011010111; // vC= -297 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101101; // iC= 2029 
// vC = 14'b1111111101111101; // vC= -131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000011; // iC= 2115 
// vC = 14'b1111111111101110; // vC=  -18 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b1111111110100010; // vC=  -94 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b1111111100100001; // vC= -223 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000101; // iC= 1989 
// vC = 14'b1111111111110111; // vC=   -9 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111001; // iC= 2105 
// vC = 14'b1111111111011001; // vC=  -39 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001011; // iC= 2123 
// vC = 14'b1111111110111110; // vC=  -66 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001010; // iC= 1866 
// vC = 14'b1111111101110011; // vC= -141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b0000000000010000; // vC=   16 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101111; // iC= 1967 
// vC = 14'b0000000000000010; // vC=    2 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000111; // iC= 2183 
// vC = 14'b1111111110001001; // vC= -119 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b1111111101111110; // vC= -130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b0000000000010001; // vC=   17 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111111100111001; // vC= -199 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111110; // iC= 1982 
// vC = 14'b1111111101010111; // vC= -169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b1111111111100111; // vC=  -25 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110000; // iC= 2096 
// vC = 14'b1111111111111111; // vC=   -1 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111111110010011; // vC= -109 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101111; // iC= 2095 
// vC = 14'b0000000000010011; // vC=   19 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b0000000001010001; // vC=   81 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111011; // iC= 1851 
// vC = 14'b0000000000011100; // vC=   28 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b0000000001000001; // vC=   65 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001001; // iC= 2057 
// vC = 14'b1111111111010011; // vC=  -45 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100111; // iC= 2151 
// vC = 14'b1111111110011111; // vC=  -97 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111000; // iC= 1976 
// vC = 14'b0000000000101100; // vC=   44 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100000; // iC= 2080 
// vC = 14'b0000000010110011; // vC=  179 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110001; // iC= 1905 
// vC = 14'b1111111111001110; // vC=  -50 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110001; // iC= 1841 
// vC = 14'b0000000001101101; // vC=  109 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b0000000001011100; // vC=   92 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b0000000001001000; // vC=   72 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111111111000101; // vC=  -59 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b0000000001001101; // vC=   77 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100001; // iC= 2145 
// vC = 14'b0000000011000010; // vC=  194 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001111; // iC= 2063 
// vC = 14'b0000000000100001; // vC=   33 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b0000000010111010; // vC=  186 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b0000000010001111; // vC=  143 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b0000000000010000; // vC=   16 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b0000000010101111; // vC=  175 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011111; // iC= 2015 
// vC = 14'b0000000100101010; // vC=  298 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101110; // iC= 2030 
// vC = 14'b0000000010000000; // vC=  128 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010001; // iC= 1937 
// vC = 14'b0000000001001000; // vC=   72 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b0000000010000010; // vC=  130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b0000000010001011; // vC=  139 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b0000000100100011; // vC=  291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000011; // iC= 1859 
// vC = 14'b0000000000110001; // vC=   49 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b0000000011111001; // vC=  249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b0000000100011001; // vC=  281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b0000000101010110; // vC=  342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b0000000101000101; // vC=  325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000011; // iC= 2115 
// vC = 14'b0000000101000111; // vC=  327 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000000; // iC= 1984 
// vC = 14'b0000000100000001; // vC=  257 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b0000000101101001; // vC=  361 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011100; // iC= 1820 
// vC = 14'b0000000101010100; // vC=  340 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b0000000110110101; // vC=  437 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111011; // iC= 1787 
// vC = 14'b0000000101001100; // vC=  332 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101100; // iC= 1900 
// vC = 14'b0000000011100011; // vC=  227 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001011; // iC= 1995 
// vC = 14'b0000000101011011; // vC=  347 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b0000000100101011; // vC=  299 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000000; // iC= 1856 
// vC = 14'b0000000101101101; // vC=  365 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000011; // iC= 2051 
// vC = 14'b0000000110100100; // vC=  420 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b0000000110100111; // vC=  423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110111; // iC= 1783 
// vC = 14'b0000000111110100; // vC=  500 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b0000000110101111; // vC=  431 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110100; // iC= 1780 
// vC = 14'b0000000110110010; // vC=  434 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100110; // iC= 2086 
// vC = 14'b0000000111011101; // vC=  477 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100100; // iC= 1892 
// vC = 14'b0000001000001100; // vC=  524 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010110; // iC= 1878 
// vC = 14'b0000000101111101; // vC=  381 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101011; // iC= 1771 
// vC = 14'b0000000110001100; // vC=  396 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010111; // iC= 1879 
// vC = 14'b0000000101110111; // vC=  375 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000000111000101; // vC=  453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000011; // iC= 2051 
// vC = 14'b0000000111011010; // vC=  474 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101011; // iC= 1899 
// vC = 14'b0000000101011011; // vC=  347 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110001; // iC= 1841 
// vC = 14'b0000001001010100; // vC=  596 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b0000000111000100; // vC=  452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b0000000101000000; // vC=  320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000001; // iC= 1921 
// vC = 14'b0000001000011100; // vC=  540 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000010; // iC= 1922 
// vC = 14'b0000000111000010; // vC=  450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b0000000100111110; // vC=  318 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b0000000101111110; // vC=  382 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b0000000111000111; // vC=  455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011110; // iC= 1822 
// vC = 14'b0000000110110011; // vC=  435 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b0000001000101100; // vC=  556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000100; // iC= 1924 
// vC = 14'b0000001001011011; // vC=  603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b0000000101110011; // vC=  371 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011000; // iC= 1880 
// vC = 14'b0000001010100101; // vC=  677 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101101; // iC= 1901 
// vC = 14'b0000001011000111; // vC=  711 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101110; // iC= 2030 
// vC = 14'b0000001010111001; // vC=  697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111100; // iC= 1724 
// vC = 14'b0000001000110110; // vC=  566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001111; // iC= 1743 
// vC = 14'b0000000110111001; // vC=  441 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b0000001000111111; // vC=  575 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b0000001010100110; // vC=  678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b0000000110111011; // vC=  443 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001111; // iC= 1743 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000101; // iC= 1925 
// vC = 14'b0000001001101100; // vC=  620 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110010; // iC= 1714 
// vC = 14'b0000000111010001; // vC=  465 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011001; // iC= 1817 
// vC = 14'b0000000111101001; // vC=  489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110001; // iC= 1713 
// vC = 14'b0000001100000011; // vC=  771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111110; // iC= 1726 
// vC = 14'b0000001100010001; // vC=  785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000001; // iC= 1729 
// vC = 14'b0000001010110111; // vC=  695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b0000001011111011; // vC=  763 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010110; // iC= 1686 
// vC = 14'b0000000111111010; // vC=  506 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110110; // iC= 1718 
// vC = 14'b0000001010111001; // vC=  697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b0000001011000101; // vC=  709 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b0000001000010011; // vC=  531 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010110; // iC= 1878 
// vC = 14'b0000001101010101; // vC=  853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b0000001001100110; // vC=  614 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b0000001011100100; // vC=  740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010001; // iC= 1937 
// vC = 14'b0000001101000101; // vC=  837 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001011; // iC= 1675 
// vC = 14'b0000001001100110; // vC=  614 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001100; // iC= 1740 
// vC = 14'b0000001010111010; // vC=  698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010110; // iC= 1750 
// vC = 14'b0000001001000110; // vC=  582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011011; // iC= 1627 
// vC = 14'b0000001010000100; // vC=  644 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b0000001001100110; // vC=  614 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110111; // iC= 1847 
// vC = 14'b0000001100010001; // vC=  785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100101; // iC= 1765 
// vC = 14'b0000001101010011; // vC=  851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101100; // iC= 1900 
// vC = 14'b0000001011101110; // vC=  750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111111; // iC= 1855 
// vC = 14'b0000001100000000; // vC=  768 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110101; // iC= 1781 
// vC = 14'b0000001001111100; // vC=  636 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010100; // iC= 1684 
// vC = 14'b0000001110100110; // vC=  934 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011001; // iC= 1817 
// vC = 14'b0000001100010000; // vC=  784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011111; // iC= 1759 
// vC = 14'b0000001111010000; // vC=  976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000101; // iC= 1861 
// vC = 14'b0000001011101001; // vC=  745 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111010; // iC= 1786 
// vC = 14'b0000001101001110; // vC=  846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111101; // iC= 1661 
// vC = 14'b0000001010111101; // vC=  701 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001001; // iC= 1737 
// vC = 14'b0000001101001110; // vC=  846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100100; // iC= 1892 
// vC = 14'b0000001011100100; // vC=  740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000110; // iC= 1606 
// vC = 14'b0000001101110001; // vC=  881 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100000; // iC= 1568 
// vC = 14'b0000001110011100; // vC=  924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111100; // iC= 1660 
// vC = 14'b0000001100000110; // vC=  774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010001; // iC= 1745 
// vC = 14'b0000001101011101; // vC=  861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111011; // iC= 1595 
// vC = 14'b0000001100001111; // vC=  783 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001101; // iC= 1741 
// vC = 14'b0000001100001010; // vC=  778 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110001; // iC= 1713 
// vC = 14'b0000001011110001; // vC=  753 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101000; // iC= 1768 
// vC = 14'b0000001111010010; // vC=  978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111101; // iC= 1661 
// vC = 14'b0000001110000000; // vC=  896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b0000001111101110; // vC= 1006 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001111; // iC= 1615 
// vC = 14'b0000001101011100; // vC=  860 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101101; // iC= 1773 
// vC = 14'b0000001101001101; // vC=  845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101110; // iC= 1710 
// vC = 14'b0000001111100010; // vC=  994 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000011; // iC= 1667 
// vC = 14'b0000010001000011; // vC= 1091 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001010; // iC= 1674 
// vC = 14'b0000010000001001; // vC= 1033 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011110; // iC= 1758 
// vC = 14'b0000001110101111; // vC=  943 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110101; // iC= 1589 
// vC = 14'b0000001101001000; // vC=  840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010001; // iC= 1553 
// vC = 14'b0000001111001101; // vC=  973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011110; // iC= 1566 
// vC = 14'b0000001111000110; // vC=  966 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111001; // iC= 1785 
// vC = 14'b0000001110010000; // vC=  912 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001001; // iC= 1609 
// vC = 14'b0000010001100110; // vC= 1126 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101111; // iC= 1647 
// vC = 14'b0000010000000100; // vC= 1028 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011011; // iC= 1627 
// vC = 14'b0000010000111101; // vC= 1085 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100110; // iC= 1510 
// vC = 14'b0000010000111111; // vC= 1087 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011111; // iC= 1695 
// vC = 14'b0000010010001010; // vC= 1162 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010100; // iC= 1492 
// vC = 14'b0000010001101001; // vC= 1129 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110110; // iC= 1590 
// vC = 14'b0000010010101001; // vC= 1193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001110; // iC= 1614 
// vC = 14'b0000001110101001; // vC=  937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101101; // iC= 1773 
// vC = 14'b0000001110010001; // vC=  913 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011101; // iC= 1693 
// vC = 14'b0000001111000111; // vC=  967 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111101; // iC= 1469 
// vC = 14'b0000010010100001; // vC= 1185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101101; // iC= 1773 
// vC = 14'b0000010001111010; // vC= 1146 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110110; // iC= 1462 
// vC = 14'b0000001110111011; // vC=  955 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110010; // iC= 1522 
// vC = 14'b0000010000001011; // vC= 1035 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111000; // iC= 1592 
// vC = 14'b0000010011010111; // vC= 1239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010000; // iC= 1552 
// vC = 14'b0000010011101101; // vC= 1261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000110; // iC= 1606 
// vC = 14'b0000010010100001; // vC= 1185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100101; // iC= 1573 
// vC = 14'b0000010001100111; // vC= 1127 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101010; // iC= 1450 
// vC = 14'b0000001111110000; // vC= 1008 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100000; // iC= 1696 
// vC = 14'b0000001111001111; // vC=  975 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111001; // iC= 1657 
// vC = 14'b0000010010101100; // vC= 1196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011100; // iC= 1500 
// vC = 14'b0000010100011010; // vC= 1306 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010100; // iC= 1492 
// vC = 14'b0000010010111010; // vC= 1210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100111; // iC= 1447 
// vC = 14'b0000010000001111; // vC= 1039 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101011; // iC= 1579 
// vC = 14'b0000010011111100; // vC= 1276 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011111; // iC= 1503 
// vC = 14'b0000010001100010; // vC= 1122 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110011; // iC= 1523 
// vC = 14'b0000010011011100; // vC= 1244 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101101; // iC= 1517 
// vC = 14'b0000010100000100; // vC= 1284 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001000; // iC= 1608 
// vC = 14'b0000010011000110; // vC= 1222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100010; // iC= 1442 
// vC = 14'b0000010011000110; // vC= 1222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000000; // iC= 1536 
// vC = 14'b0000010001111011; // vC= 1147 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111000; // iC= 1592 
// vC = 14'b0000010100001101; // vC= 1293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110011; // iC= 1651 
// vC = 14'b0000010010110101; // vC= 1205 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011001; // iC= 1497 
// vC = 14'b0000010100010011; // vC= 1299 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011101; // iC= 1629 
// vC = 14'b0000010011010101; // vC= 1237 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100001; // iC= 1377 
// vC = 14'b0000010010110100; // vC= 1204 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111110; // iC= 1534 
// vC = 14'b0000010100110001; // vC= 1329 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111011; // iC= 1403 
// vC = 14'b0000010100000001; // vC= 1281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111011; // iC= 1467 
// vC = 14'b0000010001101111; // vC= 1135 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100001; // iC= 1569 
// vC = 14'b0000010011011000; // vC= 1240 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000111; // iC= 1351 
// vC = 14'b0000010010010100; // vC= 1172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111101; // iC= 1597 
// vC = 14'b0000010101101011; // vC= 1387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101010; // iC= 1322 
// vC = 14'b0000010110000011; // vC= 1411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000111; // iC= 1607 
// vC = 14'b0000010100111010; // vC= 1338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101111; // iC= 1391 
// vC = 14'b0000010011011101; // vC= 1245 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001100; // iC= 1356 
// vC = 14'b0000010011110000; // vC= 1264 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111010; // iC= 1466 
// vC = 14'b0000010100110110; // vC= 1334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001100; // iC= 1292 
// vC = 14'b0000010101011101; // vC= 1373 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001010; // iC= 1546 
// vC = 14'b0000010100100011; // vC= 1315 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000101; // iC= 1477 
// vC = 14'b0000010010000110; // vC= 1158 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100001; // iC= 1441 
// vC = 14'b0000010100000101; // vC= 1285 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110100; // iC= 1524 
// vC = 14'b0000010110010011; // vC= 1427 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111110; // iC= 1278 
// vC = 14'b0000010100001101; // vC= 1293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001101; // iC= 1357 
// vC = 14'b0000010111011100; // vC= 1500 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010000; // iC= 1552 
// vC = 14'b0000010010110010; // vC= 1202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110010; // iC= 1266 
// vC = 14'b0000010010101100; // vC= 1196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010011; // iC= 1427 
// vC = 14'b0000010100000111; // vC= 1287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000110; // iC= 1286 
// vC = 14'b0000010110111001; // vC= 1465 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001100; // iC= 1420 
// vC = 14'b0000010110111101; // vC= 1469 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010001; // iC= 1425 
// vC = 14'b0000010100000101; // vC= 1285 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010000; // iC= 1424 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101101; // iC= 1261 
// vC = 14'b0000010110000111; // vC= 1415 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101101; // iC= 1261 
// vC = 14'b0000011000001010; // vC= 1546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000110; // iC= 1478 
// vC = 14'b0000010111111011; // vC= 1531 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101011; // iC= 1259 
// vC = 14'b0000010101011101; // vC= 1373 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100101; // iC= 1445 
// vC = 14'b0000010111000011; // vC= 1475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010001; // iC= 1233 
// vC = 14'b0000011000010100; // vC= 1556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000000; // iC= 1216 
// vC = 14'b0000010110111000; // vC= 1464 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000001; // iC= 1281 
// vC = 14'b0000011000110010; // vC= 1586 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110110; // iC= 1270 
// vC = 14'b0000010111110011; // vC= 1523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011001; // iC= 1241 
// vC = 14'b0000010111000101; // vC= 1477 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100011; // iC= 1187 
// vC = 14'b0000011000000110; // vC= 1542 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001010; // iC= 1354 
// vC = 14'b0000010110110011; // vC= 1459 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101110; // iC= 1198 
// vC = 14'b0000010100110000; // vC= 1328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001011; // iC= 1227 
// vC = 14'b0000010101101000; // vC= 1384 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111100; // iC= 1212 
// vC = 14'b0000010110001110; // vC= 1422 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111101; // iC= 1149 
// vC = 14'b0000010110010110; // vC= 1430 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100101; // iC= 1253 
// vC = 14'b0000010110100110; // vC= 1446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110101; // iC= 1141 
// vC = 14'b0000010101010010; // vC= 1362 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010110; // iC= 1238 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101101; // iC= 1325 
// vC = 14'b0000010101011010; // vC= 1370 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100000; // iC= 1184 
// vC = 14'b0000011000101011; // vC= 1579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101001; // iC= 1193 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111100; // iC= 1148 
// vC = 14'b0000011000110101; // vC= 1589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010001; // iC= 1169 
// vC = 14'b0000011000010000; // vC= 1552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110011; // iC= 1331 
// vC = 14'b0000011001001000; // vC= 1608 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001110; // iC= 1230 
// vC = 14'b0000010111000100; // vC= 1476 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110101; // iC= 1077 
// vC = 14'b0000011010001000; // vC= 1672 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000110; // iC= 1222 
// vC = 14'b0000010101111110; // vC= 1406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110011; // iC= 1331 
// vC = 14'b0000011001011010; // vC= 1626 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101000; // iC= 1128 
// vC = 14'b0000011010101100; // vC= 1708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111010; // iC= 1210 
// vC = 14'b0000011010011100; // vC= 1692 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101001; // iC= 1257 
// vC = 14'b0000011001101011; // vC= 1643 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001100; // iC= 1356 
// vC = 14'b0000011010001101; // vC= 1677 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100110; // iC= 1318 
// vC = 14'b0000010110101000; // vC= 1448 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100011; // iC= 1123 
// vC = 14'b0000010111111110; // vC= 1534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100101; // iC= 1061 
// vC = 14'b0000011011001010; // vC= 1738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100011; // iC= 1059 
// vC = 14'b0000011000100111; // vC= 1575 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000101; // iC= 1093 
// vC = 14'b0000011010000011; // vC= 1667 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111101; // iC= 1085 
// vC = 14'b0000011010000000; // vC= 1664 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010101; // iC= 1237 
// vC = 14'b0000011001011100; // vC= 1628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011111; // iC= 1247 
// vC = 14'b0000010110110000; // vC= 1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101011; // iC= 1067 
// vC = 14'b0000010111111100; // vC= 1532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000111; // iC= 1287 
// vC = 14'b0000010110101101; // vC= 1453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000111; // iC= 1159 
// vC = 14'b0000011000011010; // vC= 1562 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000101; // iC= 1029 
// vC = 14'b0000011011010000; // vC= 1744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000011; // iC= 1091 
// vC = 14'b0000011000110111; // vC= 1591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111000; // iC= 1208 
// vC = 14'b0000011010101000; // vC= 1704 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001000; // iC= 1096 
// vC = 14'b0000011000011101; // vC= 1565 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000101; // iC=  965 
// vC = 14'b0000011001010001; // vC= 1617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101110; // iC= 1006 
// vC = 14'b0000011001110010; // vC= 1650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010101; // iC=  981 
// vC = 14'b0000011010011110; // vC= 1694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100000; // iC= 1056 
// vC = 14'b0000010111011011; // vC= 1499 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101100; // iC= 1132 
// vC = 14'b0000011000110011; // vC= 1587 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001010; // iC= 1098 
// vC = 14'b0000011100000110; // vC= 1798 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010100; // iC= 1172 
// vC = 14'b0000011001011000; // vC= 1624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101000; // iC= 1192 
// vC = 14'b0000011001110111; // vC= 1655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000110; // iC= 1158 
// vC = 14'b0000011001010100; // vC= 1620 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001011; // iC=  971 
// vC = 14'b0000011000101110; // vC= 1582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100010; // iC= 1186 
// vC = 14'b0000011000010110; // vC= 1558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000110; // iC= 1158 
// vC = 14'b0000011000110001; // vC= 1585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111110; // iC= 1150 
// vC = 14'b0000011100011000; // vC= 1816 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011001; // iC=  921 
// vC = 14'b0000011001000011; // vC= 1603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001111; // iC=  975 
// vC = 14'b0000011001101001; // vC= 1641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111011; // iC=  955 
// vC = 14'b0000011010110111; // vC= 1719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010000; // iC= 1040 
// vC = 14'b0000011010101001; // vC= 1705 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111110; // iC= 1150 
// vC = 14'b0000011100011101; // vC= 1821 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100111; // iC= 1063 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100000; // iC= 1056 
// vC = 14'b0000011001000011; // vC= 1603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011110; // iC=  990 
// vC = 14'b0000011011100011; // vC= 1763 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100011; // iC= 1059 
// vC = 14'b0000011000100101; // vC= 1573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001101; // iC=  973 
// vC = 14'b0000011100001010; // vC= 1802 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110111; // iC= 1079 
// vC = 14'b0000011010010010; // vC= 1682 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011110; // iC= 1054 
// vC = 14'b0000011001010000; // vC= 1616 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011001; // iC= 1049 
// vC = 14'b0000011010111010; // vC= 1722 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011110; // iC=  926 
// vC = 14'b0000011010000101; // vC= 1669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001010; // iC= 1098 
// vC = 14'b0000011100011111; // vC= 1823 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010101; // iC=  917 
// vC = 14'b0000011000111110; // vC= 1598 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001011; // iC=  843 
// vC = 14'b0000011100011001; // vC= 1817 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111100; // iC= 1084 
// vC = 14'b0000011011000111; // vC= 1735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011101; // iC=  989 
// vC = 14'b0000011011011100; // vC= 1756 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100001; // iC=  929 
// vC = 14'b0000011100110011; // vC= 1843 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110001; // iC=  817 
// vC = 14'b0000011011010010; // vC= 1746 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100100; // iC=  868 
// vC = 14'b0000011001010010; // vC= 1618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000100; // iC=  900 
// vC = 14'b0000011100011110; // vC= 1822 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011101; // iC= 1053 
// vC = 14'b0000011010110010; // vC= 1714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100000; // iC=  992 
// vC = 14'b0000011110010100; // vC= 1940 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000110; // iC=  838 
// vC = 14'b0000011011101010; // vC= 1770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110001; // iC= 1009 
// vC = 14'b0000011100011000; // vC= 1816 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000011; // iC= 1027 
// vC = 14'b0000011101011110; // vC= 1886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101111; // iC=  943 
// vC = 14'b0000011100100111; // vC= 1831 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000100; // iC=  964 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010011; // iC=  723 
// vC = 14'b0000011110100001; // vC= 1953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101010; // iC=  810 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001001; // iC=  969 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010011; // iC=  851 
// vC = 14'b0000011101011010; // vC= 1882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011101; // iC=  989 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101011; // iC=  811 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100011; // iC=  931 
// vC = 14'b0000011110011101; // vC= 1949 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111011; // iC=  827 
// vC = 14'b0000011110011010; // vC= 1946 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111100; // iC=  892 
// vC = 14'b0000011101011110; // vC= 1886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111111; // iC=  959 
// vC = 14'b0000011110111100; // vC= 1980 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011000; // iC=  728 
// vC = 14'b0000011110101001; // vC= 1961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111011; // iC=  763 
// vC = 14'b0000011011010110; // vC= 1750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011010; // iC=  858 
// vC = 14'b0000011110011100; // vC= 1948 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000000; // iC=  768 
// vC = 14'b0000011011011111; // vC= 1759 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111011; // iC=  763 
// vC = 14'b0000011110010111; // vC= 1943 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100000; // iC=  672 
// vC = 14'b0000011010111100; // vC= 1724 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000111; // iC=  647 
// vC = 14'b0000011011110101; // vC= 1781 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100001; // iC=  737 
// vC = 14'b0000011110000001; // vC= 1921 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100110; // iC=  870 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110000; // iC=  880 
// vC = 14'b0000011110110110; // vC= 1974 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b0000011011000011; // vC= 1731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010000; // iC=  720 
// vC = 14'b0000011111011000; // vC= 2008 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111100; // iC=  636 
// vC = 14'b0000011101110000; // vC= 1904 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001110; // iC=  718 
// vC = 14'b0000011101111011; // vC= 1915 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010000; // iC=  720 
// vC = 14'b0000011100101001; // vC= 1833 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000010; // iC=  578 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111100; // iC=  764 
// vC = 14'b0000011111100011; // vC= 2019 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111100; // iC=  572 
// vC = 14'b0000011111110100; // vC= 2036 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110001; // iC=  561 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101100; // iC=  748 
// vC = 14'b0000011100011011; // vC= 1819 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000101; // iC=  709 
// vC = 14'b0000011011110001; // vC= 1777 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010101; // iC=  789 
// vC = 14'b0000011111100011; // vC= 2019 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000100; // iC=  516 
// vC = 14'b0000100000001001; // vC= 2057 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011001; // iC=  729 
// vC = 14'b0000011111111111; // vC= 2047 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010110; // iC=  662 
// vC = 14'b0000011110000000; // vC= 1920 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000000; // iC=  768 
// vC = 14'b0000011110111000; // vC= 1976 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011100; // iC=  476 
// vC = 14'b0000011101100100; // vC= 1892 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111101; // iC=  637 
// vC = 14'b0000011110110010; // vC= 1970 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011110; // iC=  606 
// vC = 14'b0000011101101001; // vC= 1897 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000100; // iC=  772 
// vC = 14'b0000011110011001; // vC= 1945 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001001; // iC=  585 
// vC = 14'b0000100000010001; // vC= 2065 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100101; // iC=  549 
// vC = 14'b0000011101100010; // vC= 1890 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010000; // iC=  592 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001101; // iC=  525 
// vC = 14'b0000011100101011; // vC= 1835 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101011; // iC=  555 
// vC = 14'b0000100000011001; // vC= 2073 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011011; // iC=  411 
// vC = 14'b0000011111100000; // vC= 2016 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010110; // iC=  534 
// vC = 14'b0000011110101010; // vC= 1962 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001111; // iC=  527 
// vC = 14'b0000011111000010; // vC= 1986 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001011; // iC=  651 
// vC = 14'b0000011011101111; // vC= 1775 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010011; // iC=  595 
// vC = 14'b0000011110001001; // vC= 1929 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110111; // iC=  567 
// vC = 14'b0000011101011110; // vC= 1886 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011011; // iC=  603 
// vC = 14'b0000011101101000; // vC= 1896 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010000; // iC=  400 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010101; // iC=  469 
// vC = 14'b0000011100111001; // vC= 1849 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000100; // iC=  388 
// vC = 14'b0000011110000000; // vC= 1920 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110100; // iC=  308 
// vC = 14'b0000100000110011; // vC= 2099 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000100; // iC=  324 
// vC = 14'b0000100000000111; // vC= 2055 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000100; // iC=  388 
// vC = 14'b0000011110001100; // vC= 1932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111111; // iC=  383 
// vC = 14'b0000011110000100; // vC= 1924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000011; // iC=  323 
// vC = 14'b0000011101110000; // vC= 1904 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011010; // iC=  282 
// vC = 14'b0000011111101111; // vC= 2031 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111101; // iC=  445 
// vC = 14'b0000100000101000; // vC= 2088 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011101; // iC=  285 
// vC = 14'b0000011110111000; // vC= 1976 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001010; // iC=  202 
// vC = 14'b0000011110101001; // vC= 1961 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111000; // iC=  184 
// vC = 14'b0000011111100111; // vC= 2023 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100101; // iC=  293 
// vC = 14'b0000100000000000; // vC= 2048 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010011; // iC=  211 
// vC = 14'b0000011110110111; // vC= 1975 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000011; // iC=  259 
// vC = 14'b0000011101110101; // vC= 1909 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011000; // iC=   88 
// vC = 14'b0000100000101101; // vC= 2093 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000101; // iC=  325 
// vC = 14'b0000011111100101; // vC= 2021 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011100; // iC=  284 
// vC = 14'b0000100000101110; // vC= 2094 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001110; // iC=  206 
// vC = 14'b0000011111101110; // vC= 2030 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110001; // iC=  113 
// vC = 14'b0000011100010001; // vC= 1809 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100010; // iC=  162 
// vC = 14'b0000011110000011; // vC= 1923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100000; // iC=   96 
// vC = 14'b0000011100101100; // vC= 1836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110011; // iC=  243 
// vC = 14'b0000011101111010; // vC= 1914 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001000111; // iC=   71 
// vC = 14'b0000011101111010; // vC= 1914 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010101; // iC=   85 
// vC = 14'b0000100001001100; // vC= 2124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111111; // iC=  191 
// vC = 14'b0000011100001101; // vC= 1805 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101011; // iC=  107 
// vC = 14'b0000011111111110; // vC= 2046 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010000; // iC= -112 
// vC = 14'b0000011110111011; // vC= 1979 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010010; // iC= -174 
// vC = 14'b0000011100011110; // vC= 1822 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100011; // iC=   35 
// vC = 14'b0000100000000110; // vC= 2054 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011010; // iC=   90 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100011; // iC= -157 
// vC = 14'b0000011101111010; // vC= 1914 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101001; // iC=   41 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111101; // iC= -131 
// vC = 14'b0000100000110001; // vC= 2097 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100100; // iC= -220 
// vC = 14'b0000011110010011; // vC= 1939 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100001; // iC=  -95 
// vC = 14'b0000011101010011; // vC= 1875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010010; // iC= -302 
// vC = 14'b0000011100000101; // vC= 1797 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001110; // iC= -242 
// vC = 14'b0000011100011010; // vC= 1818 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011100010; // iC= -286 
// vC = 14'b0000011101000001; // vC= 1857 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011011; // iC= -357 
// vC = 14'b0000011111101000; // vC= 2024 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011100; // iC= -356 
// vC = 14'b0000011111010010; // vC= 2002 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110001; // iC= -335 
// vC = 14'b0000100000110101; // vC= 2101 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110100; // iC= -204 
// vC = 14'b0000100000010000; // vC= 2064 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011100101; // iC= -283 
// vC = 14'b0000011100110010; // vC= 1842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101101; // iC= -403 
// vC = 14'b0000011111101010; // vC= 2026 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010111; // iC= -425 
// vC = 14'b0000100000101100; // vC= 2092 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000011; // iC= -573 
// vC = 14'b0000011111111000; // vC= 2040 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101010; // iC= -470 
// vC = 14'b0000011110011001; // vC= 1945 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101101; // iC= -467 
// vC = 14'b0000011100110100; // vC= 1844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101110; // iC= -466 
// vC = 14'b0000011111000111; // vC= 1991 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000111; // iC= -377 
// vC = 14'b0000011110011100; // vC= 1948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101001; // iC= -535 
// vC = 14'b0000011101010001; // vC= 1873 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000100; // iC= -636 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010010; // iC= -750 
// vC = 14'b0000011110101010; // vC= 1962 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000000101; // iC= -507 
// vC = 14'b0000011110011101; // vC= 1949 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011011; // iC= -741 
// vC = 14'b0000100000010001; // vC= 2065 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000010; // iC= -574 
// vC = 14'b0000011100111100; // vC= 1852 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010110; // iC= -618 
// vC = 14'b0000011111110100; // vC= 2036 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111111; // iC= -769 
// vC = 14'b0000011011011101; // vC= 1757 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111000; // iC= -712 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110000; // iC= -784 
// vC = 14'b0000011011001101; // vC= 1741 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101110; // iC= -658 
// vC = 14'b0000011110110100; // vC= 1972 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110010; // iC= -846 
// vC = 14'b0000011101000101; // vC= 1861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110101; // iC= -971 
// vC = 14'b0000011101101010; // vC= 1898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101001; // iC= -919 
// vC = 14'b0000011100001100; // vC= 1804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101001; // iC= -727 
// vC = 14'b0000011101010010; // vC= 1874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101100; // iC= -980 
// vC = 14'b0000011101101100; // vC= 1900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010001; // iC= -751 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101101; // iC=-1043 
// vC = 14'b0000011110001110; // vC= 1934 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100100; // iC=-1052 
// vC = 14'b0000011110101101; // vC= 1965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001101; // iC= -947 
// vC = 14'b0000011111010001; // vC= 2001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100000; // iC=-1120 
// vC = 14'b0000011010101001; // vC= 1705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001111; // iC= -881 
// vC = 14'b0000011110100001; // vC= 1953 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010010; // iC= -942 
// vC = 14'b0000011110100011; // vC= 1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101100; // iC=-1108 
// vC = 14'b0000011111010001; // vC= 2001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000101; // iC=-1083 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110000; // iC=-1168 
// vC = 14'b0000011010110001; // vC= 1713 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111101; // iC=-1091 
// vC = 14'b0000011100101111; // vC= 1839 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110110; // iC=-1098 
// vC = 14'b0000011010010101; // vC= 1685 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101000; // iC=-1048 
// vC = 14'b0000011110110110; // vC= 1974 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101001; // iC=-1047 
// vC = 14'b0000011101101010; // vC= 1898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110001; // iC=-1039 
// vC = 14'b0000011011011100; // vC= 1756 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001001; // iC=-1335 
// vC = 14'b0000011100010110; // vC= 1814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010001; // iC=-1263 
// vC = 14'b0000011100110011; // vC= 1843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110001; // iC=-1167 
// vC = 14'b0000011010111000; // vC= 1720 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111001; // iC=-1159 
// vC = 14'b0000011010010111; // vC= 1687 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001111; // iC=-1201 
// vC = 14'b0000011010111011; // vC= 1723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101101; // iC=-1363 
// vC = 14'b0000011011000010; // vC= 1730 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001111; // iC=-1329 
// vC = 14'b0000011100111011; // vC= 1851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010110; // iC=-1194 
// vC = 14'b0000011001100000; // vC= 1632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110101; // iC=-1291 
// vC = 14'b0000011011110100; // vC= 1780 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110010; // iC=-1358 
// vC = 14'b0000011001110001; // vC= 1649 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110100; // iC=-1548 
// vC = 14'b0000011100100010; // vC= 1826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100110; // iC=-1370 
// vC = 14'b0000011010100000; // vC= 1696 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010011; // iC=-1453 
// vC = 14'b0000011100001001; // vC= 1801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010110; // iC=-1450 
// vC = 14'b0000011011011001; // vC= 1753 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111111; // iC=-1473 
// vC = 14'b0000011001111010; // vC= 1658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100011; // iC=-1373 
// vC = 14'b0000011100101000; // vC= 1832 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100011; // iC=-1437 
// vC = 14'b0000011100111110; // vC= 1854 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011000; // iC=-1576 
// vC = 14'b0000011100000000; // vC= 1792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101010; // iC=-1622 
// vC = 14'b0000011011101001; // vC= 1769 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011101; // iC=-1635 
// vC = 14'b0000011000101010; // vC= 1578 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011101; // iC=-1699 
// vC = 14'b0000011001011001; // vC= 1625 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011110; // iC=-1634 
// vC = 14'b0000011000100111; // vC= 1575 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000000; // iC=-1472 
// vC = 14'b0000011001010001; // vC= 1617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100000; // iC=-1504 
// vC = 14'b0000010111100001; // vC= 1505 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010110; // iC=-1642 
// vC = 14'b0000010111111101; // vC= 1533 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100010; // iC=-1566 
// vC = 14'b0000011000111000; // vC= 1592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010100; // iC=-1516 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000111; // iC=-1785 
// vC = 14'b0000011011110111; // vC= 1783 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b0000011011000101; // vC= 1733 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100011; // iC=-1757 
// vC = 14'b0000011011011111; // vC= 1759 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111110; // iC=-1666 
// vC = 14'b0000011000001001; // vC= 1545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001011; // iC=-1717 
// vC = 14'b0000010111000001; // vC= 1473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011100; // iC=-1636 
// vC = 14'b0000011010001111; // vC= 1679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b0000011010100100; // vC= 1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101011; // iC=-1685 
// vC = 14'b0000011000111011; // vC= 1595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100101; // iC=-1691 
// vC = 14'b0000010111101100; // vC= 1516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100111; // iC=-1689 
// vC = 14'b0000010110000000; // vC= 1408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111011; // iC=-1733 
// vC = 14'b0000011000011011; // vC= 1563 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b0000010111110000; // vC= 1520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b0000010110100010; // vC= 1442 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100010; // iC=-1630 
// vC = 14'b0000010110100111; // vC= 1447 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001110; // iC=-1778 
// vC = 14'b0000011000110111; // vC= 1591 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000010110111111; // vC= 1471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000101; // iC=-1659 
// vC = 14'b0000011001010000; // vC= 1616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010111; // iC=-1961 
// vC = 14'b0000010110000000; // vC= 1408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000101; // iC=-1915 
// vC = 14'b0000010111101001; // vC= 1513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b0000011001100010; // vC= 1634 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000011000001010; // vC= 1546 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110010; // iC=-1806 
// vC = 14'b0000010101000001; // vC= 1345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b0000010101001111; // vC= 1359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110010; // iC=-1870 
// vC = 14'b0000010100011111; // vC= 1311 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100110; // iC=-1818 
// vC = 14'b0000011000011011; // vC= 1563 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001100; // iC=-1908 
// vC = 14'b0000010111000011; // vC= 1475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100110; // iC=-1754 
// vC = 14'b0000010111000001; // vC= 1473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000011; // iC=-1789 
// vC = 14'b0000010101011011; // vC= 1371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000010; // iC=-1854 
// vC = 14'b0000010110001011; // vC= 1419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b0000010101011110; // vC= 1374 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001001; // iC=-1847 
// vC = 14'b0000010011011100; // vC= 1244 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101101; // iC=-2067 
// vC = 14'b0000010011001111; // vC= 1231 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110111; // iC=-1865 
// vC = 14'b0000010101011111; // vC= 1375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110000; // iC=-1872 
// vC = 14'b0000010101111001; // vC= 1401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010111; // iC=-1833 
// vC = 14'b0000010111000110; // vC= 1478 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011110; // iC=-2018 
// vC = 14'b0000010101011011; // vC= 1371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b0000010101010011; // vC= 1363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b0000010011010000; // vC= 1232 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011101; // iC=-2083 
// vC = 14'b0000010011101000; // vC= 1256 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010111; // iC=-2089 
// vC = 14'b0000010100011000; // vC= 1304 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101010; // iC=-1814 
// vC = 14'b0000010101010001; // vC= 1361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100001; // iC=-1887 
// vC = 14'b0000010010001011; // vC= 1163 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b0000010001110110; // vC= 1142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b0000010100110000; // vC= 1328 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000010100100111; // vC= 1319 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001010; // iC=-1910 
// vC = 14'b0000010101101100; // vC= 1388 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b0000010010100101; // vC= 1189 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011011; // iC=-1829 
// vC = 14'b0000010011101101; // vC= 1261 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000010; // iC=-1918 
// vC = 14'b0000010010010011; // vC= 1171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100000; // iC=-1824 
// vC = 14'b0000010011111101; // vC= 1277 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101001; // iC=-2135 
// vC = 14'b0000010010101001; // vC= 1193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b0000010100010110; // vC= 1302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000110; // iC=-2106 
// vC = 14'b0000010100010111; // vC= 1303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100111; // iC=-2009 
// vC = 14'b0000010001010111; // vC= 1111 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101000; // iC=-1880 
// vC = 14'b0000010001001100; // vC= 1100 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b0000010010011001; // vC= 1177 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111111; // iC=-2049 
// vC = 14'b0000010100100011; // vC= 1315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b0000010011110101; // vC= 1269 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010111; // iC=-1961 
// vC = 14'b0000010011110110; // vC= 1270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000010011011011; // vC= 1243 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000111; // iC=-1977 
// vC = 14'b0000001110111110; // vC=  958 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b0000010011001111; // vC= 1231 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011010; // iC=-2022 
// vC = 14'b0000001111000011; // vC=  963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011010; // iC=-2022 
// vC = 14'b0000010011100000; // vC= 1248 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000001; // iC=-1919 
// vC = 14'b0000010010110000; // vC= 1200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011100; // iC=-1956 
// vC = 14'b0000010001000111; // vC= 1095 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000010001101110; // vC= 1134 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b0000001110100101; // vC=  933 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000001110110001; // vC=  945 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100001; // iC=-2143 
// vC = 14'b0000010001000111; // vC= 1095 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b0000010010001000; // vC= 1160 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b0000001110110101; // vC=  949 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100101; // iC=-2011 
// vC = 14'b0000010000111001; // vC= 1081 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101100; // iC=-2068 
// vC = 14'b0000001110101110; // vC=  942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111001; // iC=-2119 
// vC = 14'b0000010000011100; // vC= 1052 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001111; // iC=-2097 
// vC = 14'b0000010000111111; // vC= 1087 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b0000010001110010; // vC= 1138 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101010; // iC=-2070 
// vC = 14'b0000001101100001; // vC=  865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b0000001101111011; // vC=  891 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b0000001111100100; // vC=  996 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000001111101110; // vC= 1006 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b0000001100101010; // vC=  810 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010111; // iC=-2025 
// vC = 14'b0000001111101010; // vC= 1002 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000001100000110; // vC=  774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110001; // iC=-1935 
// vC = 14'b0000001110100010; // vC=  930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000001101001011; // vC=  843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101100; // iC=-2068 
// vC = 14'b0000001110001011; // vC=  907 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110010; // iC=-1998 
// vC = 14'b0000001110101100; // vC=  940 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101010; // iC=-2070 
// vC = 14'b0000001111101001; // vC= 1001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111000; // iC=-2056 
// vC = 14'b0000001111111001; // vC= 1017 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b0000001101101010; // vC=  874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b0000001010111000; // vC=  696 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b0000001011000000; // vC=  704 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000110; // iC=-2170 
// vC = 14'b0000001110000101; // vC=  901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111110; // iC=-2178 
// vC = 14'b0000001110011100; // vC=  924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011010; // iC=-1894 
// vC = 14'b0000001010010010; // vC=  658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111111; // iC=-2177 
// vC = 14'b0000001100011100; // vC=  796 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b0000001101010001; // vC=  849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011101; // iC=-2083 
// vC = 14'b0000001100101010; // vC=  810 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110010; // iC=-1998 
// vC = 14'b0000001101101011; // vC=  875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110111; // iC=-2121 
// vC = 14'b0000001010100011; // vC=  675 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b0000001001100001; // vC=  609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011000; // iC=-2152 
// vC = 14'b0000001010111111; // vC=  703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b0000001010010010; // vC=  658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000110; // iC=-2170 
// vC = 14'b0000001100110011; // vC=  819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011111; // iC=-2209 
// vC = 14'b0000001100001110; // vC=  782 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001110; // iC=-2226 
// vC = 14'b0000001001011000; // vC=  600 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b0000001010010101; // vC=  661 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010001; // iC=-2159 
// vC = 14'b0000001100100010; // vC=  802 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110010; // iC=-2190 
// vC = 14'b0000001001111010; // vC=  634 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010100; // iC=-2092 
// vC = 14'b0000001011101010; // vC=  746 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b0000000111111010; // vC=  506 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b0000001100010010; // vC=  786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000001000111111; // vC=  575 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b0000001010100110; // vC=  678 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110010; // iC=-1998 
// vC = 14'b0000000111110101; // vC=  501 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b0000001011111011; // vC=  763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000001000001000; // vC=  520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000101; // iC=-2171 
// vC = 14'b0000001001100011; // vC=  611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b0000000111001110; // vC=  462 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111011; // iC=-2117 
// vC = 14'b0000001000110111; // vC=  567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010110; // iC=-2026 
// vC = 14'b0000000110011000; // vC=  408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b0000001011000100; // vC=  708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b0000001011000111; // vC=  711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b0000001001101100; // vC=  620 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000010; // iC=-2174 
// vC = 14'b0000001010000010; // vC=  642 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111110; // iC=-1922 
// vC = 14'b0000001001000011; // vC=  579 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b0000001001000111; // vC=  583 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011000; // iC=-2216 
// vC = 14'b0000001001101101; // vC=  621 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b0000000101111111; // vC=  383 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100011; // iC=-1949 
// vC = 14'b0000001001111000; // vC=  632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111111; // iC=-2049 
// vC = 14'b0000000101000011; // vC=  323 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010111; // iC=-2089 
// vC = 14'b0000001001110000; // vC=  624 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b0000001000100000; // vC=  544 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101011; // iC=-2197 
// vC = 14'b0000000110101101; // vC=  429 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b0000000111111000; // vC=  504 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010101; // iC=-2027 
// vC = 14'b0000000101001110; // vC=  334 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001111; // iC=-2161 
// vC = 14'b0000000100011100; // vC=  284 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b0000000101011001; // vC=  345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101001; // iC=-2135 
// vC = 14'b0000000100001010; // vC=  266 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011000; // iC=-2024 
// vC = 14'b0000000110011101; // vC=  413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010111; // iC=-2089 
// vC = 14'b0000001000000001; // vC=  513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100111; // iC=-2009 
// vC = 14'b0000000100010001; // vC=  273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000000011011110; // vC=  222 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000000111000110; // vC=  454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000100; // iC=-2172 
// vC = 14'b0000000101100101; // vC=  357 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b0000000110010110; // vC=  406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000000111011100; // vC=  476 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000000100010110; // vC=  278 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010101; // iC=-2155 
// vC = 14'b0000000111010110; // vC=  470 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000101; // iC=-2107 
// vC = 14'b0000000110011101; // vC=  413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b0000000101111011; // vC=  379 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000110; // iC=-2106 
// vC = 14'b0000000011110000; // vC=  240 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001110; // iC=-1906 
// vC = 14'b0000000011110000; // vC=  240 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100101; // iC=-2075 
// vC = 14'b0000000101001101; // vC=  333 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110100; // iC=-2124 
// vC = 14'b0000000101001010; // vC=  330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b0000000101101111; // vC=  367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b0000000100110111; // vC=  311 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111110; // iC=-1922 
// vC = 14'b0000000100111011; // vC=  315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010100; // iC=-2092 
// vC = 14'b0000000101101000; // vC=  360 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110111; // iC=-2121 
// vC = 14'b0000000011000101; // vC=  197 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000000011000011; // vC=  195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b0000000100111001; // vC=  313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110100; // iC=-2124 
// vC = 14'b0000000001010000; // vC=   80 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010000; // iC=-2096 
// vC = 14'b0000000100110101; // vC=  309 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011100; // iC=-2148 
// vC = 14'b0000000011001000; // vC=  200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110111; // iC=-2121 
// vC = 14'b0000000100011001; // vC=  281 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001011; // iC=-2165 
// vC = 14'b1111111111110011; // vC=  -13 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b0000000011100111; // vC=  231 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b1111111111110100; // vC=  -12 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000000000111111; // vC=   63 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000000100010001; // vC=  273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110111; // iC=-2185 
// vC = 14'b0000000000010010; // vC=   18 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000000; // iC=-2176 
// vC = 14'b0000000011110110; // vC=  246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b1111111111100001; // vC=  -31 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001011; // iC=-2165 
// vC = 14'b0000000001100010; // vC=   98 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000000000111111; // vC=   63 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110100; // iC=-2188 
// vC = 14'b1111111110110010; // vC=  -78 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b0000000000001011; // vC=   11 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111110; // iC=-2050 
// vC = 14'b0000000010001010; // vC=  138 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b0000000010100101; // vC=  165 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000000000111111; // vC=   63 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b1111111101111110; // vC= -130 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b0000000000100111; // vC=   39 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000000000110011; // vC=   51 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011110; // iC=-2146 
// vC = 14'b1111111110101111; // vC=  -81 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011001; // iC=-2151 
// vC = 14'b1111111111010100; // vC=  -44 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b1111111101010110; // vC= -170 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100000; // iC=-2016 
// vC = 14'b1111111101011110; // vC= -162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b1111111110101001; // vC=  -87 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b1111111110000100; // vC= -124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111100; // iC=-2180 
// vC = 14'b1111111101010111; // vC= -169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b1111111100110000; // vC= -208 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b1111111111001110; // vC=  -50 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b0000000000101110; // vC=   46 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000111; // iC=-2105 
// vC = 14'b1111111100010101; // vC= -235 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011011; // iC=-2085 
// vC = 14'b1111111111000100; // vC=  -60 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b1111111110100001; // vC=  -95 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b1111111011110100; // vC= -268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001111; // iC=-1905 
// vC = 14'b1111111011011111; // vC= -289 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b1111111011101000; // vC= -280 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b1111111111000001; // vC=  -63 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b1111111100101011; // vC= -213 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110010; // iC=-2062 
// vC = 14'b1111111101010011; // vC= -173 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b1111111100110101; // vC= -203 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b1111111100100010; // vC= -222 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b1111111101101001; // vC= -151 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b1111111010101011; // vC= -341 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b1111111010100110; // vC= -346 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b1111111101000111; // vC= -185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101001; // iC=-1879 
// vC = 14'b1111111100001010; // vC= -246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100000; // iC=-1824 
// vC = 14'b1111111011111111; // vC= -257 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b1111111100100101; // vC= -219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111111100010011; // vC= -237 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b1111111101001110; // vC= -178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b1111111010010001; // vC= -367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b1111111010100111; // vC= -345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b1111111011000100; // vC= -316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110010; // iC=-1806 
// vC = 14'b1111111101110111; // vC= -137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b1111111101010011; // vC= -173 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b1111111001100000; // vC= -416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011010; // iC=-2022 
// vC = 14'b1111111000101010; // vC= -470 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111101; // iC=-1859 
// vC = 14'b1111111010001000; // vC= -376 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b1111111100100001; // vC= -223 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000100; // iC=-1980 
// vC = 14'b1111111101000100; // vC= -188 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b1111111001010000; // vC= -432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100101; // iC=-1819 
// vC = 14'b1111111100001001; // vC= -247 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b1111110111110000; // vC= -528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011110; // iC=-1826 
// vC = 14'b1111111001011010; // vC= -422 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010011; // iC=-2093 
// vC = 14'b1111111001000100; // vC= -444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101001; // iC=-2007 
// vC = 14'b1111111010010010; // vC= -366 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011110; // iC=-2082 
// vC = 14'b1111110111101000; // vC= -536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011001; // iC=-1831 
// vC = 14'b1111111011001000; // vC= -312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000111; // iC=-1977 
// vC = 14'b1111111001001111; // vC= -433 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110010; // iC=-1934 
// vC = 14'b1111111000100101; // vC= -475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b1111111001000000; // vC= -448 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b1111111011001101; // vC= -307 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b1111111001010011; // vC= -429 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b1111111011001001; // vC= -311 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111100; // iC=-1988 
// vC = 14'b1111111010001111; // vC= -369 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100101; // iC=-1819 
// vC = 14'b1111110111010001; // vC= -559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110010; // iC=-1934 
// vC = 14'b1111111000000011; // vC= -509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b1111111010111000; // vC= -328 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b1111110111000001; // vC= -575 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000010; // iC=-1854 
// vC = 14'b1111110110001001; // vC= -631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010110; // iC=-1962 
// vC = 14'b1111110101101010; // vC= -662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111110; // iC=-2050 
// vC = 14'b1111111001100111; // vC= -409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b1111111000100011; // vC= -477 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b1111110101011000; // vC= -680 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b1111110110100010; // vC= -606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b1111111000111011; // vC= -453 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b1111111001001101; // vC= -435 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b1111110110010001; // vC= -623 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000001; // iC=-1791 
// vC = 14'b1111110100101011; // vC= -725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110001; // iC=-1807 
// vC = 14'b1111111000000101; // vC= -507 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000001; // iC=-1855 
// vC = 14'b1111110111001000; // vC= -568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010110; // iC=-1962 
// vC = 14'b1111111000001100; // vC= -500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b1111111000001100; // vC= -500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100010; // iC=-1822 
// vC = 14'b1111110110000010; // vC= -638 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111100; // iC=-1924 
// vC = 14'b1111110101110010; // vC= -654 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b1111110101101000; // vC= -664 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b1111110100111111; // vC= -705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b1111110110101011; // vC= -597 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001111; // iC=-1841 
// vC = 14'b1111110110110000; // vC= -592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b1111110101100011; // vC= -669 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b1111110011001111; // vC= -817 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b1111110110110101; // vC= -587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011000; // iC=-1768 
// vC = 14'b1111110110001110; // vC= -626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100111; // iC=-1881 
// vC = 14'b1111110100101000; // vC= -728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110010; // iC=-1742 
// vC = 14'b1111110010100010; // vC= -862 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110000; // iC=-1744 
// vC = 14'b1111110100011111; // vC= -737 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101101; // iC=-1683 
// vC = 14'b1111110011110110; // vC= -778 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000010; // iC=-1918 
// vC = 14'b1111110010011011; // vC= -869 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111001; // iC=-1863 
// vC = 14'b1111110110011101; // vC= -611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b1111110001111101; // vC= -899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110101; // iC=-1803 
// vC = 14'b1111110110100001; // vC= -607 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110101; // iC=-1675 
// vC = 14'b1111110100010111; // vC= -745 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b1111110100001010; // vC= -758 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011111; // iC=-1825 
// vC = 14'b1111110100000001; // vC= -767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011111; // iC=-1761 
// vC = 14'b1111110010010101; // vC= -875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000101; // iC=-1787 
// vC = 14'b1111110010000111; // vC= -889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001100; // iC=-1716 
// vC = 14'b1111110100100000; // vC= -736 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b1111110011100111; // vC= -793 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011010; // iC=-1702 
// vC = 14'b1111110001001110; // vC= -946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b1111110011000111; // vC= -825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001100; // iC=-1908 
// vC = 14'b1111110011100110; // vC= -794 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b1111110101011001; // vC= -679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b1111110011111011; // vC= -773 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100000; // iC=-1696 
// vC = 14'b1111110000110110; // vC= -970 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011111; // iC=-1825 
// vC = 14'b1111110000100100; // vC= -988 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b1111110010000010; // vC= -894 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b1111110000011000; // vC=-1000 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011001; // iC=-1831 
// vC = 14'b1111110011100001; // vC= -799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001110; // iC=-1842 
// vC = 14'b1111110001010000; // vC= -944 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000010; // iC=-1662 
// vC = 14'b1111110001101101; // vC= -915 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b1111110000101100; // vC= -980 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111001; // iC=-1799 
// vC = 14'b1111110100011000; // vC= -744 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011111; // iC=-1633 
// vC = 14'b1111110100001011; // vC= -757 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b1111110011101011; // vC= -789 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b1111110010001010; // vC= -886 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000101; // iC=-1723 
// vC = 14'b1111110011101000; // vC= -792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100011; // iC=-1757 
// vC = 14'b1111101111010001; // vC=-1071 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111111; // iC=-1601 
// vC = 14'b1111110011100011; // vC= -797 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011001; // iC=-1767 
// vC = 14'b1111110000011010; // vC= -998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010110; // iC=-1834 
// vC = 14'b1111101111110000; // vC=-1040 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011011; // iC=-1573 
// vC = 14'b1111101111000001; // vC=-1087 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b1111110010100110; // vC= -858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010111; // iC=-1769 
// vC = 14'b1111101111001001; // vC=-1079 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000111; // iC=-1657 
// vC = 14'b1111110010111100; // vC= -836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001001; // iC=-1655 
// vC = 14'b1111101110110000; // vC=-1104 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010111; // iC=-1769 
// vC = 14'b1111110001101100; // vC= -916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000000; // iC=-1664 
// vC = 14'b1111110010001100; // vC= -884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010010; // iC=-1646 
// vC = 14'b1111110001000110; // vC= -954 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101100; // iC=-1556 
// vC = 14'b1111101101011001; // vC=-1191 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100110; // iC=-1818 
// vC = 14'b1111110001011110; // vC= -930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001011; // iC=-1589 
// vC = 14'b1111110000001011; // vC=-1013 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000001; // iC=-1727 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011001; // iC=-1703 
// vC = 14'b1111110000110010; // vC= -974 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b1111101101100010; // vC=-1182 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111011; // iC=-1669 
// vC = 14'b1111110000111111; // vC= -961 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000101; // iC=-1659 
// vC = 14'b1111101100111010; // vC=-1222 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011111; // iC=-1569 
// vC = 14'b1111101111110000; // vC=-1040 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001001; // iC=-1783 
// vC = 14'b1111101101110110; // vC=-1162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011111; // iC=-1697 
// vC = 14'b1111110000100000; // vC= -992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011111; // iC=-1633 
// vC = 14'b1111110000111010; // vC= -966 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111001; // iC=-1671 
// vC = 14'b1111101100001001; // vC=-1271 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100010; // iC=-1502 
// vC = 14'b1111101101101000; // vC=-1176 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100001; // iC=-1631 
// vC = 14'b1111101101000101; // vC=-1211 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101001; // iC=-1687 
// vC = 14'b1111101101011101; // vC=-1187 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010101; // iC=-1515 
// vC = 14'b1111101100010111; // vC=-1257 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001101; // iC=-1459 
// vC = 14'b1111101101010011; // vC=-1197 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110111; // iC=-1545 
// vC = 14'b1111101111100100; // vC=-1052 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111001; // iC=-1735 
// vC = 14'b1111101100010010; // vC=-1262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000000; // iC=-1536 
// vC = 14'b1111101011110111; // vC=-1289 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100100; // iC=-1564 
// vC = 14'b1111101100000111; // vC=-1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000111; // iC=-1657 
// vC = 14'b1111101100100110; // vC=-1242 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010101; // iC=-1579 
// vC = 14'b1111101111110100; // vC=-1036 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110011; // iC=-1485 
// vC = 14'b1111101100001001; // vC=-1271 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111100; // iC=-1540 
// vC = 14'b1111101110111010; // vC=-1094 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110101; // iC=-1483 
// vC = 14'b1111101101001011; // vC=-1205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010001; // iC=-1455 
// vC = 14'b1111101011100011; // vC=-1309 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110101; // iC=-1547 
// vC = 14'b1111101010111111; // vC=-1345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010111; // iC=-1577 
// vC = 14'b1111101101010000; // vC=-1200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111111; // iC=-1601 
// vC = 14'b1111101100001111; // vC=-1265 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100111; // iC=-1497 
// vC = 14'b1111101101000001; // vC=-1215 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100100; // iC=-1500 
// vC = 14'b1111101101101001; // vC=-1175 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101010; // iC=-1430 
// vC = 14'b1111101011010110; // vC=-1322 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000011; // iC=-1597 
// vC = 14'b1111101010011100; // vC=-1380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111000; // iC=-1544 
// vC = 14'b1111101100001011; // vC=-1269 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100001; // iC=-1439 
// vC = 14'b1111101011111101; // vC=-1283 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010000; // iC=-1392 
// vC = 14'b1111101100001010; // vC=-1270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011111; // iC=-1441 
// vC = 14'b1111101001100111; // vC=-1433 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110011; // iC=-1549 
// vC = 14'b1111101100101010; // vC=-1238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010001; // iC=-1455 
// vC = 14'b1111101011011101; // vC=-1315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011011; // iC=-1509 
// vC = 14'b1111101110010001; // vC=-1135 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110110; // iC=-1418 
// vC = 14'b1111101100001011; // vC=-1269 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100101; // iC=-1499 
// vC = 14'b1111101101100110; // vC=-1178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101000; // iC=-1560 
// vC = 14'b1111101001110011; // vC=-1421 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000010; // iC=-1470 
// vC = 14'b1111101101100011; // vC=-1181 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100000; // iC=-1568 
// vC = 14'b1111101010000101; // vC=-1403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100101; // iC=-1307 
// vC = 14'b1111101001000011; // vC=-1469 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111111; // iC=-1537 
// vC = 14'b1111101001001110; // vC=-1458 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010110; // iC=-1386 
// vC = 14'b1111101001000000; // vC=-1472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001101; // iC=-1459 
// vC = 14'b1111101100110101; // vC=-1227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001000; // iC=-1528 
// vC = 14'b1111101001000111; // vC=-1465 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010010; // iC=-1454 
// vC = 14'b1111101001000000; // vC=-1472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110011; // iC=-1357 
// vC = 14'b1111101000000101; // vC=-1531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100000; // iC=-1376 
// vC = 14'b1111101001011100; // vC=-1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110100; // iC=-1292 
// vC = 14'b1111101100000001; // vC=-1279 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100100; // iC=-1244 
// vC = 14'b1111101011001110; // vC=-1330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001110; // iC=-1330 
// vC = 14'b1111101001111000; // vC=-1416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110110; // iC=-1546 
// vC = 14'b1111101011100101; // vC=-1307 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011001; // iC=-1255 
// vC = 14'b1111101001001101; // vC=-1459 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110101; // iC=-1291 
// vC = 14'b1111101011100100; // vC=-1308 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000000; // iC=-1216 
// vC = 14'b1111101011111010; // vC=-1286 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101101; // iC=-1363 
// vC = 14'b1111101000101010; // vC=-1494 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001011; // iC=-1397 
// vC = 14'b1111101011010000; // vC=-1328 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111010; // iC=-1286 
// vC = 14'b1111101000100010; // vC=-1502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111111; // iC=-1281 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010111; // iC=-1513 
// vC = 14'b1111101010110100; // vC=-1356 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000001; // iC=-1279 
// vC = 14'b1111101000111101; // vC=-1475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101000; // iC=-1432 
// vC = 14'b1111101010101111; // vC=-1361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100011; // iC=-1373 
// vC = 14'b1111100111101000; // vC=-1560 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001010; // iC=-1270 
// vC = 14'b1111101010000010; // vC=-1406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110111; // iC=-1289 
// vC = 14'b1111101010100101; // vC=-1371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010011; // iC=-1389 
// vC = 14'b1111101000010101; // vC=-1515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000111; // iC=-1273 
// vC = 14'b1111100110101111; // vC=-1617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111011; // iC=-1349 
// vC = 14'b1111101000011010; // vC=-1510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111001; // iC=-1223 
// vC = 14'b1111100111011001; // vC=-1575 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000101; // iC=-1339 
// vC = 14'b1111100111001110; // vC=-1586 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010110; // iC=-1322 
// vC = 14'b1111101001111001; // vC=-1415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110011; // iC=-1229 
// vC = 14'b1111100111110011; // vC=-1549 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101101; // iC=-1235 
// vC = 14'b1111100111001110; // vC=-1586 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000111; // iC=-1273 
// vC = 14'b1111100110100000; // vC=-1632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100010; // iC=-1374 
// vC = 14'b1111101010000101; // vC=-1403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011011; // iC=-1317 
// vC = 14'b1111101010010101; // vC=-1387 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111101; // iC=-1219 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010100; // iC=-1260 
// vC = 14'b1111101010100001; // vC=-1375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111011; // iC=-1157 
// vC = 14'b1111101001000001; // vC=-1471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001000; // iC=-1400 
// vC = 14'b1111100110010111; // vC=-1641 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010100; // iC=-1388 
// vC = 14'b1111100110000111; // vC=-1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101010; // iC=-1174 
// vC = 14'b1111101000011101; // vC=-1507 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110101; // iC=-1355 
// vC = 14'b1111100110001010; // vC=-1654 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100100; // iC=-1372 
// vC = 14'b1111100110000101; // vC=-1659 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010111; // iC=-1193 
// vC = 14'b1111100110110011; // vC=-1613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010100; // iC=-1132 
// vC = 14'b1111100111111000; // vC=-1544 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111000; // iC=-1288 
// vC = 14'b1111101001011100; // vC=-1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000000; // iC=-1344 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101011; // iC=-1301 
// vC = 14'b1111101000111000; // vC=-1480 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011000; // iC=-1256 
// vC = 14'b1111100110100010; // vC=-1630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010001; // iC=-1263 
// vC = 14'b1111100111100010; // vC=-1566 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101001; // iC=-1175 
// vC = 14'b1111101000011010; // vC=-1510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101010; // iC=-1238 
// vC = 14'b1111101000001001; // vC=-1527 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110111; // iC=-1289 
// vC = 14'b1111101000111000; // vC=-1480 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101010; // iC=-1302 
// vC = 14'b1111101001001101; // vC=-1459 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110000; // iC=-1168 
// vC = 14'b1111100110110110; // vC=-1610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100011; // iC=-1309 
// vC = 14'b1111100101011000; // vC=-1704 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110001; // iC=-1231 
// vC = 14'b1111100111100011; // vC=-1565 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100110; // iC= -986 
// vC = 14'b1111100111011110; // vC=-1570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111010; // iC=-1094 
// vC = 14'b1111101000001101; // vC=-1523 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010110; // iC=-1130 
// vC = 14'b1111100111001010; // vC=-1590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110001; // iC=-1039 
// vC = 14'b1111100100101010; // vC=-1750 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001001; // iC=-1015 
// vC = 14'b1111101000000100; // vC=-1532 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111101; // iC=-1219 
// vC = 14'b1111100110110000; // vC=-1616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011101; // iC=-1187 
// vC = 14'b1111100100110110; // vC=-1738 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100101; // iC=-1179 
// vC = 14'b1111100110001100; // vC=-1652 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100110; // iC=-1178 
// vC = 14'b1111100110011101; // vC=-1635 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000111; // iC=-1145 
// vC = 14'b1111100100111010; // vC=-1734 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000001; // iC=-1151 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100010; // iC= -926 
// vC = 14'b1111100101101101; // vC=-1683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110000; // iC=-1168 
// vC = 14'b1111100111000100; // vC=-1596 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000010; // iC=-1022 
// vC = 14'b1111100011001011; // vC=-1845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000001; // iC=-1023 
// vC = 14'b1111100101101010; // vC=-1686 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101111; // iC=-1169 
// vC = 14'b1111100011100111; // vC=-1817 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000000; // iC= -960 
// vC = 14'b1111100110110000; // vC=-1616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110110; // iC= -906 
// vC = 14'b1111100011000101; // vC=-1851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001010; // iC= -950 
// vC = 14'b1111100011111001; // vC=-1799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001110; // iC=-1138 
// vC = 14'b1111100101000000; // vC=-1728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000100; // iC= -956 
// vC = 14'b1111100100110010; // vC=-1742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101001; // iC= -855 
// vC = 14'b1111100010110111; // vC=-1865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001001; // iC=-1015 
// vC = 14'b1111100010100101; // vC=-1883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000000; // iC= -896 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101101; // iC= -915 
// vC = 14'b1111100110001110; // vC=-1650 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011000; // iC= -872 
// vC = 14'b1111100100111110; // vC=-1730 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101001; // iC=-1047 
// vC = 14'b1111100111000010; // vC=-1598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100110; // iC= -922 
// vC = 14'b1111100110111000; // vC=-1608 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010011; // iC=-1069 
// vC = 14'b1111100100011111; // vC=-1761 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111010; // iC=-1094 
// vC = 14'b1111100011101000; // vC=-1816 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111011; // iC=-1029 
// vC = 14'b1111100110111000; // vC=-1608 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001001; // iC= -887 
// vC = 14'b1111100001111011; // vC=-1925 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111101; // iC= -835 
// vC = 14'b1111100101100000; // vC=-1696 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110010; // iC=-1038 
// vC = 14'b1111100011100100; // vC=-1820 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111100; // iC=-1092 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010001; // iC= -815 
// vC = 14'b1111100101011011; // vC=-1701 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000000; // iC= -960 
// vC = 14'b1111100101100111; // vC=-1689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000011; // iC= -765 
// vC = 14'b1111100001111100; // vC=-1924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001111; // iC= -753 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011111; // iC= -929 
// vC = 14'b1111100001101001; // vC=-1943 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010100; // iC=-1004 
// vC = 14'b1111100101010111; // vC=-1705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101010; // iC= -918 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111101; // iC= -963 
// vC = 14'b1111100010010011; // vC=-1901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101000; // iC= -856 
// vC = 14'b1111100010010011; // vC=-1901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101111; // iC= -913 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100110; // iC= -794 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011110; // iC= -866 
// vC = 14'b1111100010001011; // vC=-1909 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001001; // iC= -823 
// vC = 14'b1111100100101100; // vC=-1748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001010; // iC= -950 
// vC = 14'b1111100001101001; // vC=-1943 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101110; // iC= -722 
// vC = 14'b1111100011011001; // vC=-1831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000101; // iC= -763 
// vC = 14'b1111100100011000; // vC=-1768 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111011; // iC= -901 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110000; // iC= -720 
// vC = 14'b1111100011111011; // vC=-1797 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011001; // iC= -871 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111011; // iC= -645 
// vC = 14'b1111100010000010; // vC=-1918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010011; // iC= -877 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000111; // iC= -633 
// vC = 14'b1111100010101110; // vC=-1874 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111101; // iC= -771 
// vC = 14'b1111100001110101; // vC=-1931 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100100; // iC= -860 
// vC = 14'b1111100011101110; // vC=-1810 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100001; // iC= -671 
// vC = 14'b1111100100011010; // vC=-1766 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001000; // iC= -888 
// vC = 14'b1111100011111011; // vC=-1797 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110001; // iC= -655 
// vC = 14'b1111100100010011; // vC=-1773 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110101; // iC= -651 
// vC = 14'b1111100001001100; // vC=-1972 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110000; // iC= -720 
// vC = 14'b1111100011001111; // vC=-1841 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111011; // iC= -581 
// vC = 14'b1111100100000001; // vC=-1791 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011110; // iC= -610 
// vC = 14'b1111100010101001; // vC=-1879 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101010; // iC= -854 
// vC = 14'b1111100010000101; // vC=-1915 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001111; // iC= -625 
// vC = 14'b1111100010001101; // vC=-1907 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101100; // iC= -788 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000011; // iC= -701 
// vC = 14'b1111100001101110; // vC=-1938 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001010; // iC= -630 
// vC = 14'b1111100001010101; // vC=-1963 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011011; // iC= -549 
// vC = 14'b1111100011100001; // vC=-1823 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111010; // iC= -774 
// vC = 14'b1111100100001100; // vC=-1780 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110010; // iC= -654 
// vC = 14'b1111100001100111; // vC=-1945 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010010; // iC= -558 
// vC = 14'b1111100001101101; // vC=-1939 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001000; // iC= -504 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001101; // iC= -499 
// vC = 14'b1111100000010110; // vC=-2026 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110111; // iC= -713 
// vC = 14'b1111100100000010; // vC=-1790 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111000; // iC= -520 
// vC = 14'b1111100100011010; // vC=-1766 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101011; // iC= -725 
// vC = 14'b1111100001001101; // vC=-1971 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100111; // iC= -473 
// vC = 14'b1111100000001010; // vC=-2038 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110110; // iC= -714 
// vC = 14'b1111100011001010; // vC=-1846 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110111; // iC= -585 
// vC = 14'b1111100001001101; // vC=-1971 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001011; // iC= -501 
// vC = 14'b1111100011010001; // vC=-1839 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101111; // iC= -657 
// vC = 14'b1111100001111001; // vC=-1927 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111111; // iC= -449 
// vC = 14'b1111100011010010; // vC=-1838 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100011; // iC= -669 
// vC = 14'b1111100011111011; // vC=-1797 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000111; // iC= -441 
// vC = 14'b1111011111101101; // vC=-2067 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111000; // iC= -584 
// vC = 14'b1111011111011011; // vC=-2085 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100110; // iC= -474 
// vC = 14'b1111011111100101; // vC=-2075 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100011; // iC= -413 
// vC = 14'b1111100001111011; // vC=-1925 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110011; // iC= -397 
// vC = 14'b1111100011001101; // vC=-1843 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111100; // iC= -516 
// vC = 14'b1111100001110110; // vC=-1930 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101110; // iC= -402 
// vC = 14'b1111100000101101; // vC=-2003 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010011; // iC= -429 
// vC = 14'b1111100011010010; // vC=-1838 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010001; // iC= -303 
// vC = 14'b1111100000011110; // vC=-2018 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010010; // iC= -494 
// vC = 14'b1111100011100100; // vC=-1820 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100110; // iC= -346 
// vC = 14'b1111100000010001; // vC=-2031 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110111; // iC= -201 
// vC = 14'b1111100010110010; // vC=-1870 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001101; // iC= -179 
// vC = 14'b1111100011100111; // vC=-1817 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111000; // iC= -456 
// vC = 14'b1111100011101111; // vC=-1809 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111000; // iC= -392 
// vC = 14'b1111100011101001; // vC=-1815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111011; // iC= -197 
// vC = 14'b1111100011100100; // vC=-1820 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101111; // iC= -401 
// vC = 14'b1111100000010000; // vC=-2032 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101011; // iC= -149 
// vC = 14'b1111011110111101; // vC=-2115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011001; // iC= -359 
// vC = 14'b1111011111111101; // vC=-2051 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000111; // iC= -185 
// vC = 14'b1111100000111111; // vC=-1985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010111; // iC= -233 
// vC = 14'b1111100001111010; // vC=-1926 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101110; // iC= -146 
// vC = 14'b1111100000111111; // vC=-1985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001011; // iC= -245 
// vC = 14'b1111011111101111; // vC=-2065 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010010; // iC= -302 
// vC = 14'b1111100001110000; // vC=-1936 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111000; // iC= -200 
// vC = 14'b1111100011110100; // vC=-1804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011010; // iC=   26 
// vC = 14'b1111100000000111; // vC=-2041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010011; // iC=  -45 
// vC = 14'b1111100011100101; // vC=-1819 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001000; // iC=  -56 
// vC = 14'b1111100010100011; // vC=-1885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000110; // iC= -122 
// vC = 14'b1111100000000010; // vC=-2046 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010100; // iC=   20 
// vC = 14'b1111011111111010; // vC=-2054 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100101; // iC=  -91 
// vC = 14'b1111100010001100; // vC=-1908 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100111; // iC=  103 
// vC = 14'b1111100001110011; // vC=-1933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111010; // iC=  122 
// vC = 14'b1111011111010010; // vC=-2094 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000000; // iC=  -64 
// vC = 14'b1111100000111111; // vC=-1985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111011101; // iC=  -35 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110000; // iC=  240 
// vC = 14'b1111011110111011; // vC=-2117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000010; // iC=  130 
// vC = 14'b1111100010001100; // vC=-1908 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001110; // iC=   14 
// vC = 14'b1111100010011101; // vC=-1891 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000111001; // iC=   57 
// vC = 14'b1111100011111010; // vC=-1798 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111111; // iC=  255 
// vC = 14'b1111100000111100; // vC=-1988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000111000; // iC=   56 
// vC = 14'b1111100011000101; // vC=-1851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010101; // iC=  213 
// vC = 14'b1111100000010101; // vC=-2027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111000; // iC=  184 
// vC = 14'b1111100001001000; // vC=-1976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011100; // iC=  412 
// vC = 14'b1111100010011111; // vC=-1889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111110; // iC=  254 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011011; // iC=  411 
// vC = 14'b1111100001100100; // vC=-1948 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100101; // iC=  229 
// vC = 14'b1111100001001011; // vC=-1973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100010; // iC=  418 
// vC = 14'b1111100010000100; // vC=-1916 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000101; // iC=  453 
// vC = 14'b1111100000100101; // vC=-2011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001000; // iC=  520 
// vC = 14'b1111100010111001; // vC=-1863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011011; // iC=  347 
// vC = 14'b1111100001000001; // vC=-1983 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100010; // iC=  546 
// vC = 14'b1111100010000100; // vC=-1916 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100000; // iC=  544 
// vC = 14'b1111100010101001; // vC=-1879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010100; // iC=  660 
// vC = 14'b1111100001000001; // vC=-1983 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000001; // iC=  577 
// vC = 14'b1111100010000000; // vC=-1920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010111; // iC=  471 
// vC = 14'b1111100000101101; // vC=-2003 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101111; // iC=  623 
// vC = 14'b1111100010100000; // vC=-1888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111100; // iC=  444 
// vC = 14'b1111100010100101; // vC=-1883 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011110; // iC=  606 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111011; // iC=  635 
// vC = 14'b1111100100100000; // vC=-1760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111110; // iC=  766 
// vC = 14'b1111100000101111; // vC=-2001 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000001; // iC=  833 
// vC = 14'b1111100010011110; // vC=-1890 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100111; // iC=  807 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110100; // iC=  692 
// vC = 14'b1111100100001011; // vC=-1781 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001100; // iC=  652 
// vC = 14'b1111100100110110; // vC=-1738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111000; // iC=  888 
// vC = 14'b1111100011111000; // vC=-1800 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110001; // iC=  881 
// vC = 14'b1111100000111010; // vC=-1990 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000110; // iC=  710 
// vC = 14'b1111100101001001; // vC=-1719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100111; // iC=  807 
// vC = 14'b1111100011011111; // vC=-1825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100111; // iC=  743 
// vC = 14'b1111100011001100; // vC=-1844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001110; // iC=  782 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111000; // iC=  760 
// vC = 14'b1111100100010111; // vC=-1769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001010; // iC= 1034 
// vC = 14'b1111100100010111; // vC=-1769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001010; // iC= 1098 
// vC = 14'b1111100001011110; // vC=-1954 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110011; // iC= 1011 
// vC = 14'b1111100001100001; // vC=-1951 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111101; // iC= 1021 
// vC = 14'b1111100000111100; // vC=-1988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101100; // iC= 1068 
// vC = 14'b1111100001111100; // vC=-1924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111111; // iC=  959 
// vC = 14'b1111100001110000; // vC=-1936 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001010; // iC=  906 
// vC = 14'b1111100001001000; // vC=-1976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011010; // iC=  986 
// vC = 14'b1111100011100000; // vC=-1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111111; // iC=  959 
// vC = 14'b1111100011010111; // vC=-1833 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100010; // iC= 1122 
// vC = 14'b1111100001111010; // vC=-1926 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000001; // iC= 1217 
// vC = 14'b1111100101011111; // vC=-1697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010011; // iC= 1235 
// vC = 14'b1111100001001101; // vC=-1971 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001001; // iC= 1225 
// vC = 14'b1111100011011011; // vC=-1829 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010111; // iC= 1047 
// vC = 14'b1111100100101101; // vC=-1747 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010101; // iC= 1301 
// vC = 14'b1111100110010001; // vC=-1647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000011; // iC= 1219 
// vC = 14'b1111100110000000; // vC=-1664 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110111; // iC= 1143 
// vC = 14'b1111100110101101; // vC=-1619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100101; // iC= 1125 
// vC = 14'b1111100010100011; // vC=-1885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100010; // iC= 1378 
// vC = 14'b1111100011110100; // vC=-1804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111101; // iC= 1149 
// vC = 14'b1111100010000111; // vC=-1913 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001101; // iC= 1357 
// vC = 14'b1111100010000011; // vC=-1917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110001; // iC= 1393 
// vC = 14'b1111100101100001; // vC=-1695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100100; // iC= 1380 
// vC = 14'b1111100011001000; // vC=-1848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010011; // iC= 1427 
// vC = 14'b1111100011001010; // vC=-1846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010101; // iC= 1493 
// vC = 14'b1111100100100000; // vC=-1760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100010; // iC= 1250 
// vC = 14'b1111100011011011; // vC=-1829 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000010; // iC= 1410 
// vC = 14'b1111100110111000; // vC=-1608 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101100; // iC= 1452 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000111; // iC= 1479 
// vC = 14'b1111100110110011; // vC=-1613 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110110; // iC= 1590 
// vC = 14'b1111100111110111; // vC=-1545 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110111; // iC= 1399 
// vC = 14'b1111100111010010; // vC=-1582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001010; // iC= 1354 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100110; // iC= 1510 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110101; // iC= 1397 
// vC = 14'b1111100110100011; // vC=-1629 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000111; // iC= 1607 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101011; // iC= 1515 
// vC = 14'b1111100101010011; // vC=-1709 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111011; // iC= 1723 
// vC = 14'b1111100111110010; // vC=-1550 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101111; // iC= 1711 
// vC = 14'b1111100110000000; // vC=-1664 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011111; // iC= 1695 
// vC = 14'b1111100110100101; // vC=-1627 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000100; // iC= 1476 
// vC = 14'b1111100101110010; // vC=-1678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101000; // iC= 1512 
// vC = 14'b1111101000110100; // vC=-1484 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101101; // iC= 1581 
// vC = 14'b1111100111010111; // vC=-1577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111101; // iC= 1533 
// vC = 14'b1111100111100101; // vC=-1563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110000; // iC= 1584 
// vC = 14'b1111100111000111; // vC=-1593 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011101; // iC= 1565 
// vC = 14'b1111101000100110; // vC=-1498 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b1111101001000000; // vC=-1472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111010; // iC= 1722 
// vC = 14'b1111101000011111; // vC=-1505 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011111; // iC= 1631 
// vC = 14'b1111101001100101; // vC=-1435 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110110; // iC= 1654 
// vC = 14'b1111101001100100; // vC=-1436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b1111101001011001; // vC=-1447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b1111100101101000; // vC=-1688 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111101; // iC= 1661 
// vC = 14'b1111101010000000; // vC=-1408 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000100; // iC= 1796 
// vC = 14'b1111100111100001; // vC=-1567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001010; // iC= 1674 
// vC = 14'b1111101000110010; // vC=-1486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100100; // iC= 1636 
// vC = 14'b1111101010010011; // vC=-1389 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001010; // iC= 1802 
// vC = 14'b1111100111101001; // vC=-1559 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b1111101001100010; // vC=-1438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100011; // iC= 1699 
// vC = 14'b1111101010100110; // vC=-1370 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001110; // iC= 1806 
// vC = 14'b1111101010001101; // vC=-1395 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011011; // iC= 1755 
// vC = 14'b1111100111010101; // vC=-1579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111101000010000; // vC=-1520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000100; // iC= 1988 
// vC = 14'b1111101010010010; // vC=-1390 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111011; // iC= 1851 
// vC = 14'b1111101001011000; // vC=-1448 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b1111101000110001; // vC=-1487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100010; // iC= 1890 
// vC = 14'b1111101000010011; // vC=-1517 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110000; // iC= 1968 
// vC = 14'b1111100111101101; // vC=-1555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011010; // iC= 1754 
// vC = 14'b1111101010010110; // vC=-1386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001001; // iC= 1865 
// vC = 14'b1111101011110000; // vC=-1296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100101; // iC= 1829 
// vC = 14'b1111101010100101; // vC=-1371 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b1111101011000010; // vC=-1342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001111; // iC= 2063 
// vC = 14'b1111101000000111; // vC=-1529 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101001; // iC= 1897 
// vC = 14'b1111101100011000; // vC=-1256 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111101; // iC= 1789 
// vC = 14'b1111101000101000; // vC=-1496 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001111; // iC= 1871 
// vC = 14'b1111101101000010; // vC=-1214 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010111; // iC= 1815 
// vC = 14'b1111101000111010; // vC=-1478 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101111; // iC= 1903 
// vC = 14'b1111101011010000; // vC=-1328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111101100101000; // vC=-1240 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000000; // iC= 2112 
// vC = 14'b1111101100010100; // vC=-1260 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b1111101001111000; // vC=-1416 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111101010101100; // vC=-1364 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011110; // iC= 1822 
// vC = 14'b1111101011000010; // vC=-1342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101110; // iC= 1966 
// vC = 14'b1111101010111010; // vC=-1350 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011000; // iC= 2136 
// vC = 14'b1111101100010001; // vC=-1263 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b1111101011111001; // vC=-1287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011110; // iC= 2014 
// vC = 14'b1111101011011101; // vC=-1315 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b1111101101010010; // vC=-1198 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001101; // iC= 1997 
// vC = 14'b1111101011110010; // vC=-1294 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b1111101101101111; // vC=-1169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b1111101101110000; // vC=-1168 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b1111101110000001; // vC=-1151 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001000; // iC= 1864 
// vC = 14'b1111101111100001; // vC=-1055 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b1111101010111100; // vC=-1348 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010110; // iC= 2134 
// vC = 14'b1111101100100001; // vC=-1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000100; // iC= 2116 
// vC = 14'b1111101111110100; // vC=-1036 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b1111101110111001; // vC=-1095 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b1111101011110101; // vC=-1291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101110; // iC= 2094 
// vC = 14'b1111101111011110; // vC=-1058 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b1111101100110010; // vC=-1230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b1111101111100101; // vC=-1051 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b1111101100010110; // vC=-1258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111110; // iC= 2046 
// vC = 14'b1111101101000001; // vC=-1215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b1111101101100100; // vC=-1180 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110111; // iC= 1911 
// vC = 14'b1111101100111100; // vC=-1220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010101; // iC= 1877 
// vC = 14'b1111101100111011; // vC=-1221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000000; // iC= 2112 
// vC = 14'b1111110000001000; // vC=-1016 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b1111101111111100; // vC=-1028 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100001; // iC= 2145 
// vC = 14'b1111101101110101; // vC=-1163 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111101111011101; // vC=-1059 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111110; // iC= 2046 
// vC = 14'b1111101111110110; // vC=-1034 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001011; // iC= 2123 
// vC = 14'b1111101110101010; // vC=-1110 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b1111110000101110; // vC= -978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010100; // iC= 2132 
// vC = 14'b1111101111101000; // vC=-1048 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011010; // iC= 2138 
// vC = 14'b1111101111000110; // vC=-1082 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101010; // iC= 1898 
// vC = 14'b1111101111010010; // vC=-1070 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b1111101111011101; // vC=-1059 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111110; // iC= 2174 
// vC = 14'b1111101110101010; // vC=-1110 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111101110010100; // vC=-1132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000100; // iC= 1988 
// vC = 14'b1111101111110110; // vC=-1034 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110011; // iC= 2163 
// vC = 14'b1111110001101111; // vC= -913 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101100; // iC= 1900 
// vC = 14'b1111110000110111; // vC= -969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010111; // iC= 2199 
// vC = 14'b1111110010101111; // vC= -849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b1111110001010001; // vC= -943 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000011; // iC= 2051 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b1111110001011101; // vC= -931 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011001; // iC= 2137 
// vC = 14'b1111110001111011; // vC= -901 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011100; // iC= 2012 
// vC = 14'b1111110011100110; // vC= -794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010101; // iC= 2197 
// vC = 14'b1111110011000010; // vC= -830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001110; // iC= 2126 
// vC = 14'b1111110100110110; // vC= -714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b1111110100001111; // vC= -753 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100101; // iC= 2213 
// vC = 14'b1111110001000000; // vC= -960 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111110010110110; // vC= -842 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101111; // iC= 2095 
// vC = 14'b1111110100100101; // vC= -731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111111; // iC= 1983 
// vC = 14'b1111110101001011; // vC= -693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b1111110100001010; // vC= -758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000001; // iC= 2177 
// vC = 14'b1111110001011111; // vC= -929 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b1111110110000011; // vC= -637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100010; // iC= 2146 
// vC = 14'b1111110101010010; // vC= -686 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000100; // iC= 1924 
// vC = 14'b1111110011111010; // vC= -774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010101; // iC= 2133 
// vC = 14'b1111110010100000; // vC= -864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b1111110101100011; // vC= -669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011111; // iC= 2143 
// vC = 14'b1111110011011101; // vC= -803 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100101; // iC= 2149 
// vC = 14'b1111110010101000; // vC= -856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b1111110100101111; // vC= -721 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000100; // iC= 1924 
// vC = 14'b1111110010110101; // vC= -843 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011110; // iC= 2014 
// vC = 14'b1111110011011001; // vC= -807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110000; // iC= 2096 
// vC = 14'b1111110100111100; // vC= -708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b1111110010110010; // vC= -846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b1111110100110100; // vC= -716 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b1111111000000010; // vC= -510 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010101; // iC= 2133 
// vC = 14'b1111110110110000; // vC= -592 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010001; // iC= 2001 
// vC = 14'b1111110011011010; // vC= -806 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b1111110100100101; // vC= -731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111110; // iC= 2174 
// vC = 14'b1111110110010101; // vC= -619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101111; // iC= 2159 
// vC = 14'b1111110110000000; // vC= -640 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111011; // iC= 1915 
// vC = 14'b1111110100100010; // vC= -734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b1111110110011010; // vC= -614 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101000; // iC= 2216 
// vC = 14'b1111110110010010; // vC= -622 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b1111110100010001; // vC= -751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000000; // iC= 2240 
// vC = 14'b1111110100101011; // vC= -725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111110110001100; // vC= -628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b1111110111110110; // vC= -522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101001; // iC= 2217 
// vC = 14'b1111110111001010; // vC= -566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010001; // iC= 2065 
// vC = 14'b1111111001000000; // vC= -448 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010010; // iC= 2002 
// vC = 14'b1111110110100000; // vC= -608 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100011; // iC= 2147 
// vC = 14'b1111110101011101; // vC= -675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b1111110110111011; // vC= -581 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001101; // iC= 2189 
// vC = 14'b1111110111110111; // vC= -521 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101110; // iC= 2222 
// vC = 14'b1111111000100010; // vC= -478 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111110111111010; // vC= -518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111111010001001; // vC= -375 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b1111110110001010; // vC= -630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011110; // iC= 2142 
// vC = 14'b1111111001010100; // vC= -428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111110110111000; // vC= -584 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100010; // iC= 2146 
// vC = 14'b1111111011000000; // vC= -320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000101; // iC= 2117 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010001; // iC= 2001 
// vC = 14'b1111110110110011; // vC= -589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111110111001101; // vC= -563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110101; // iC= 2037 
// vC = 14'b1111111010101000; // vC= -344 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b1111111001010110; // vC= -426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b1111111011000100; // vC= -316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b1111111001000110; // vC= -442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100111; // iC= 2087 
// vC = 14'b1111111000010001; // vC= -495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001101; // iC= 2189 
// vC = 14'b1111111010101001; // vC= -343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111111001100000; // vC= -416 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110000; // iC= 2032 
// vC = 14'b1111111000100010; // vC= -478 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100000; // iC= 2016 
// vC = 14'b1111111001101111; // vC= -401 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b1111111010001101; // vC= -371 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000101; // iC= 2053 
// vC = 14'b1111111010101111; // vC= -337 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b1111111001101011; // vC= -405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b1111111101011000; // vC= -168 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b1111111011101001; // vC= -279 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111001; // iC= 2169 
// vC = 14'b1111111100100010; // vC= -222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111111010000111; // vC= -377 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111111001011111; // vC= -417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b1111111011110011; // vC= -269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b1111111100110110; // vC= -202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110011; // iC= 1971 
// vC = 14'b1111111011000101; // vC= -315 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101001; // iC= 2217 
// vC = 14'b1111111010010110; // vC= -362 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b1111111100000010; // vC= -254 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110110; // iC= 1910 
// vC = 14'b1111111010110100; // vC= -332 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b1111111110011000; // vC= -104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b1111111010110011; // vC= -333 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001011; // iC= 2123 
// vC = 14'b1111111011110010; // vC= -270 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110110; // iC= 2038 
// vC = 14'b1111111111011010; // vC=  -38 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b1111111100111111; // vC= -193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110001; // iC= 2097 
// vC = 14'b1111111100001000; // vC= -248 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000000; // iC= 2176 
// vC = 14'b1111111100111010; // vC= -198 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011000; // iC= 2072 
// vC = 14'b1111111110101110; // vC=  -82 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b1111111100101101; // vC= -211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010000; // iC= 2192 
// vC = 14'b1111111110000011; // vC= -125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011100; // iC= 2140 
// vC = 14'b1111111100010101; // vC= -235 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010011; // iC= 2067 
// vC = 14'b0000000000101100; // vC=   44 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b1111111110010010; // vC= -110 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110001; // iC= 2097 
// vC = 14'b0000000000001110; // vC=   14 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001011; // iC= 2123 
// vC = 14'b1111111111100111; // vC=  -25 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b0000000000100010; // vC=   34 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001000; // iC= 2120 
// vC = 14'b0000000000101011; // vC=   43 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b1111111110000100; // vC= -124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110101; // iC= 2101 
// vC = 14'b1111111101111110; // vC= -130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b0000000000111010; // vC=   58 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101000; // iC= 2024 
// vC = 14'b1111111101100111; // vC= -153 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011001; // iC= 2137 
// vC = 14'b1111111110001110; // vC= -114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b0000000001011111; // vC=   95 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000100; // iC= 1988 
// vC = 14'b0000000010010110; // vC=  150 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011000; // iC= 1880 
// vC = 14'b0000000001100010; // vC=   98 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111000; // iC= 1912 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b1111111111010001; // vC=  -47 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b0000000000010110; // vC=   22 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100011; // iC= 2083 
// vC = 14'b1111111110111111; // vC=  -65 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100111; // iC= 1895 
// vC = 14'b0000000001011111; // vC=   95 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111100; // iC= 1980 
// vC = 14'b1111111111100100; // vC=  -28 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b0000000010000100; // vC=  132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101001; // iC= 1897 
// vC = 14'b0000000001111000; // vC=  120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b0000000000010101; // vC=   21 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b0000000000000100; // vC=    4 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111000; // iC= 2168 
// vC = 14'b0000000001000011; // vC=   67 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b0000000100010110; // vC=  278 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b0000000011110110; // vC=  246 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111000; // iC= 1976 
// vC = 14'b0000000011101001; // vC=  233 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b0000000000111011; // vC=   59 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111000; // iC= 2104 
// vC = 14'b0000000011110110; // vC=  246 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b0000000001000110; // vC=   70 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111110; // iC= 1854 
// vC = 14'b0000000001111111; // vC=  127 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011111; // iC= 1887 
// vC = 14'b0000000000100011; // vC=   35 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b0000000001100000; // vC=   96 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b0000000011011000; // vC=  216 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010110; // iC= 2070 
// vC = 14'b0000000011101010; // vC=  234 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b0000000001101110; // vC=  110 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011011; // iC= 2075 
// vC = 14'b0000000011110000; // vC=  240 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111110; // iC= 2110 
// vC = 14'b0000000001110011; // vC=  115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b0000000101011000; // vC=  344 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010001; // iC= 1937 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000100; // iC= 2116 
// vC = 14'b0000000010110100; // vC=  180 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b0000000101101000; // vC=  360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b0000000101010010; // vC=  338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b0000000101001111; // vC=  335 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000000; // iC= 1984 
// vC = 14'b0000000010011111; // vC=  159 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010100; // iC= 2068 
// vC = 14'b0000000011111111; // vC=  255 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b0000000110101011; // vC=  427 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b0000000100110001; // vC=  305 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b0000000111100000; // vC=  480 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000011; // iC= 1923 
// vC = 14'b0000000111001100; // vC=  460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b0000000011100110; // vC=  230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b0000000111010001; // vC=  465 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b0000000011111001; // vC=  249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b0000000111110001; // vC=  497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101001; // iC= 1897 
// vC = 14'b0000000100011000; // vC=  280 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110000; // iC= 2032 
// vC = 14'b0000000100110111; // vC=  311 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b0000000100011011; // vC=  283 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b0000001000010110; // vC=  534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001000; // iC= 1928 
// vC = 14'b0000001000110100; // vC=  564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000101; // iC= 1861 
// vC = 14'b0000000111011011; // vC=  475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000110; // iC= 1798 
// vC = 14'b0000000100010111; // vC=  279 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011100; // iC= 2076 
// vC = 14'b0000000111100110; // vC=  486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b0000000111000011; // vC=  451 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b0000000101110000; // vC=  368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111000; // iC= 1784 
// vC = 14'b0000000110001010; // vC=  394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010111; // iC= 1815 
// vC = 14'b0000001000111101; // vC=  573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b0000000111010111; // vC=  471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b0000000101001011; // vC=  331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b0000000101011101; // vC=  349 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b0000000101010101; // vC=  341 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b0000000101110010; // vC=  370 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110000; // iC= 1776 
// vC = 14'b0000000110101001; // vC=  425 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b0000001000000011; // vC=  515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b0000000110110110; // vC=  438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011111; // iC= 1759 
// vC = 14'b0000001000011111; // vC=  543 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b0000001000101100; // vC=  556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b0000000110001101; // vC=  397 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000110; // iC= 1798 
// vC = 14'b0000001000011010; // vC=  538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110111; // iC= 2039 
// vC = 14'b0000000111111010; // vC=  506 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b0000001001001010; // vC=  586 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010111; // iC= 1879 
// vC = 14'b0000001001101001; // vC=  617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000001; // iC= 1857 
// vC = 14'b0000001000001111; // vC=  527 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110101; // iC= 1781 
// vC = 14'b0000001001101011; // vC=  619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001100; // iC= 1804 
// vC = 14'b0000001011101101; // vC=  749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010011; // iC= 1875 
// vC = 14'b0000000111110110; // vC=  502 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101101; // iC= 1773 
// vC = 14'b0000001000010001; // vC=  529 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b0000001010100010; // vC=  674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100110; // iC= 1830 
// vC = 14'b0000001000000001; // vC=  513 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010011; // iC= 1747 
// vC = 14'b0000001011001001; // vC=  713 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101010; // iC= 1898 
// vC = 14'b0000001000000111; // vC=  519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b0000001000001010; // vC=  522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101110; // iC= 1838 
// vC = 14'b0000001000100011; // vC=  547 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100111; // iC= 1703 
// vC = 14'b0000001011001101; // vC=  717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011010; // iC= 1818 
// vC = 14'b0000001101001000; // vC=  840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101010; // iC= 1770 
// vC = 14'b0000001001110111; // vC=  631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001101; // iC= 1741 
// vC = 14'b0000001011001010; // vC=  714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001100; // iC= 1676 
// vC = 14'b0000001100011111; // vC=  799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b0000001010110011; // vC=  691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010101; // iC= 1749 
// vC = 14'b0000001001101100; // vC=  620 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100011; // iC= 1955 
// vC = 14'b0000001001001110; // vC=  590 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110011; // iC= 1971 
// vC = 14'b0000001110000110; // vC=  902 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101011; // iC= 1899 
// vC = 14'b0000001100001101; // vC=  781 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101110; // iC= 1966 
// vC = 14'b0000001011000010; // vC=  706 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001000; // iC= 1800 
// vC = 14'b0000001110010110; // vC=  918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101001; // iC= 1833 
// vC = 14'b0000001110000010; // vC=  898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b0000001010011001; // vC=  665 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101100; // iC= 1900 
// vC = 14'b0000001010001011; // vC=  651 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101101; // iC= 1773 
// vC = 14'b0000001010010111; // vC=  663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b0000001101101010; // vC=  874 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100111; // iC= 1639 
// vC = 14'b0000001110001000; // vC=  904 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b0000001110000100; // vC=  900 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010111; // iC= 1687 
// vC = 14'b0000001100001010; // vC=  778 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001011; // iC= 1739 
// vC = 14'b0000001010100011; // vC=  675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110100; // iC= 1780 
// vC = 14'b0000001010111010; // vC=  698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100111; // iC= 1895 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100100; // iC= 1636 
// vC = 14'b0000001011000110; // vC=  710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110101; // iC= 1909 
// vC = 14'b0000001100011100; // vC=  796 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111001; // iC= 1721 
// vC = 14'b0000001011011111; // vC=  735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001010; // iC= 1610 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110110; // iC= 1718 
// vC = 14'b0000001100000001; // vC=  769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011010; // iC= 1818 
// vC = 14'b0000001100000011; // vC=  771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111111; // iC= 1791 
// vC = 14'b0000001101110101; // vC=  885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000110; // iC= 1734 
// vC = 14'b0000001101100001; // vC=  865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000001; // iC= 1601 
// vC = 14'b0000001101001000; // vC=  840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001101; // iC= 1677 
// vC = 14'b0000001110100101; // vC=  933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111010; // iC= 1722 
// vC = 14'b0000001100011101; // vC=  797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000010; // iC= 1666 
// vC = 14'b0000001100010101; // vC=  789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001111; // iC= 1615 
// vC = 14'b0000001111010000; // vC=  976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110001; // iC= 1585 
// vC = 14'b0000010000011000; // vC= 1048 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110011; // iC= 1715 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000110; // iC= 1734 
// vC = 14'b0000010000010100; // vC= 1044 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011010; // iC= 1754 
// vC = 14'b0000001111101101; // vC= 1005 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110011; // iC= 1715 
// vC = 14'b0000001110000010; // vC=  898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000011; // iC= 1603 
// vC = 14'b0000001110001011; // vC=  907 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001001; // iC= 1609 
// vC = 14'b0000001110011100; // vC=  924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101101; // iC= 1645 
// vC = 14'b0000001110111011; // vC=  955 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011101; // iC= 1821 
// vC = 14'b0000010001001011; // vC= 1099 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001101; // iC= 1549 
// vC = 14'b0000001110111100; // vC=  956 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110000; // iC= 1840 
// vC = 14'b0000001110001001; // vC=  905 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b0000010000001000; // vC= 1032 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111101; // iC= 1661 
// vC = 14'b0000010001100100; // vC= 1124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111101; // iC= 1597 
// vC = 14'b0000010000111010; // vC= 1082 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100001; // iC= 1633 
// vC = 14'b0000001111000100; // vC=  964 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001100; // iC= 1548 
// vC = 14'b0000010001111100; // vC= 1148 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010001; // iC= 1681 
// vC = 14'b0000001110101000; // vC=  936 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101001; // iC= 1577 
// vC = 14'b0000010010010100; // vC= 1172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001000; // iC= 1800 
// vC = 14'b0000010000010111; // vC= 1047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011000; // iC= 1752 
// vC = 14'b0000010011010101; // vC= 1237 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000101; // iC= 1733 
// vC = 14'b0000010010110001; // vC= 1201 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000010; // iC= 1730 
// vC = 14'b0000001111010000; // vC=  976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011000; // iC= 1752 
// vC = 14'b0000010010111011; // vC= 1211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100001; // iC= 1569 
// vC = 14'b0000010011001010; // vC= 1226 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111111; // iC= 1471 
// vC = 14'b0000001111111100; // vC= 1020 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111000; // iC= 1464 
// vC = 14'b0000010100000010; // vC= 1282 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100111; // iC= 1703 
// vC = 14'b0000010001111011; // vC= 1147 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110000; // iC= 1456 
// vC = 14'b0000010000101000; // vC= 1064 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001110; // iC= 1678 
// vC = 14'b0000010000000001; // vC= 1025 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111000; // iC= 1528 
// vC = 14'b0000010100011111; // vC= 1311 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010110; // iC= 1686 
// vC = 14'b0000010100101010; // vC= 1322 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101010; // iC= 1514 
// vC = 14'b0000010011001111; // vC= 1231 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001100; // iC= 1548 
// vC = 14'b0000010010000110; // vC= 1158 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100110; // iC= 1574 
// vC = 14'b0000010100011110; // vC= 1310 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011000; // iC= 1432 
// vC = 14'b0000010101000110; // vC= 1350 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111001; // iC= 1657 
// vC = 14'b0000010010111111; // vC= 1215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000100; // iC= 1412 
// vC = 14'b0000010010110000; // vC= 1200 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011010; // iC= 1434 
// vC = 14'b0000010010101100; // vC= 1196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100000; // iC= 1440 
// vC = 14'b0000010010110010; // vC= 1202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101011; // iC= 1579 
// vC = 14'b0000010100010110; // vC= 1302 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011111; // iC= 1695 
// vC = 14'b0000010011011001; // vC= 1241 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011101; // iC= 1693 
// vC = 14'b0000010010110010; // vC= 1202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010001; // iC= 1425 
// vC = 14'b0000010001000111; // vC= 1095 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011001; // iC= 1561 
// vC = 14'b0000010001010100; // vC= 1108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010000; // iC= 1424 
// vC = 14'b0000010010111001; // vC= 1209 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111001; // iC= 1401 
// vC = 14'b0000010101001101; // vC= 1357 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001101; // iC= 1613 
// vC = 14'b0000010010000110; // vC= 1158 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000011; // iC= 1411 
// vC = 14'b0000010101001110; // vC= 1358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110111; // iC= 1655 
// vC = 14'b0000010001111111; // vC= 1151 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001101; // iC= 1485 
// vC = 14'b0000010100001001; // vC= 1289 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100101; // iC= 1573 
// vC = 14'b0000010100110111; // vC= 1335 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100101; // iC= 1445 
// vC = 14'b0000010100101101; // vC= 1325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000010; // iC= 1602 
// vC = 14'b0000010100011011; // vC= 1307 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011001; // iC= 1433 
// vC = 14'b0000010010111110; // vC= 1214 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000000; // iC= 1344 
// vC = 14'b0000010011001111; // vC= 1231 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000011; // iC= 1539 
// vC = 14'b0000010100101110; // vC= 1326 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001000; // iC= 1544 
// vC = 14'b0000010011011010; // vC= 1242 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011011; // iC= 1563 
// vC = 14'b0000010100111000; // vC= 1336 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000100; // iC= 1476 
// vC = 14'b0000010110111111; // vC= 1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001011; // iC= 1611 
// vC = 14'b0000010110110001; // vC= 1457 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010010; // iC= 1490 
// vC = 14'b0000010011110111; // vC= 1271 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110001; // iC= 1585 
// vC = 14'b0000010100100100; // vC= 1316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000100; // iC= 1412 
// vC = 14'b0000010110100100; // vC= 1444 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100100; // iC= 1572 
// vC = 14'b0000010111111011; // vC= 1531 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011110; // iC= 1502 
// vC = 14'b0000010101000001; // vC= 1345 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101000; // iC= 1320 
// vC = 14'b0000010111000101; // vC= 1477 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011011; // iC= 1563 
// vC = 14'b0000010100101100; // vC= 1324 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000100; // iC= 1348 
// vC = 14'b0000010100111101; // vC= 1341 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111011; // iC= 1403 
// vC = 14'b0000010110110101; // vC= 1461 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001000; // iC= 1416 
// vC = 14'b0000010101000101; // vC= 1349 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110101; // iC= 1525 
// vC = 14'b0000010101010100; // vC= 1364 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010011; // iC= 1491 
// vC = 14'b0000010101101011; // vC= 1387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011011; // iC= 1371 
// vC = 14'b0000010111011000; // vC= 1496 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100111; // iC= 1511 
// vC = 14'b0000010100100110; // vC= 1318 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110001; // iC= 1457 
// vC = 14'b0000010110111011; // vC= 1467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110010; // iC= 1522 
// vC = 14'b0000010111110000; // vC= 1520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000100; // iC= 1476 
// vC = 14'b0000010101110011; // vC= 1395 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111011; // iC= 1211 
// vC = 14'b0000010111111100; // vC= 1532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111101; // iC= 1277 
// vC = 14'b0000010111010011; // vC= 1491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001111; // iC= 1423 
// vC = 14'b0000010111110011; // vC= 1523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010001; // iC= 1233 
// vC = 14'b0000010111110011; // vC= 1523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101101; // iC= 1389 
// vC = 14'b0000011000101011; // vC= 1579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110001; // iC= 1265 
// vC = 14'b0000010101011000; // vC= 1368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001111; // iC= 1295 
// vC = 14'b0000010110110101; // vC= 1461 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001010; // iC= 1418 
// vC = 14'b0000011000110010; // vC= 1586 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000011; // iC= 1475 
// vC = 14'b0000010110111000; // vC= 1464 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101011; // iC= 1323 
// vC = 14'b0000010101011101; // vC= 1373 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010111; // iC= 1175 
// vC = 14'b0000010101011000; // vC= 1368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b0000010110001111; // vC= 1423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000110; // iC= 1222 
// vC = 14'b0000010101001010; // vC= 1354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111001; // iC= 1337 
// vC = 14'b0000011000011110; // vC= 1566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101110; // iC= 1390 
// vC = 14'b0000010101111010; // vC= 1402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101010; // iC= 1322 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000011; // iC= 1155 
// vC = 14'b0000011010000001; // vC= 1665 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010001; // iC= 1361 
// vC = 14'b0000011001011110; // vC= 1630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011110; // iC= 1246 
// vC = 14'b0000010111000101; // vC= 1477 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000001; // iC= 1409 
// vC = 14'b0000011000001110; // vC= 1550 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111010; // iC= 1402 
// vC = 14'b0000011000001011; // vC= 1547 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000011; // iC= 1411 
// vC = 14'b0000011000010011; // vC= 1555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110110; // iC= 1142 
// vC = 14'b0000011001000001; // vC= 1601 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110000; // iC= 1328 
// vC = 14'b0000011010110010; // vC= 1714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000111; // iC= 1351 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100011; // iC= 1379 
// vC = 14'b0000011010000010; // vC= 1666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100111; // iC= 1319 
// vC = 14'b0000011011010101; // vC= 1749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011101; // iC= 1373 
// vC = 14'b0000010111100101; // vC= 1509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101101; // iC= 1261 
// vC = 14'b0000010110100111; // vC= 1447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011000; // iC= 1048 
// vC = 14'b0000011000010101; // vC= 1557 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110111; // iC= 1335 
// vC = 14'b0000011010110000; // vC= 1712 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010111; // iC= 1111 
// vC = 14'b0000011010000100; // vC= 1668 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000111; // iC= 1159 
// vC = 14'b0000010110111010; // vC= 1466 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100111; // iC= 1127 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100100; // iC= 1252 
// vC = 14'b0000011010101110; // vC= 1710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111011; // iC= 1019 
// vC = 14'b0000011000010000; // vC= 1552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010001; // iC= 1297 
// vC = 14'b0000011001100010; // vC= 1634 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111000; // iC= 1208 
// vC = 14'b0000011001011000; // vC= 1624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001100; // iC= 1100 
// vC = 14'b0000011011101111; // vC= 1775 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101110; // iC= 1134 
// vC = 14'b0000011000010011; // vC= 1555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001011; // iC= 1163 
// vC = 14'b0000011001001101; // vC= 1613 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001101; // iC= 1037 
// vC = 14'b0000011000001111; // vC= 1551 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001000; // iC= 1288 
// vC = 14'b0000011000001100; // vC= 1548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110100; // iC= 1012 
// vC = 14'b0000011000111100; // vC= 1596 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000001; // iC= 1089 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011110; // iC= 1118 
// vC = 14'b0000011010011001; // vC= 1689 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110101; // iC= 1077 
// vC = 14'b0000011000000100; // vC= 1540 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100011; // iC= 1187 
// vC = 14'b0000011001101101; // vC= 1645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011011; // iC= 1243 
// vC = 14'b0000011100000101; // vC= 1797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000010; // iC=  962 
// vC = 14'b0000011010001001; // vC= 1673 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001010; // iC= 1098 
// vC = 14'b0000011100111100; // vC= 1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000111; // iC= 1031 
// vC = 14'b0000011000110011; // vC= 1587 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110100; // iC= 1140 
// vC = 14'b0000011100101001; // vC= 1833 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111111; // iC= 1215 
// vC = 14'b0000011010001110; // vC= 1678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010000; // iC=  976 
// vC = 14'b0000011101001000; // vC= 1864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011001; // iC= 1177 
// vC = 14'b0000011001100100; // vC= 1636 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100111; // iC=  935 
// vC = 14'b0000011100100011; // vC= 1827 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010110; // iC=  918 
// vC = 14'b0000011001000101; // vC= 1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111001; // iC=  953 
// vC = 14'b0000011001101001; // vC= 1641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000100; // iC=  964 
// vC = 14'b0000011101000010; // vC= 1858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110000; // iC= 1072 
// vC = 14'b0000011100101001; // vC= 1833 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000001; // iC= 1153 
// vC = 14'b0000011010011000; // vC= 1688 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000101; // iC= 1093 
// vC = 14'b0000011100010011; // vC= 1811 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010100; // iC=  980 
// vC = 14'b0000011101100100; // vC= 1892 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010010; // iC=  850 
// vC = 14'b0000011010111000; // vC= 1720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110010; // iC= 1138 
// vC = 14'b0000011010001000; // vC= 1672 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110010; // iC=  946 
// vC = 14'b0000011010101010; // vC= 1706 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000010; // iC= 1090 
// vC = 14'b0000011010100001; // vC= 1697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100011; // iC=  995 
// vC = 14'b0000011011000011; // vC= 1731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011000; // iC= 1048 
// vC = 14'b0000011100000111; // vC= 1799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011010; // iC=  858 
// vC = 14'b0000011001010010; // vC= 1618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100100; // iC=  804 
// vC = 14'b0000011011100001; // vC= 1761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011110; // iC=  990 
// vC = 14'b0000011011010111; // vC= 1751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001011; // iC= 1099 
// vC = 14'b0000011100001101; // vC= 1805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001001; // iC= 1097 
// vC = 14'b0000011100110000; // vC= 1840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110110; // iC=  822 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111001; // iC=  953 
// vC = 14'b0000011110001001; // vC= 1929 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001001; // iC=  777 
// vC = 14'b0000011100011100; // vC= 1820 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001000; // iC=  904 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101011; // iC= 1067 
// vC = 14'b0000011110111000; // vC= 1976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011100; // iC=  860 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011100; // iC=  732 
// vC = 14'b0000011100000110; // vC= 1798 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011110; // iC=  734 
// vC = 14'b0000011100111101; // vC= 1853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000001; // iC=  833 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100111; // iC=  807 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001000; // iC=  840 
// vC = 14'b0000011011110011; // vC= 1779 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001111; // iC=  911 
// vC = 14'b0000011101001101; // vC= 1869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001000; // iC=  840 
// vC = 14'b0000011111001000; // vC= 1992 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100001; // iC=  801 
// vC = 14'b0000011100111110; // vC= 1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111011; // iC=  891 
// vC = 14'b0000011010010111; // vC= 1687 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101101; // iC=  813 
// vC = 14'b0000011111010100; // vC= 2004 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011001; // iC=  921 
// vC = 14'b0000011110001111; // vC= 1935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011111; // iC=  799 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101001; // iC=  809 
// vC = 14'b0000011101101111; // vC= 1903 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110001; // iC=  689 
// vC = 14'b0000011101111111; // vC= 1919 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111011; // iC=  955 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110100; // iC=  820 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001000; // iC=  904 
// vC = 14'b0000011111000111; // vC= 1991 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110001; // iC=  753 
// vC = 14'b0000011100100111; // vC= 1831 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110001; // iC=  817 
// vC = 14'b0000011111110100; // vC= 2036 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110110; // iC=  822 
// vC = 14'b0000011101001101; // vC= 1869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100101; // iC=  613 
// vC = 14'b0000011111111101; // vC= 2045 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000011; // iC=  771 
// vC = 14'b0000011110001011; // vC= 1931 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000110; // iC=  710 
// vC = 14'b0000011101101001; // vC= 1897 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110100; // iC=  820 
// vC = 14'b0000011110011000; // vC= 1944 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001100; // iC=  780 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101011; // iC=  683 
// vC = 14'b0000011110010001; // vC= 1937 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110011; // iC=  627 
// vC = 14'b0000011100010101; // vC= 1813 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100111; // iC=  807 
// vC = 14'b0000011011100110; // vC= 1766 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100001; // iC=  801 
// vC = 14'b0000011100010110; // vC= 1814 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000000; // iC=  576 
// vC = 14'b0000011111100011; // vC= 2019 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010001; // iC=  721 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110101; // iC=  757 
// vC = 14'b0000011100111000; // vC= 1848 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010010; // iC=  658 
// vC = 14'b0000100000000010; // vC= 2050 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000010; // iC=  642 
// vC = 14'b0000011101000101; // vC= 1861 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000011; // iC=  579 
// vC = 14'b0000100000100101; // vC= 2085 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000010; // iC=  706 
// vC = 14'b0000011110010010; // vC= 1938 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100110; // iC=  678 
// vC = 14'b0000100000011001; // vC= 2073 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101010; // iC=  554 
// vC = 14'b0000011111111010; // vC= 2042 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100111; // iC=  807 
// vC = 14'b0000011110100101; // vC= 1957 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001010; // iC=  714 
// vC = 14'b0000011100000111; // vC= 1799 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111011; // iC=  699 
// vC = 14'b0000100000010011; // vC= 2067 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101100; // iC=  620 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010100; // iC=  660 
// vC = 14'b0000011101111011; // vC= 1915 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010001; // iC=  721 
// vC = 14'b0000011100010001; // vC= 1809 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001100; // iC=  460 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010100; // iC=  660 
// vC = 14'b0000011110001101; // vC= 1933 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011010; // iC=  410 
// vC = 14'b0000011100010111; // vC= 1815 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111100; // iC=  700 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010100; // iC=  596 
// vC = 14'b0000011111010100; // vC= 2004 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000110; // iC=  582 
// vC = 14'b0000011111101001; // vC= 2025 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100100; // iC=  356 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001011; // iC=  331 
// vC = 14'b0000011101111110; // vC= 1918 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110110; // iC=  374 
// vC = 14'b0000100000000111; // vC= 2055 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100100; // iC=  420 
// vC = 14'b0000011111000001; // vC= 1985 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011101; // iC=  477 
// vC = 14'b0000011111010110; // vC= 2006 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110001; // iC=  305 
// vC = 14'b0000011111101001; // vC= 2025 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000101; // iC=  325 
// vC = 14'b0000011110011001; // vC= 1945 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010100; // iC=  276 
// vC = 14'b0000011100010001; // vC= 1809 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110101; // iC=  373 
// vC = 14'b0000011101010001; // vC= 1873 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111000; // iC=  376 
// vC = 14'b0000100000100100; // vC= 2084 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100010; // iC=  418 
// vC = 14'b0000100001001101; // vC= 2125 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101111; // iC=  495 
// vC = 14'b0000011110111001; // vC= 1977 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100110; // iC=  294 
// vC = 14'b0000011100110011; // vC= 1843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011110; // iC=  350 
// vC = 14'b0000011110111010; // vC= 1978 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111100; // iC=  188 
// vC = 14'b0000011101111001; // vC= 1913 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011111; // iC=  159 
// vC = 14'b0000011101001111; // vC= 1871 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010111; // iC=  279 
// vC = 14'b0000011110101011; // vC= 1963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110101; // iC=  245 
// vC = 14'b0000011100011011; // vC= 1819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111100; // iC=  124 
// vC = 14'b0000100000001001; // vC= 2057 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001100; // iC=   76 
// vC = 14'b0000011111110100; // vC= 2036 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100111; // iC=  167 
// vC = 14'b0000011110100011; // vC= 1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100101; // iC=  101 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001001; // iC=  137 
// vC = 14'b0000011111010001; // vC= 2001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100110; // iC=  166 
// vC = 14'b0000011110111010; // vC= 1978 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101111; // iC=  -17 
// vC = 14'b0000011100100100; // vC= 1828 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101110; // iC=   46 
// vC = 14'b0000100000110000; // vC= 2096 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001010; // iC=  138 
// vC = 14'b0000011110001011; // vC= 1931 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010010; // iC=  -46 
// vC = 14'b0000100000100111; // vC= 2087 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111010; // iC=   -6 
// vC = 14'b0000011111010000; // vC= 2000 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011110; // iC=   94 
// vC = 14'b0000011100110000; // vC= 1840 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101110111; // iC= -137 
// vC = 14'b0000011101101010; // vC= 1898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100101; // iC=  -91 
// vC = 14'b0000011100111011; // vC= 1851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101000; // iC=  -24 
// vC = 14'b0000011110111001; // vC= 1977 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001010; // iC=   10 
// vC = 14'b0000100000111000; // vC= 2104 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100101; // iC=  -91 
// vC = 14'b0000011110100100; // vC= 1956 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010100; // iC= -236 
// vC = 14'b0000011111110111; // vC= 2039 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011100; // iC= -100 
// vC = 14'b0000011100100100; // vC= 1828 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111110101; // iC=  -11 
// vC = 14'b0000011101000000; // vC= 1856 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110110010; // iC=  -78 
// vC = 14'b0000011111010101; // vC= 2005 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000000; // iC= -256 
// vC = 14'b0000011111101100; // vC= 2028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001100; // iC= -308 
// vC = 14'b0000100000100100; // vC= 2084 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101000; // iC= -216 
// vC = 14'b0000011101101110; // vC= 1902 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110100; // iC= -396 
// vC = 14'b0000011100110101; // vC= 1845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111000; // iC= -392 
// vC = 14'b0000100000010011; // vC= 2067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100101; // iC= -219 
// vC = 14'b0000011111111111; // vC= 2047 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011010; // iC= -422 
// vC = 14'b0000011110001111; // vC= 1935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001100; // iC= -436 
// vC = 14'b0000011110100110; // vC= 1958 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101110; // iC= -466 
// vC = 14'b0000011110111100; // vC= 1980 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011010; // iC= -358 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110110; // iC= -394 
// vC = 14'b0000011111100011; // vC= 2019 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011101; // iC= -291 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010001; // iC= -367 
// vC = 14'b0000100000100111; // vC= 2087 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110011; // iC= -461 
// vC = 14'b0000011110100101; // vC= 1957 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000111; // iC= -633 
// vC = 14'b0000011110001111; // vC= 1935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100000; // iC= -416 
// vC = 14'b0000011110010001; // vC= 1937 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101111; // iC= -593 
// vC = 14'b0000011111000001; // vC= 1985 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001010; // iC= -694 
// vC = 14'b0000011100010111; // vC= 1815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100110; // iC= -666 
// vC = 14'b0000011100001010; // vC= 1802 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100100; // iC= -732 
// vC = 14'b0000011100001100; // vC= 1804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110110; // iC= -586 
// vC = 14'b0000011111001010; // vC= 1994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111110010; // iC= -526 
// vC = 14'b0000011111010111; // vC= 2007 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010100; // iC= -556 
// vC = 14'b0000011101001001; // vC= 1865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011111; // iC= -801 
// vC = 14'b0000011101101101; // vC= 1901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101011; // iC= -917 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010111; // iC= -617 
// vC = 14'b0000100000001011; // vC= 2059 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001111; // iC= -945 
// vC = 14'b0000011111100000; // vC= 2016 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101001; // iC= -983 
// vC = 14'b0000100000010010; // vC= 2066 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100100; // iC= -860 
// vC = 14'b0000011111000111; // vC= 1991 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001110; // iC= -946 
// vC = 14'b0000011101011001; // vC= 1881 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000010; // iC= -766 
// vC = 14'b0000011110000011; // vC= 1923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111011; // iC= -837 
// vC = 14'b0000011100101101; // vC= 1837 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111101; // iC= -835 
// vC = 14'b0000011100001011; // vC= 1803 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100111; // iC=-1049 
// vC = 14'b0000011111010000; // vC= 2000 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000101; // iC= -955 
// vC = 14'b0000011011010100; // vC= 1748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101001; // iC=-1047 
// vC = 14'b0000011011000101; // vC= 1733 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101111; // iC=-1105 
// vC = 14'b0000011101100111; // vC= 1895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110100; // iC= -908 
// vC = 14'b0000011111001000; // vC= 1992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101000; // iC=-1048 
// vC = 14'b0000011100010110; // vC= 1814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110010; // iC=-1230 
// vC = 14'b0000011011010101; // vC= 1749 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110011; // iC=-1165 
// vC = 14'b0000011110010011; // vC= 1939 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110111; // iC=-1225 
// vC = 14'b0000011010101111; // vC= 1711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111100; // iC=-1284 
// vC = 14'b0000011110110001; // vC= 1969 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110010; // iC=-1038 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111001; // iC=-1287 
// vC = 14'b0000011111001000; // vC= 1992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010100; // iC=-1324 
// vC = 14'b0000011010111110; // vC= 1726 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111010; // iC=-1158 
// vC = 14'b0000011011101101; // vC= 1773 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011110; // iC=-1314 
// vC = 14'b0000011110101000; // vC= 1960 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101010; // iC=-1174 
// vC = 14'b0000011001111000; // vC= 1656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111110; // iC=-1282 
// vC = 14'b0000011100101010; // vC= 1834 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100100; // iC=-1436 
// vC = 14'b0000011110010010; // vC= 1938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111111; // iC=-1345 
// vC = 14'b0000011100110100; // vC= 1844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010000; // iC=-1264 
// vC = 14'b0000011010000011; // vC= 1667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100011; // iC=-1373 
// vC = 14'b0000011001101001; // vC= 1641 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000101; // iC=-1211 
// vC = 14'b0000011110001111; // vC= 1935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011100; // iC=-1316 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000011; // iC=-1341 
// vC = 14'b0000011100110011; // vC= 1843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011100; // iC=-1572 
// vC = 14'b0000011001001001; // vC= 1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100010; // iC=-1566 
// vC = 14'b0000011001110000; // vC= 1648 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000010; // iC=-1342 
// vC = 14'b0000011101011000; // vC= 1880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000011; // iC=-1533 
// vC = 14'b0000011100000101; // vC= 1797 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000101; // iC=-1339 
// vC = 14'b0000011101000001; // vC= 1857 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100001; // iC=-1631 
// vC = 14'b0000011001001100; // vC= 1612 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010110; // iC=-1514 
// vC = 14'b0000011101000111; // vC= 1863 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101011; // iC=-1685 
// vC = 14'b0000011000011101; // vC= 1565 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001100; // iC=-1396 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001101; // iC=-1587 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000000; // iC=-1600 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100101; // iC=-1691 
// vC = 14'b0000011010101110; // vC= 1710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000011; // iC=-1597 
// vC = 14'b0000011001111111; // vC= 1663 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111110; // iC=-1602 
// vC = 14'b0000011010111011; // vC= 1723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111110; // iC=-1730 
// vC = 14'b0000011010111110; // vC= 1726 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110100; // iC=-1484 
// vC = 14'b0000011010110011; // vC= 1715 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100001; // iC=-1695 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100000; // iC=-1824 
// vC = 14'b0000011001110001; // vC= 1649 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110110; // iC=-1610 
// vC = 14'b0000011000101000; // vC= 1576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111001; // iC=-1735 
// vC = 14'b0000011010110001; // vC= 1713 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110011; // iC=-1677 
// vC = 14'b0000010111101001; // vC= 1513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b0000011010011011; // vC= 1691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110111; // iC=-1673 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b0000011010001010; // vC= 1674 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011001; // iC=-1639 
// vC = 14'b0000011000101000; // vC= 1576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100110; // iC=-1818 
// vC = 14'b0000011001100100; // vC= 1636 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b0000010111001110; // vC= 1486 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101111; // iC=-1681 
// vC = 14'b0000011001111101; // vC= 1661 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100010; // iC=-1694 
// vC = 14'b0000011001010001; // vC= 1617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110001; // iC=-1743 
// vC = 14'b0000010111000100; // vC= 1476 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b0000011010000001; // vC= 1665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111101; // iC=-1859 
// vC = 14'b0000011001100001; // vC= 1633 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001011; // iC=-1973 
// vC = 14'b0000011000110101; // vC= 1589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000100; // iC=-1788 
// vC = 14'b0000010111000111; // vC= 1479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110000; // iC=-2000 
// vC = 14'b0000010101011100; // vC= 1372 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011001; // iC=-1831 
// vC = 14'b0000010110000110; // vC= 1414 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110001; // iC=-1935 
// vC = 14'b0000010111011110; // vC= 1502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100011; // iC=-1949 
// vC = 14'b0000011001010111; // vC= 1623 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b0000011000100010; // vC= 1570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b0000010111010100; // vC= 1492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000010101101000; // vC= 1384 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000010100000011; // vC= 1283 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000100; // iC=-1916 
// vC = 14'b0000011000101101; // vC= 1581 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110010; // iC=-1998 
// vC = 14'b0000010111011001; // vC= 1497 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100001; // iC=-2079 
// vC = 14'b0000010111101000; // vC= 1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010100; // iC=-1900 
// vC = 14'b0000010110100011; // vC= 1443 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b0000010100110001; // vC= 1329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001101; // iC=-2099 
// vC = 14'b0000010111110111; // vC= 1527 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b0000010111001110; // vC= 1486 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b0000010110010011; // vC= 1427 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100100; // iC=-1820 
// vC = 14'b0000010011001111; // vC= 1231 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110010; // iC=-1998 
// vC = 14'b0000010111010001; // vC= 1489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111111; // iC=-2113 
// vC = 14'b0000010101100010; // vC= 1378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b0000010101011110; // vC= 1374 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b0000010011001001; // vC= 1225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000010; // iC=-2046 
// vC = 14'b0000010001110001; // vC= 1137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110001; // iC=-1999 
// vC = 14'b0000010100010110; // vC= 1302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b0000010010110100; // vC= 1204 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011101; // iC=-1827 
// vC = 14'b0000010101010010; // vC= 1362 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100111; // iC=-2073 
// vC = 14'b0000010100010111; // vC= 1303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b0000010001011010; // vC= 1114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010011; // iC=-2093 
// vC = 14'b0000010001101011; // vC= 1131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010110; // iC=-2154 
// vC = 14'b0000010101010110; // vC= 1366 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100100; // iC=-1948 
// vC = 14'b0000010010111001; // vC= 1209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b0000010010001010; // vC= 1162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b0000010011111010; // vC= 1274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b0000010001111010; // vC= 1146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110001; // iC=-2127 
// vC = 14'b0000010010001010; // vC= 1162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100000; // iC=-2016 
// vC = 14'b0000010000100100; // vC= 1060 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b0000010011110001; // vC= 1265 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100100; // iC=-1948 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111101; // iC=-1923 
// vC = 14'b0000010011100001; // vC= 1249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000010011111111; // vC= 1279 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b0000001111100111; // vC=  999 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000010010111010; // vC= 1210 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010110; // iC=-2154 
// vC = 14'b0000001111110011; // vC= 1011 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101011; // iC=-2069 
// vC = 14'b0000001111000001; // vC=  961 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001101; // iC=-2099 
// vC = 14'b0000001111101111; // vC= 1007 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b0000010001100001; // vC= 1121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110010; // iC=-2190 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110000; // iC=-2128 
// vC = 14'b0000010000001010; // vC= 1034 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b0000010001111110; // vC= 1150 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b0000010010011000; // vC= 1176 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110100; // iC=-2060 
// vC = 14'b0000010001110110; // vC= 1142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001001; // iC=-2103 
// vC = 14'b0000010000001101; // vC= 1037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101010; // iC=-2134 
// vC = 14'b0000010001010100; // vC= 1108 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b0000001110001001; // vC=  905 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011111; // iC=-2209 
// vC = 14'b0000010001111011; // vC= 1147 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101011; // iC=-2069 
// vC = 14'b0000001111101001; // vC= 1001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110010; // iC=-2126 
// vC = 14'b0000001101101001; // vC=  873 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b0000001110110111; // vC=  951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111111; // iC=-2113 
// vC = 14'b0000001101000111; // vC=  839 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000101; // iC=-2171 
// vC = 14'b0000001101000100; // vC=  836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110011; // iC=-1997 
// vC = 14'b0000010000011001; // vC= 1049 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b0000010000100011; // vC= 1059 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b0000001101110101; // vC=  885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b0000010000110010; // vC= 1074 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011110; // iC=-2146 
// vC = 14'b0000001111111001; // vC= 1017 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001000; // iC=-2168 
// vC = 14'b0000001110111001; // vC=  953 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111001; // iC=-1927 
// vC = 14'b0000001110111011; // vC=  955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100101; // iC=-2203 
// vC = 14'b0000001100000010; // vC=  770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b0000001101110101; // vC=  885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110001; // iC=-2063 
// vC = 14'b0000001101111010; // vC=  890 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b0000001111001011; // vC=  971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111100; // iC=-2180 
// vC = 14'b0000001011000110; // vC=  710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b0000001101001111; // vC=  847 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b0000001100101000; // vC=  808 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000001; // iC=-1919 
// vC = 14'b0000001100011011; // vC=  795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000001101100100; // vC=  868 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111011; // iC=-2181 
// vC = 14'b0000001101101100; // vC=  876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000001011000111; // vC=  711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000001101100011; // vC=  867 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b0000001100000110; // vC=  774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100000; // iC=-2208 
// vC = 14'b0000001010010101; // vC=  661 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b0000001110000000; // vC=  896 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010010; // iC=-1966 
// vC = 14'b0000001010011000; // vC=  664 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001000; // iC=-2040 
// vC = 14'b0000001100100000; // vC=  800 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110010; // iC=-2126 
// vC = 14'b0000001101000111; // vC=  839 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110101; // iC=-2187 
// vC = 14'b0000001001000100; // vC=  580 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000001; // iC=-1919 
// vC = 14'b0000001010011001; // vC=  665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101000; // iC=-2200 
// vC = 14'b0000001010110101; // vC=  693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b0000001010111011; // vC=  699 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110010; // iC=-2190 
// vC = 14'b0000001100000000; // vC=  768 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b0000001101001101; // vC=  845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b0000001100011111; // vC=  799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b0000001001010111; // vC=  599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b0000001000110011; // vC=  563 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001000; // iC=-2040 
// vC = 14'b0000001100010110; // vC=  790 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b0000001001111010; // vC=  634 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b0000001001000111; // vC=  583 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000001001100101; // vC=  613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b0000001000011111; // vC=  543 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100001; // iC=-2143 
// vC = 14'b0000000111011100; // vC=  476 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001011; // iC=-2229 
// vC = 14'b0000000111001111; // vC=  463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000100; // iC=-2236 
// vC = 14'b0000001000011000; // vC=  536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101001; // iC=-2135 
// vC = 14'b0000001011001010; // vC=  714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000111; // iC=-1977 
// vC = 14'b0000001000001110; // vC=  526 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001000; // iC=-2168 
// vC = 14'b0000001010110110; // vC=  694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011110; // iC=-2146 
// vC = 14'b0000001000011000; // vC=  536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011001; // iC=-2151 
// vC = 14'b0000001001001100; // vC=  588 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111100; // iC=-1988 
// vC = 14'b0000001000111010; // vC=  570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011100; // iC=-2148 
// vC = 14'b0000000110110000; // vC=  432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010100; // iC=-2092 
// vC = 14'b0000000110111001; // vC=  441 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000011; // iC=-2237 
// vC = 14'b0000001010010101; // vC=  661 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000000110111011; // vC=  443 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010011; // iC=-2221 
// vC = 14'b0000001001001000; // vC=  584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110000; // iC=-2064 
// vC = 14'b0000001001001100; // vC=  588 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000111; // iC=-2169 
// vC = 14'b0000001000000111; // vC=  519 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100101; // iC=-2203 
// vC = 14'b0000000101001001; // vC=  329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111001; // iC=-1991 
// vC = 14'b0000000110100010; // vC=  418 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001011; // iC=-2165 
// vC = 14'b0000000111110110; // vC=  502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b0000000100001110; // vC=  270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000001000011000; // vC=  536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b0000000100101010; // vC=  298 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010101; // iC=-2027 
// vC = 14'b0000000111010111; // vC=  471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b0000000011111111; // vC=  255 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110100; // iC=-2124 
// vC = 14'b0000001000100001; // vC=  545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011001; // iC=-2087 
// vC = 14'b0000000111110010; // vC=  498 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b0000000011101111; // vC=  239 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011111; // iC=-2209 
// vC = 14'b0000000111011000; // vC=  472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000000111111111; // vC=  511 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b0000000011000111; // vC=  199 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111000; // iC=-1928 
// vC = 14'b0000000110001100; // vC=  396 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000000011100001; // vC=  225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010111; // iC=-2217 
// vC = 14'b0000000011111110; // vC=  254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b0000000111010011; // vC=  467 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b0000000011000011; // vC=  195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000000110000101; // vC=  389 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010111; // iC=-2089 
// vC = 14'b0000000010111110; // vC=  190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011011; // iC=-2149 
// vC = 14'b0000000101110011; // vC=  371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000000100001100; // vC=  268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001111; // iC=-2161 
// vC = 14'b0000000100100011; // vC=  291 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111000; // iC=-1928 
// vC = 14'b0000000110010011; // vC=  403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b0000000011000110; // vC=  198 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b0000000011111011; // vC=  251 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011110; // iC=-2018 
// vC = 14'b0000000010101001; // vC=  169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b0000000100001011; // vC=  267 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000111; // iC=-2169 
// vC = 14'b0000000100101110; // vC=  302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b0000000001010011; // vC=   83 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001101; // iC=-2227 
// vC = 14'b0000000001010011; // vC=   83 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111100; // iC=-1924 
// vC = 14'b0000000010101001; // vC=  169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100000; // iC=-2016 
// vC = 14'b0000000100110000; // vC=  304 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000010; // iC=-2046 
// vC = 14'b0000000100111000; // vC=  312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011111; // iC=-2209 
// vC = 14'b0000000010100010; // vC=  162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b0000000010000011; // vC=  131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000000001000011; // vC=   67 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010101; // iC=-2027 
// vC = 14'b0000000010101110; // vC=  174 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b0000000000100110; // vC=   38 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100110; // iC=-2138 
// vC = 14'b0000000001000110; // vC=   70 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b1111111111111111; // vC=   -1 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101111; // iC=-2193 
// vC = 14'b0000000010100011; // vC=  163 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000000001010111; // vC=   87 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011101; // iC=-2211 
// vC = 14'b0000000000101000; // vC=   40 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b1111111111001000; // vC=  -56 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b1111111110101111; // vC=  -81 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b1111111111010101; // vC=  -43 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b1111111111010100; // vC=  -44 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111110; // iC=-1922 
// vC = 14'b1111111111101100; // vC=  -20 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b1111111110111001; // vC=  -71 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010000; // iC=-2160 
// vC = 14'b0000000001111001; // vC=  121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b1111111101110011; // vC= -141 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111010; // iC=-2182 
// vC = 14'b1111111101101100; // vC= -148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010010; // iC=-1966 
// vC = 14'b0000000000011111; // vC=   31 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011000; // iC=-2024 
// vC = 14'b0000000001100010; // vC=   98 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b1111111101001011; // vC= -181 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011000; // iC=-2088 
// vC = 14'b1111111100111101; // vC= -195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010000; // iC=-2160 
// vC = 14'b1111111111000010; // vC=  -62 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b1111111100101110; // vC= -210 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b1111111111101001; // vC=  -23 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b1111111110101101; // vC=  -83 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000010; // iC=-2174 
// vC = 14'b1111111110101110; // vC=  -82 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b1111111100001010; // vC= -246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b1111111111000110; // vC=  -58 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111100; // iC=-2180 
// vC = 14'b1111111100100111; // vC= -217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101010; // iC=-2070 
// vC = 14'b1111111110111110; // vC=  -66 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b1111111100101011; // vC= -213 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b1111111100110110; // vC= -202 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110011; // iC=-1933 
// vC = 14'b1111111111000101; // vC=  -59 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b1111111110001000; // vC= -120 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b1111111110011100; // vC= -100 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010100; // iC=-2028 
// vC = 14'b1111111110010011; // vC= -109 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011001; // iC=-2087 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b1111111101001010; // vC= -182 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011001; // iC=-1895 
// vC = 14'b1111111110000010; // vC= -126 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010000; // iC=-1968 
// vC = 14'b1111111110111001; // vC=  -71 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100101; // iC=-2139 
// vC = 14'b1111111001110101; // vC= -395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000001; // iC=-1855 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111100; // iC=-1860 
// vC = 14'b1111111010101101; // vC= -339 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100001; // iC=-2079 
// vC = 14'b1111111110011111; // vC=  -97 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b1111111011101010; // vC= -278 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011111; // iC=-2081 
// vC = 14'b1111111100111000; // vC= -200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b1111111101110100; // vC= -140 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b1111111010011010; // vC= -358 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111111010110010; // vC= -334 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111100; // iC=-1860 
// vC = 14'b1111111001000101; // vC= -443 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b1111111001100100; // vC= -412 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111100; // iC=-1924 
// vC = 14'b1111111001010000; // vC= -432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b1111111000100001; // vC= -479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101001; // iC=-2071 
// vC = 14'b1111111100111111; // vC= -193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010111; // iC=-2089 
// vC = 14'b1111111001010000; // vC= -432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010000; // iC=-1968 
// vC = 14'b1111111001010011; // vC= -429 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b1111111010110100; // vC= -332 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100101; // iC=-1819 
// vC = 14'b1111111001000001; // vC= -447 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b1111111011010111; // vC= -297 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b1111111011100100; // vC= -284 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b1111111000110100; // vC= -460 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111111; // iC=-1921 
// vC = 14'b1111111011011111; // vC= -289 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111100; // iC=-1860 
// vC = 14'b1111111001110111; // vC= -393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000000; // iC=-1856 
// vC = 14'b1111111010010010; // vC= -366 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110111; // iC=-1865 
// vC = 14'b1111111010010010; // vC= -366 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b1111111011010101; // vC= -299 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010001; // iC=-2031 
// vC = 14'b1111111001110011; // vC= -397 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b1111111000010111; // vC= -489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110010; // iC=-2062 
// vC = 14'b1111111001100111; // vC= -409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b1111110111001001; // vC= -567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010111; // iC=-1769 
// vC = 14'b1111110110011101; // vC= -611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b1111111001101111; // vC= -401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b1111111001010110; // vC= -426 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110000; // iC=-1808 
// vC = 14'b1111111000111000; // vC= -456 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000101; // iC=-2043 
// vC = 14'b1111110111010001; // vC= -559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011110; // iC=-1826 
// vC = 14'b1111110111100001; // vC= -543 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000100; // iC=-1852 
// vC = 14'b1111110110010110; // vC= -618 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b1111110101011011; // vC= -677 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b1111110110001100; // vC= -628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b1111110110011001; // vC= -615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110010; // iC=-1934 
// vC = 14'b1111110111110011; // vC= -525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101011; // iC=-1749 
// vC = 14'b1111110100011011; // vC= -741 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b1111110100100010; // vC= -734 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b1111110111101011; // vC= -533 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b1111110101101100; // vC= -660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b1111110111110000; // vC= -528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b1111110110100111; // vC= -601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b1111110100111100; // vC= -708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b1111110011110110; // vC= -778 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b1111110100101010; // vC= -726 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b1111110111110011; // vC= -525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b1111110111000111; // vC= -569 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110011; // iC=-1869 
// vC = 14'b1111111000000011; // vC= -509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010101; // iC=-1707 
// vC = 14'b1111110101011001; // vC= -679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011001; // iC=-1767 
// vC = 14'b1111110111010011; // vC= -557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110001; // iC=-1743 
// vC = 14'b1111110010111100; // vC= -836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011101; // iC=-1699 
// vC = 14'b1111110101110001; // vC= -655 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111000; // iC=-1928 
// vC = 14'b1111110101110000; // vC= -656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b1111110011000011; // vC= -829 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000100; // iC=-1916 
// vC = 14'b1111110100100110; // vC= -730 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b1111110100011100; // vC= -740 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001110; // iC=-1842 
// vC = 14'b1111110100010100; // vC= -748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001110; // iC=-1714 
// vC = 14'b1111110101000010; // vC= -702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b1111110100111001; // vC= -711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b1111110001111001; // vC= -903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b1111110010000000; // vC= -896 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100100; // iC=-1948 
// vC = 14'b1111110010100011; // vC= -861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110010; // iC=-1806 
// vC = 14'b1111110011000001; // vC= -831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110011; // iC=-1677 
// vC = 14'b1111110100111010; // vC= -710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001000; // iC=-1720 
// vC = 14'b1111110011100111; // vC= -793 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001011; // iC=-1781 
// vC = 14'b1111110010011100; // vC= -868 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110111; // iC=-1673 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110010; // iC=-1678 
// vC = 14'b1111110010011011; // vC= -869 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b1111110010001110; // vC= -882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110010; // iC=-1870 
// vC = 14'b1111110011010000; // vC= -816 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b1111110011001010; // vC= -822 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b1111110100110101; // vC= -715 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b1111110100001111; // vC= -753 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101010; // iC=-1750 
// vC = 14'b1111110000101011; // vC= -981 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111110010010010; // vC= -878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111010; // iC=-1734 
// vC = 14'b1111110000111000; // vC= -968 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111110; // iC=-1602 
// vC = 14'b1111110000100101; // vC= -987 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000101; // iC=-1723 
// vC = 14'b1111110000101100; // vC= -980 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111000; // iC=-1800 
// vC = 14'b1111110001111011; // vC= -901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101110; // iC=-1746 
// vC = 14'b1111110001011110; // vC= -930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111101; // iC=-1859 
// vC = 14'b1111110000111001; // vC= -967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000100; // iC=-1788 
// vC = 14'b1111101111110110; // vC=-1034 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001110; // iC=-1842 
// vC = 14'b1111110001001001; // vC= -951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010000; // iC=-1776 
// vC = 14'b1111110001000101; // vC= -955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001001; // iC=-1847 
// vC = 14'b1111110010101111; // vC= -849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010000; // iC=-1584 
// vC = 14'b1111110011001101; // vC= -819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101101; // iC=-1683 
// vC = 14'b1111101110101000; // vC=-1112 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001001; // iC=-1783 
// vC = 14'b1111101110111000; // vC=-1096 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110100; // iC=-1740 
// vC = 14'b1111110001011010; // vC= -934 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011011; // iC=-1701 
// vC = 14'b1111101110000011; // vC=-1149 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011111; // iC=-1569 
// vC = 14'b1111101110110000; // vC=-1104 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011111; // iC=-1697 
// vC = 14'b1111110001011001; // vC= -935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101111; // iC=-1553 
// vC = 14'b1111110001111011; // vC= -901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111011; // iC=-1541 
// vC = 14'b1111110010001000; // vC= -888 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000001; // iC=-1535 
// vC = 14'b1111101110101100; // vC=-1108 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110001; // iC=-1551 
// vC = 14'b1111101101101100; // vC=-1172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110110; // iC=-1674 
// vC = 14'b1111110000110010; // vC= -974 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101101; // iC=-1619 
// vC = 14'b1111110000000001; // vC=-1023 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011011; // iC=-1573 
// vC = 14'b1111101110001101; // vC=-1139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011010; // iC=-1510 
// vC = 14'b1111101110011110; // vC=-1122 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000110; // iC=-1722 
// vC = 14'b1111101101100101; // vC=-1179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111111; // iC=-1601 
// vC = 14'b1111101111110111; // vC=-1033 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001101; // iC=-1779 
// vC = 14'b1111101101001101; // vC=-1203 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100101; // iC=-1691 
// vC = 14'b1111101101001111; // vC=-1201 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111110; // iC=-1794 
// vC = 14'b1111101111000111; // vC=-1081 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111110; // iC=-1730 
// vC = 14'b1111110000010100; // vC=-1004 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100000; // iC=-1504 
// vC = 14'b1111101110001111; // vC=-1137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001111; // iC=-1521 
// vC = 14'b1111101111110110; // vC=-1034 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111000; // iC=-1672 
// vC = 14'b1111101100100010; // vC=-1246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000001; // iC=-1471 
// vC = 14'b1111101110001010; // vC=-1142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000000; // iC=-1728 
// vC = 14'b1111101011111101; // vC=-1283 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000011; // iC=-1661 
// vC = 14'b1111101011101000; // vC=-1304 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101001; // iC=-1495 
// vC = 14'b1111101101010000; // vC=-1200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000101; // iC=-1595 
// vC = 14'b1111101100000101; // vC=-1275 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100111; // iC=-1753 
// vC = 14'b1111101011100111; // vC=-1305 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010110; // iC=-1514 
// vC = 14'b1111101100111110; // vC=-1218 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111001; // iC=-1735 
// vC = 14'b1111101111000011; // vC=-1085 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011111; // iC=-1697 
// vC = 14'b1111101011011101; // vC=-1315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100001; // iC=-1695 
// vC = 14'b1111101110110001; // vC=-1103 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001010; // iC=-1590 
// vC = 14'b1111101110100000; // vC=-1120 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011110; // iC=-1442 
// vC = 14'b1111101111110000; // vC=-1040 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011111; // iC=-1505 
// vC = 14'b1111101110000101; // vC=-1147 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010100; // iC=-1580 
// vC = 14'b1111101100101110; // vC=-1234 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111011; // iC=-1605 
// vC = 14'b1111101101000110; // vC=-1210 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001000; // iC=-1656 
// vC = 14'b1111101011101010; // vC=-1302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100111; // iC=-1497 
// vC = 14'b1111101011100111; // vC=-1305 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111001; // iC=-1479 
// vC = 14'b1111101101000100; // vC=-1212 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011111; // iC=-1697 
// vC = 14'b1111101110010000; // vC=-1136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001101; // iC=-1651 
// vC = 14'b1111101010110110; // vC=-1354 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010010; // iC=-1390 
// vC = 14'b1111101001111000; // vC=-1416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100010; // iC=-1502 
// vC = 14'b1111101011001100; // vC=-1332 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111100; // iC=-1476 
// vC = 14'b1111101010110000; // vC=-1360 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110100; // iC=-1548 
// vC = 14'b1111101011101110; // vC=-1298 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100000; // iC=-1504 
// vC = 14'b1111101101011100; // vC=-1188 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100100; // iC=-1564 
// vC = 14'b1111101001111111; // vC=-1409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110001; // iC=-1423 
// vC = 14'b1111101100111111; // vC=-1217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000110; // iC=-1402 
// vC = 14'b1111101010101100; // vC=-1364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010100; // iC=-1516 
// vC = 14'b1111101010101101; // vC=-1363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101000; // iC=-1496 
// vC = 14'b1111101011001111; // vC=-1329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100000; // iC=-1504 
// vC = 14'b1111101100000111; // vC=-1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110110; // iC=-1354 
// vC = 14'b1111101101000111; // vC=-1209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110101; // iC=-1611 
// vC = 14'b1111101001100010; // vC=-1438 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100100; // iC=-1628 
// vC = 14'b1111101001111000; // vC=-1416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000100; // iC=-1596 
// vC = 14'b1111101001101010; // vC=-1430 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011010; // iC=-1382 
// vC = 14'b1111101100000101; // vC=-1275 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010110; // iC=-1322 
// vC = 14'b1111101101000010; // vC=-1214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111100; // iC=-1348 
// vC = 14'b1111101101001011; // vC=-1205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000000; // iC=-1472 
// vC = 14'b1111101010011100; // vC=-1380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000001; // iC=-1599 
// vC = 14'b1111101011110011; // vC=-1293 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010110; // iC=-1450 
// vC = 14'b1111101010000110; // vC=-1402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111001; // iC=-1543 
// vC = 14'b1111101001101000; // vC=-1432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011011; // iC=-1573 
// vC = 14'b1111101100101010; // vC=-1238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110110; // iC=-1482 
// vC = 14'b1111101000011100; // vC=-1508 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110111; // iC=-1353 
// vC = 14'b1111101000100000; // vC=-1504 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101010; // iC=-1302 
// vC = 14'b1111100111111111; // vC=-1537 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000111; // iC=-1465 
// vC = 14'b1111101000111000; // vC=-1480 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110110; // iC=-1418 
// vC = 14'b1111101001110111; // vC=-1417 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100000; // iC=-1312 
// vC = 14'b1111101011000011; // vC=-1341 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001010; // iC=-1398 
// vC = 14'b1111101010101101; // vC=-1363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101000; // iC=-1304 
// vC = 14'b1111101010000111; // vC=-1401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110110; // iC=-1546 
// vC = 14'b1111101000010110; // vC=-1514 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101101; // iC=-1491 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001101; // iC=-1267 
// vC = 14'b1111101010111111; // vC=-1345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010100; // iC=-1516 
// vC = 14'b1111100111101100; // vC=-1556 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001011; // iC=-1269 
// vC = 14'b1111101000011100; // vC=-1508 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101100; // iC=-1492 
// vC = 14'b1111101010010101; // vC=-1387 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111101; // iC=-1411 
// vC = 14'b1111100110100110; // vC=-1626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100000; // iC=-1248 
// vC = 14'b1111101000000110; // vC=-1530 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000110; // iC=-1466 
// vC = 14'b1111101000111001; // vC=-1479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111010; // iC=-1350 
// vC = 14'b1111101000101100; // vC=-1492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010110; // iC=-1322 
// vC = 14'b1111100111011010; // vC=-1574 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000000; // iC=-1216 
// vC = 14'b1111100110100110; // vC=-1626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110111; // iC=-1417 
// vC = 14'b1111101001011011; // vC=-1445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101110; // iC=-1170 
// vC = 14'b1111101001001010; // vC=-1462 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000111; // iC=-1273 
// vC = 14'b1111101000000101; // vC=-1531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001010; // iC=-1334 
// vC = 14'b1111101001000111; // vC=-1465 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110101; // iC=-1355 
// vC = 14'b1111100111111100; // vC=-1540 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110011; // iC=-1229 
// vC = 14'b1111100111100111; // vC=-1561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110101; // iC=-1355 
// vC = 14'b1111101001110100; // vC=-1420 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000011; // iC=-1277 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000111; // iC=-1145 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101010; // iC=-1174 
// vC = 14'b1111100110100110; // vC=-1626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010100; // iC=-1196 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100011; // iC=-1181 
// vC = 14'b1111100111011100; // vC=-1572 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000111; // iC=-1209 
// vC = 14'b1111100101110111; // vC=-1673 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111101; // iC=-1347 
// vC = 14'b1111100101111100; // vC=-1668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000000; // iC=-1152 
// vC = 14'b1111100101111111; // vC=-1665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101000; // iC=-1176 
// vC = 14'b1111100101011010; // vC=-1702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111101; // iC=-1219 
// vC = 14'b1111100111000001; // vC=-1599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010101; // iC=-1259 
// vC = 14'b1111100110000001; // vC=-1663 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110001; // iC=-1103 
// vC = 14'b1111100111011000; // vC=-1576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001110; // iC=-1074 
// vC = 14'b1111100110001011; // vC=-1653 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010100; // iC=-1132 
// vC = 14'b1111100111001100; // vC=-1588 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000100; // iC=-1212 
// vC = 14'b1111101001001110; // vC=-1458 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100110; // iC=-1306 
// vC = 14'b1111100100000111; // vC=-1785 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001010; // iC=-1270 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000111; // iC=-1209 
// vC = 14'b1111101000111101; // vC=-1475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111010; // iC=-1030 
// vC = 14'b1111100101101011; // vC=-1685 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011010; // iC=-1126 
// vC = 14'b1111100111001011; // vC=-1589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111100; // iC=-1156 
// vC = 14'b1111100011111100; // vC=-1796 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010011; // iC=-1197 
// vC = 14'b1111100100001100; // vC=-1780 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001001; // iC=-1271 
// vC = 14'b1111100101101100; // vC=-1684 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110100; // iC=-1164 
// vC = 14'b1111100110011010; // vC=-1638 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111001; // iC=-1223 
// vC = 14'b1111100011101011; // vC=-1813 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000101; // iC=-1019 
// vC = 14'b1111100111001110; // vC=-1586 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111110; // iC=-1090 
// vC = 14'b1111100110010101; // vC=-1643 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b1111100110000110; // vC=-1658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101010; // iC=-1110 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000111; // iC=-1273 
// vC = 14'b1111100111100100; // vC=-1564 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010100; // iC=-1196 
// vC = 14'b1111100101111000; // vC=-1672 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110011; // iC=-1165 
// vC = 14'b1111100110000010; // vC=-1662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000001; // iC=-1087 
// vC = 14'b1111100111010111; // vC=-1577 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011100; // iC=-1188 
// vC = 14'b1111100101011101; // vC=-1699 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100111; // iC=-1177 
// vC = 14'b1111100011110101; // vC=-1803 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100110; // iC=-1050 
// vC = 14'b1111100101101111; // vC=-1681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101001; // iC= -919 
// vC = 14'b1111100011100111; // vC=-1817 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111010; // iC=-1158 
// vC = 14'b1111100101000001; // vC=-1727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010010; // iC=-1134 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101010; // iC=-1174 
// vC = 14'b1111100110001011; // vC=-1653 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000110; // iC= -890 
// vC = 14'b1111100100001010; // vC=-1782 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100111; // iC= -985 
// vC = 14'b1111100011100010; // vC=-1822 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110011; // iC= -909 
// vC = 14'b1111100010010000; // vC=-1904 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001101; // iC=-1011 
// vC = 14'b1111100110010110; // vC=-1642 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100000; // iC= -928 
// vC = 14'b1111100110011111; // vC=-1633 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100011; // iC= -861 
// vC = 14'b1111100110000100; // vC=-1660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011011; // iC=-1125 
// vC = 14'b1111100101010111; // vC=-1705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110000; // iC= -848 
// vC = 14'b1111100101111011; // vC=-1669 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000010; // iC=-1086 
// vC = 14'b1111100101011011; // vC=-1701 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001101; // iC= -883 
// vC = 14'b1111100010101111; // vC=-1873 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001001; // iC=-1015 
// vC = 14'b1111100010111100; // vC=-1860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010100; // iC=-1068 
// vC = 14'b1111100110011110; // vC=-1634 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111111; // iC= -833 
// vC = 14'b1111100101000101; // vC=-1723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010100; // iC=-1068 
// vC = 14'b1111100011100110; // vC=-1818 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100110; // iC=-1114 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110110; // iC=-1098 
// vC = 14'b1111100101000111; // vC=-1721 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001101; // iC= -883 
// vC = 14'b1111100101011100; // vC=-1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101001; // iC= -855 
// vC = 14'b1111100010110000; // vC=-1872 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011101; // iC= -803 
// vC = 14'b1111100011110101; // vC=-1803 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011100; // iC=-1060 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110101; // iC=-1035 
// vC = 14'b1111100010010100; // vC=-1900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001100; // iC= -820 
// vC = 14'b1111100010110001; // vC=-1871 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010000; // iC= -752 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101100; // iC= -852 
// vC = 14'b1111100010110011; // vC=-1869 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011011; // iC= -933 
// vC = 14'b1111100001101010; // vC=-1942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010010; // iC= -878 
// vC = 14'b1111100101010110; // vC=-1706 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101000; // iC= -984 
// vC = 14'b1111100011011110; // vC=-1826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010101; // iC= -747 
// vC = 14'b1111100001001001; // vC=-1975 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001111; // iC= -817 
// vC = 14'b1111100101100011; // vC=-1693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101010; // iC= -854 
// vC = 14'b1111100011010100; // vC=-1836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001110; // iC= -818 
// vC = 14'b1111100011111000; // vC=-1800 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011110; // iC= -802 
// vC = 14'b1111100010100011; // vC=-1885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101000; // iC= -984 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110011; // iC= -845 
// vC = 14'b1111100001110001; // vC=-1935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010011; // iC= -941 
// vC = 14'b1111100100101011; // vC=-1749 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011100; // iC= -932 
// vC = 14'b1111100011011010; // vC=-1830 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000111; // iC= -761 
// vC = 14'b1111100001110001; // vC=-1935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001010; // iC= -758 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100100; // iC= -924 
// vC = 14'b1111100010000010; // vC=-1918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100001; // iC= -735 
// vC = 14'b1111100001110101; // vC=-1931 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011001; // iC= -679 
// vC = 14'b1111100001011111; // vC=-1953 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000001; // iC= -767 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101110; // iC= -658 
// vC = 14'b1111100010011011; // vC=-1893 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000110; // iC= -890 
// vC = 14'b1111100000101111; // vC=-2001 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010010; // iC= -750 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001011; // iC= -693 
// vC = 14'b1111100000011010; // vC=-2022 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110011; // iC= -845 
// vC = 14'b1111100011101110; // vC=-1810 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111000; // iC= -904 
// vC = 14'b1111100011001111; // vC=-1841 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000111; // iC= -761 
// vC = 14'b1111100000111101; // vC=-1987 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101001; // iC= -663 
// vC = 14'b1111100001101111; // vC=-1937 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101111; // iC= -849 
// vC = 14'b1111100011101000; // vC=-1816 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000011; // iC= -573 
// vC = 14'b1111100001010101; // vC=-1963 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010000; // iC= -688 
// vC = 14'b1111100011000001; // vC=-1855 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111001; // iC= -839 
// vC = 14'b1111100000010001; // vC=-2031 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000111; // iC= -761 
// vC = 14'b1111100001100101; // vC=-1947 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011111; // iC= -865 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001010; // iC= -566 
// vC = 14'b1111100011011010; // vC=-1830 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111010; // iC= -774 
// vC = 14'b1111100000001011; // vC=-2037 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111100; // iC= -644 
// vC = 14'b1111011111010100; // vC=-2092 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111001; // iC= -775 
// vC = 14'b1111100001101000; // vC=-1944 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101000; // iC= -536 
// vC = 14'b1111100000010010; // vC=-2030 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000000; // iC= -640 
// vC = 14'b1111100001101011; // vC=-1941 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110101; // iC= -779 
// vC = 14'b1111011111001011; // vC=-2101 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001000; // iC= -632 
// vC = 14'b1111100011100111; // vC=-1817 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001010; // iC= -694 
// vC = 14'b1111100001001101; // vC=-1971 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011101; // iC= -611 
// vC = 14'b1111011111011001; // vC=-2087 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110101; // iC= -651 
// vC = 14'b1111100000111010; // vC=-1990 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111101; // iC= -579 
// vC = 14'b1111100011000001; // vC=-1855 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111110; // iC= -514 
// vC = 14'b1111100000000010; // vC=-2046 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101011; // iC= -405 
// vC = 14'b1111100010000101; // vC=-1915 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110111; // iC= -457 
// vC = 14'b1111100001010000; // vC=-1968 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001111; // iC= -369 
// vC = 14'b1111100000111000; // vC=-1992 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000010; // iC= -638 
// vC = 14'b1111100010111011; // vC=-1861 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100111; // iC= -537 
// vC = 14'b1111100000110111; // vC=-1993 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011110; // iC= -354 
// vC = 14'b1111011110111101; // vC=-2115 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110000; // iC= -592 
// vC = 14'b1111100000000111; // vC=-2041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100011; // iC= -477 
// vC = 14'b1111100000001110; // vC=-2034 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010101011; // iC= -341 
// vC = 14'b1111100010110111; // vC=-1865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010010; // iC= -494 
// vC = 14'b1111100010110001; // vC=-1871 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011111000; // iC= -264 
// vC = 14'b1111100010111000; // vC=-1864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111000; // iC= -392 
// vC = 14'b1111100000001101; // vC=-2035 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110001; // iC= -399 
// vC = 14'b1111011111010101; // vC=-2091 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100001; // iC= -415 
// vC = 14'b1111100011100001; // vC=-1823 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010110; // iC= -362 
// vC = 14'b1111011111101011; // vC=-2069 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001010; // iC= -246 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000011; // iC= -317 
// vC = 14'b1111011110101100; // vC=-2132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001010; // iC= -374 
// vC = 14'b1111100010000010; // vC=-1918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010101111; // iC= -337 
// vC = 14'b1111100010110001; // vC=-1871 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110010; // iC= -206 
// vC = 14'b1111100001100101; // vC=-1947 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011111; // iC= -289 
// vC = 14'b1111011111011111; // vC=-2081 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010001; // iC= -367 
// vC = 14'b1111100010010111; // vC=-1897 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000011; // iC= -125 
// vC = 14'b1111011110110010; // vC=-2126 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001000; // iC=  -56 
// vC = 14'b1111100010101001; // vC=-1879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011001; // iC= -295 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101110010; // iC= -142 
// vC = 14'b1111011110110011; // vC=-2125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110001; // iC= -207 
// vC = 14'b1111011111101110; // vC=-2066 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000001; // iC= -255 
// vC = 14'b1111100011000111; // vC=-1849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001001; // iC= -119 
// vC = 14'b1111100010111110; // vC=-1858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001011; // iC= -181 
// vC = 14'b1111011110111101; // vC=-2115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111011; // iC= -133 
// vC = 14'b1111100000001001; // vC=-2039 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111010; // iC=  122 
// vC = 14'b1111100010100010; // vC=-1886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010110; // iC= -106 
// vC = 14'b1111100000000111; // vC=-2041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110111; // iC=  119 
// vC = 14'b1111100001000101; // vC=-1979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101111; // iC=  175 
// vC = 14'b1111011111000110; // vC=-2106 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000111000; // iC=   56 
// vC = 14'b1111100010101000; // vC=-1880 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101110; // iC=  238 
// vC = 14'b1111100001100001; // vC=-1951 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000101; // iC=  197 
// vC = 14'b1111100000110010; // vC=-1998 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110100; // iC=  180 
// vC = 14'b1111100000000111; // vC=-2041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001000; // iC=   72 
// vC = 14'b1111100000101101; // vC=-2003 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111011; // iC=  187 
// vC = 14'b1111100011100010; // vC=-1822 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011110; // iC=  286 
// vC = 14'b1111100010011011; // vC=-1893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111010; // iC=  186 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100010; // iC=  354 
// vC = 14'b1111100000001111; // vC=-2033 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000010; // iC=  386 
// vC = 14'b1111100001110001; // vC=-1935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110111; // iC=  311 
// vC = 14'b1111011111101001; // vC=-2071 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000000; // iC=  320 
// vC = 14'b1111100010111011; // vC=-1861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101100; // iC=  236 
// vC = 14'b1111100001000001; // vC=-1983 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111100; // iC=  380 
// vC = 14'b1111100010100011; // vC=-1885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100000; // iC=  416 
// vC = 14'b1111100000110101; // vC=-1995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000101; // iC=  261 
// vC = 14'b1111100011000100; // vC=-1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111001; // iC=  441 
// vC = 14'b1111100000000001; // vC=-2047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100100; // iC=  612 
// vC = 14'b1111100010100011; // vC=-1885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010111; // iC=  407 
// vC = 14'b1111100001110011; // vC=-1933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011000; // iC=  408 
// vC = 14'b1111100001000011; // vC=-1981 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101010; // iC=  490 
// vC = 14'b1111100010101000; // vC=-1880 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010011; // iC=  467 
// vC = 14'b1111100011001110; // vC=-1842 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110111; // iC=  695 
// vC = 14'b1111100000111011; // vC=-1989 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110111; // iC=  759 
// vC = 14'b1111100001000111; // vC=-1977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001100; // iC=  652 
// vC = 14'b1111011111010111; // vC=-2089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100001; // iC=  609 
// vC = 14'b1111100000011111; // vC=-2017 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011111; // iC=  799 
// vC = 14'b1111100001001011; // vC=-1973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100000; // iC=  608 
// vC = 14'b1111011111110000; // vC=-2064 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010011; // iC=  851 
// vC = 14'b1111100001010011; // vC=-1965 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111100; // iC=  764 
// vC = 14'b1111100010110100; // vC=-1868 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110101; // iC=  821 
// vC = 14'b1111100001010111; // vC=-1961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000100; // iC=  836 
// vC = 14'b1111100000111100; // vC=-1988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101000; // iC=  744 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000010; // iC=  962 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001101; // iC=  973 
// vC = 14'b1111100100010111; // vC=-1769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110111; // iC=  951 
// vC = 14'b1111100010010010; // vC=-1902 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101101; // iC= 1005 
// vC = 14'b1111100001101111; // vC=-1937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111010; // iC=  762 
// vC = 14'b1111100010000011; // vC=-1917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101110; // iC= 1006 
// vC = 14'b1111100100011111; // vC=-1761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011101; // iC= 1117 
// vC = 14'b1111100010010000; // vC=-1904 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100100; // iC=  868 
// vC = 14'b1111100001001110; // vC=-1970 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011110; // iC=  990 
// vC = 14'b1111100001110010; // vC=-1934 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011100; // iC= 1052 
// vC = 14'b1111100100010011; // vC=-1773 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010100; // iC=  916 
// vC = 14'b1111100011111010; // vC=-1798 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010011; // iC=  915 
// vC = 14'b1111100010010001; // vC=-1903 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101000; // iC= 1192 
// vC = 14'b1111100000011100; // vC=-2020 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011000; // iC= 1112 
// vC = 14'b1111100001010110; // vC=-1962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110100; // iC= 1012 
// vC = 14'b1111100100000101; // vC=-1787 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001010; // iC= 1162 
// vC = 14'b1111100010000000; // vC=-1920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010011; // iC= 1299 
// vC = 14'b1111100011101011; // vC=-1813 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000010; // iC= 1218 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000111; // iC= 1223 
// vC = 14'b1111100010110101; // vC=-1867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110111; // iC= 1335 
// vC = 14'b1111100011101010; // vC=-1814 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111101; // iC= 1341 
// vC = 14'b1111100100010111; // vC=-1769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110000; // iC= 1328 
// vC = 14'b1111100010111101; // vC=-1859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000111; // iC= 1287 
// vC = 14'b1111100011001011; // vC=-1845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101111; // iC= 1263 
// vC = 14'b1111100010010010; // vC=-1902 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000110; // iC= 1286 
// vC = 14'b1111100011100000; // vC=-1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101101; // iC= 1197 
// vC = 14'b1111100011100100; // vC=-1820 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100110; // iC= 1446 
// vC = 14'b1111100010111011; // vC=-1861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110010; // iC= 1394 
// vC = 14'b1111100100110110; // vC=-1738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001011; // iC= 1547 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110111; // iC= 1399 
// vC = 14'b1111100110001010; // vC=-1654 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010111; // iC= 1303 
// vC = 14'b1111100011010001; // vC=-1839 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101101; // iC= 1389 
// vC = 14'b1111100011001000; // vC=-1848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111110; // iC= 1598 
// vC = 14'b1111100010001100; // vC=-1908 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100101; // iC= 1317 
// vC = 14'b1111100110000100; // vC=-1660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101111; // iC= 1455 
// vC = 14'b1111100101100110; // vC=-1690 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111001; // iC= 1401 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001011; // iC= 1675 
// vC = 14'b1111100100100110; // vC=-1754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001111; // iC= 1615 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100111; // iC= 1511 
// vC = 14'b1111100010111001; // vC=-1863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000111; // iC= 1415 
// vC = 14'b1111100100101011; // vC=-1749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110010; // iC= 1586 
// vC = 14'b1111100111101110; // vC=-1554 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010110; // iC= 1686 
// vC = 14'b1111100011111010; // vC=-1798 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100110; // iC= 1702 
// vC = 14'b1111100101111100; // vC=-1668 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000000; // iC= 1664 
// vC = 14'b1111101000001001; // vC=-1527 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000100; // iC= 1796 
// vC = 14'b1111100110011011; // vC=-1637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100000; // iC= 1632 
// vC = 14'b1111100100011010; // vC=-1766 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110011; // iC= 1523 
// vC = 14'b1111100101110000; // vC=-1680 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111111; // iC= 1791 
// vC = 14'b1111100101100000; // vC=-1696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100010; // iC= 1762 
// vC = 14'b1111100110011100; // vC=-1636 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100000; // iC= 1760 
// vC = 14'b1111100111110101; // vC=-1547 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111000; // iC= 1592 
// vC = 14'b1111100101000101; // vC=-1723 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011100; // iC= 1820 
// vC = 14'b1111101001010001; // vC=-1455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100010; // iC= 1890 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111111; // iC= 1855 
// vC = 14'b1111100111110011; // vC=-1549 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111011; // iC= 1851 
// vC = 14'b1111101001000001; // vC=-1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000100; // iC= 1860 
// vC = 14'b1111101001010101; // vC=-1451 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110010; // iC= 1650 
// vC = 14'b1111100110011001; // vC=-1639 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000111; // iC= 1671 
// vC = 14'b1111100111011011; // vC=-1573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000001; // iC= 1793 
// vC = 14'b1111101001011001; // vC=-1447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010001; // iC= 1681 
// vC = 14'b1111101001110000; // vC=-1424 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001110; // iC= 1678 
// vC = 14'b1111100110110110; // vC=-1610 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011010; // iC= 1818 
// vC = 14'b1111101001100111; // vC=-1433 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b1111100110101010; // vC=-1622 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b1111101001000110; // vC=-1466 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111011; // iC= 1723 
// vC = 14'b1111101010011111; // vC=-1377 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010011; // iC= 1747 
// vC = 14'b1111101010101001; // vC=-1367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001000; // iC= 1736 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001000; // iC= 1864 
// vC = 14'b1111101011000101; // vC=-1339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b1111101011011111; // vC=-1313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111100; // iC= 1788 
// vC = 14'b1111101010000101; // vC=-1403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001001; // iC= 2057 
// vC = 14'b1111101000101001; // vC=-1495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100101; // iC= 1829 
// vC = 14'b1111100111011111; // vC=-1569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001001; // iC= 1801 
// vC = 14'b1111101011000010; // vC=-1342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011111; // iC= 1823 
// vC = 14'b1111100111010010; // vC=-1582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b1111100111111001; // vC=-1543 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b1111101000001110; // vC=-1522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b1111101100100011; // vC=-1245 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001111; // iC= 1807 
// vC = 14'b1111101010000111; // vC=-1401 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000111; // iC= 2055 
// vC = 14'b1111101010001101; // vC=-1395 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001101; // iC= 1805 
// vC = 14'b1111101001011110; // vC=-1442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001000; // iC= 1864 
// vC = 14'b1111101001101110; // vC=-1426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010011; // iC= 2067 
// vC = 14'b1111101001100111; // vC=-1433 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b1111101101100000; // vC=-1184 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b1111101101101000; // vC=-1176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000000; // iC= 2048 
// vC = 14'b1111101001011111; // vC=-1441 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111101010110100; // vC=-1356 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b1111101001100001; // vC=-1439 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101111; // iC= 1903 
// vC = 14'b1111101001100010; // vC=-1438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101010; // iC= 2090 
// vC = 14'b1111101110000011; // vC=-1149 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001110; // iC= 1934 
// vC = 14'b1111101100011100; // vC=-1252 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b1111101010001011; // vC=-1397 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b1111101011001010; // vC=-1334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101110; // iC= 2158 
// vC = 14'b1111101101001100; // vC=-1204 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111101111000011; // vC=-1085 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001010; // iC= 1994 
// vC = 14'b1111101101111011; // vC=-1157 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111101; // iC= 2109 
// vC = 14'b1111101101111001; // vC=-1159 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001111; // iC= 2127 
// vC = 14'b1111101101011110; // vC=-1186 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110001; // iC= 1905 
// vC = 14'b1111101100000000; // vC=-1280 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000111; // iC= 2183 
// vC = 14'b1111101101101101; // vC=-1171 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b1111101111110000; // vC=-1040 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001101; // iC= 2189 
// vC = 14'b1111101100001011; // vC=-1269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b1111101011111000; // vC=-1288 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101101; // iC= 2157 
// vC = 14'b1111101110001111; // vC=-1137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b1111101110001000; // vC=-1144 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111101; // iC= 2109 
// vC = 14'b1111101111101100; // vC=-1044 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010110; // iC= 2134 
// vC = 14'b1111101100000010; // vC=-1278 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b1111101011111010; // vC=-1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b1111101101001110; // vC=-1202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000001; // iC= 2049 
// vC = 14'b1111110001001100; // vC= -948 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101011; // iC= 1963 
// vC = 14'b1111101111100111; // vC=-1049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111101100101000; // vC=-1240 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b1111110000000011; // vC=-1021 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b1111110000011010; // vC= -998 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b1111110000110000; // vC= -976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111101; // iC= 2173 
// vC = 14'b1111101101111001; // vC=-1159 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111110001110101; // vC= -907 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000001; // iC= 1921 
// vC = 14'b1111101111001111; // vC=-1073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101100; // iC= 2156 
// vC = 14'b1111101111000111; // vC=-1081 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110100; // iC= 2036 
// vC = 14'b1111101110111011; // vC=-1093 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000101; // iC= 2181 
// vC = 14'b1111101111011110; // vC=-1058 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101100; // iC= 2156 
// vC = 14'b1111110001100101; // vC= -923 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111110010000000; // vC= -896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110101; // iC= 2101 
// vC = 14'b1111101110110001; // vC=-1103 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000101; // iC= 2117 
// vC = 14'b1111101111110000; // vC=-1040 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111101; // iC= 2173 
// vC = 14'b1111110000100010; // vC= -990 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100110; // iC= 2214 
// vC = 14'b1111110001111100; // vC= -900 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110001; // iC= 2161 
// vC = 14'b1111110010100100; // vC= -860 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111110011011011; // vC= -805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111111; // iC= 2111 
// vC = 14'b1111110000110111; // vC= -969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100111; // iC= 2151 
// vC = 14'b1111110000100010; // vC= -990 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000011; // iC= 2051 
// vC = 14'b1111110000001101; // vC=-1011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011010; // iC= 2202 
// vC = 14'b1111110011110010; // vC= -782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111010; // iC= 2106 
// vC = 14'b1111110001001110; // vC= -946 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110011; // iC= 2163 
// vC = 14'b1111101111111011; // vC=-1029 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b1111110100110011; // vC= -717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000100; // iC= 1924 
// vC = 14'b1111110011100101; // vC= -795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b1111110100010010; // vC= -750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001101; // iC= 2189 
// vC = 14'b1111110100001011; // vC= -757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100011; // iC= 1955 
// vC = 14'b1111110011110100; // vC= -780 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001000; // iC= 2184 
// vC = 14'b1111110000110101; // vC= -971 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011011; // iC= 2075 
// vC = 14'b1111110011111001; // vC= -775 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111110100100101; // vC= -731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b1111110101101100; // vC= -660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b1111110010101111; // vC= -849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b1111110010110011; // vC= -845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000111; // iC= 2247 
// vC = 14'b1111110010000000; // vC= -896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b1111110011011010; // vC= -806 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001001; // iC= 2185 
// vC = 14'b1111110011000110; // vC= -826 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111100; // iC= 2108 
// vC = 14'b1111110011001011; // vC= -821 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111110011100100; // vC= -796 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000111; // iC= 2055 
// vC = 14'b1111110111000001; // vC= -575 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101111; // iC= 2095 
// vC = 14'b1111110011000001; // vC= -831 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b1111110100100011; // vC= -733 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100010; // iC= 1954 
// vC = 14'b1111110110011111; // vC= -609 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101010; // iC= 2090 
// vC = 14'b1111110011111101; // vC= -771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000100; // iC= 2244 
// vC = 14'b1111110010110111; // vC= -841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b1111110100101101; // vC= -723 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b1111111000000000; // vC= -512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111110100011001; // vC= -743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010011; // iC= 2131 
// vC = 14'b1111110111010001; // vC= -559 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011101; // iC= 2205 
// vC = 14'b1111110011101000; // vC= -792 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000101; // iC= 1989 
// vC = 14'b1111110100110010; // vC= -718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101100; // iC= 2092 
// vC = 14'b1111110100110011; // vC= -717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110011; // iC= 2227 
// vC = 14'b1111111000001011; // vC= -501 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110000; // iC= 2032 
// vC = 14'b1111110111011111; // vC= -545 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011001; // iC= 2137 
// vC = 14'b1111110110001000; // vC= -632 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110111; // iC= 2039 
// vC = 14'b1111110111100011; // vC= -541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001111; // iC= 2127 
// vC = 14'b1111110111001100; // vC= -564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b1111111001100001; // vC= -415 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010111; // iC= 2199 
// vC = 14'b1111110111010010; // vC= -558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100010; // iC= 1954 
// vC = 14'b1111111000010111; // vC= -489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b1111111000100001; // vC= -479 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011010; // iC= 2202 
// vC = 14'b1111110101100110; // vC= -666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101111; // iC= 2159 
// vC = 14'b1111110111111000; // vC= -520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011010; // iC= 2074 
// vC = 14'b1111111001010100; // vC= -428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101011; // iC= 1963 
// vC = 14'b1111110111101001; // vC= -535 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001110; // iC= 2126 
// vC = 14'b1111110110000001; // vC= -639 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b1111110111100011; // vC= -541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100001; // iC= 2209 
// vC = 14'b1111110111010100; // vC= -556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000111; // iC= 2055 
// vC = 14'b1111110111010100; // vC= -556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110000; // iC= 2224 
// vC = 14'b1111111001001001; // vC= -439 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111010; // iC= 1978 
// vC = 14'b1111110111100101; // vC= -539 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b1111110111101110; // vC= -530 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110001; // iC= 2161 
// vC = 14'b1111111001111000; // vC= -392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001011; // iC= 2251 
// vC = 14'b1111111011100001; // vC= -287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100001; // iC= 2017 
// vC = 14'b1111111011011000; // vC= -296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b1111111000001110; // vC= -498 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b1111111011101010; // vC= -278 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000100; // iC= 2116 
// vC = 14'b1111111010110101; // vC= -331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b1111111100110010; // vC= -206 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111110; // iC= 2238 
// vC = 14'b1111111011011010; // vC= -294 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001001; // iC= 2249 
// vC = 14'b1111111001001010; // vC= -438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110000; // iC= 2224 
// vC = 14'b1111111010111001; // vC= -327 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001001; // iC= 2121 
// vC = 14'b1111111001101011; // vC= -405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110110; // iC= 1974 
// vC = 14'b1111111001101000; // vC= -408 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011000; // iC= 2136 
// vC = 14'b1111111001100011; // vC= -413 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101111; // iC= 2095 
// vC = 14'b1111111101101110; // vC= -146 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110110; // iC= 2102 
// vC = 14'b1111111100011100; // vC= -228 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111111; // iC= 2239 
// vC = 14'b1111111010001111; // vC= -369 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010010; // iC= 2066 
// vC = 14'b1111111100111110; // vC= -194 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110001; // iC= 1969 
// vC = 14'b1111111010101101; // vC= -339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011111; // iC= 2207 
// vC = 14'b1111111101010111; // vC= -169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b1111111010110011; // vC= -333 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001001; // iC= 2249 
// vC = 14'b1111111010011010; // vC= -358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110010; // iC= 2034 
// vC = 14'b1111111101001011; // vC= -181 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b1111111010010110; // vC= -362 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110101; // iC= 2229 
// vC = 14'b1111111011011011; // vC= -293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b1111111101010000; // vC= -176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100000; // iC= 2208 
// vC = 14'b1111111110001010; // vC= -118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111111101111010; // vC= -134 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110101; // iC= 2165 
// vC = 14'b1111111011111000; // vC= -264 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100001; // iC= 2017 
// vC = 14'b1111111111011011; // vC=  -37 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000011; // iC= 1923 
// vC = 14'b1111111011010111; // vC= -297 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b1111111101000011; // vC= -189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b1111111110111100; // vC=  -68 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b1111111110111001; // vC=  -71 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111111110011000; // vC= -104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110101; // iC= 2165 
// vC = 14'b1111111100110101; // vC= -203 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b0000000000010111; // vC=   23 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110111; // iC= 2231 
// vC = 14'b1111111100010101; // vC= -235 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100010; // iC= 2082 
// vC = 14'b1111111100010011; // vC= -237 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001110; // iC= 2126 
// vC = 14'b1111111100010010; // vC= -238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101010; // iC= 2218 
// vC = 14'b1111111101100001; // vC= -159 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110110; // iC= 1974 
// vC = 14'b1111111100100110; // vC= -218 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b1111111101110111; // vC= -137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101101; // iC= 2157 
// vC = 14'b0000000001111000; // vC=  120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010001; // iC= 2129 
// vC = 14'b0000000010001001; // vC=  137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001011; // iC= 2187 
// vC = 14'b1111111110110100; // vC=  -76 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111010; // iC= 1914 
// vC = 14'b1111111110101111; // vC=  -81 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b0000000010010110; // vC=  150 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111111111010111; // vC=  -41 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b0000000000010001; // vC=   17 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101011; // iC= 1899 
// vC = 14'b1111111111100000; // vC=  -32 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001000; // iC= 1928 
// vC = 14'b1111111111100001; // vC=  -31 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b0000000011010101; // vC=  213 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b0000000011010111; // vC=  215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111010; // iC= 2170 
// vC = 14'b0000000011100011; // vC=  227 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b1111111111000111; // vC=  -57 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001010; // iC= 2186 
// vC = 14'b0000000000101010; // vC=   42 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b0000000001110110; // vC=  118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110000; // iC= 1904 
// vC = 14'b0000000000011100; // vC=   28 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110011; // iC= 1907 
// vC = 14'b0000000010110001; // vC=  177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001001; // iC= 1993 
// vC = 14'b0000000010010111; // vC=  151 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110011; // iC= 2099 
// vC = 14'b0000000010001111; // vC=  143 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b0000000011010010; // vC=  210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001001; // iC= 2121 
// vC = 14'b0000000010000010; // vC=  130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b0000000010100100; // vC=  164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b0000000000101011; // vC=   43 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000000; // iC= 2112 
// vC = 14'b0000000100001010; // vC=  266 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101111; // iC= 1967 
// vC = 14'b0000000000110111; // vC=   55 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b0000000000100010; // vC=   34 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111100; // iC= 1916 
// vC = 14'b0000000101010111; // vC=  343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100111; // iC= 2023 
// vC = 14'b0000000010100101; // vC=  165 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010010; // iC= 2130 
// vC = 14'b0000000101111000; // vC=  376 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b0000000100000010; // vC=  258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b0000000100111100; // vC=  316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b0000000101010110; // vC=  342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010100; // iC= 2132 
// vC = 14'b0000000100100101; // vC=  293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110101; // iC= 2101 
// vC = 14'b0000000011001010; // vC=  202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b0000000001101100; // vC=  108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100110; // iC= 2022 
// vC = 14'b0000000011001011; // vC=  203 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b0000000010101010; // vC=  170 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b0000000011011000; // vC=  216 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b0000000011000101; // vC=  197 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110011; // iC= 1907 
// vC = 14'b0000000010100110; // vC=  166 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111110; // iC= 1854 
// vC = 14'b0000000110010000; // vC=  400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011000; // iC= 2136 
// vC = 14'b0000000010101110; // vC=  174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b0000000111110010; // vC=  498 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b0000000111001101; // vC=  461 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b0000000011010100; // vC=  212 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110001; // iC= 1969 
// vC = 14'b0000000111011000; // vC=  472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001111; // iC= 2063 
// vC = 14'b0000000101101111; // vC=  367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001001; // iC= 2121 
// vC = 14'b0000001000010110; // vC=  534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b0000000110111110; // vC=  446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b0000000101011001; // vC=  345 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111011; // iC= 1915 
// vC = 14'b0000000111010011; // vC=  467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b0000001000010010; // vC=  530 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100010; // iC= 2018 
// vC = 14'b0000000101001101; // vC=  333 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b0000000111011010; // vC=  474 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b0000000110000010; // vC=  386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010111; // iC= 1815 
// vC = 14'b0000001001001100; // vC=  588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101111; // iC= 1839 
// vC = 14'b0000001000011100; // vC=  540 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101000; // iC= 1832 
// vC = 14'b0000000101100000; // vC=  352 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b0000001000100010; // vC=  546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b0000000101010100; // vC=  340 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100101; // iC= 1829 
// vC = 14'b0000000111111011; // vC=  507 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111110; // iC= 1982 
// vC = 14'b0000000110101100; // vC=  428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b0000000111100101; // vC=  485 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b0000000111101101; // vC=  493 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011101; // iC= 1885 
// vC = 14'b0000001001000111; // vC=  583 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101101; // iC= 2093 
// vC = 14'b0000000111010011; // vC=  467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111101; // iC= 1789 
// vC = 14'b0000001001110111; // vC=  631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b0000000110001101; // vC=  397 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100110; // iC= 1766 
// vC = 14'b0000000111011111; // vC=  479 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b0000001001110000; // vC=  624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b0000000111101110; // vC=  494 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001111; // iC= 1999 
// vC = 14'b0000001001101010; // vC=  618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101000; // iC= 2024 
// vC = 14'b0000000111100001; // vC=  481 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b0000001011010011; // vC=  723 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000000; // iC= 1792 
// vC = 14'b0000001010100011; // vC=  675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b0000001000100110; // vC=  550 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000000; // iC= 1792 
// vC = 14'b0000001010001100; // vC=  652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001000; // iC= 1864 
// vC = 14'b0000001010101111; // vC=  687 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011000; // iC= 1816 
// vC = 14'b0000001000100101; // vC=  549 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111101; // iC= 1789 
// vC = 14'b0000001000100100; // vC=  548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001101; // iC= 1869 
// vC = 14'b0000001011101100; // vC=  748 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110110; // iC= 1974 
// vC = 14'b0000001011001011; // vC=  715 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110111; // iC= 1911 
// vC = 14'b0000001000110001; // vC=  561 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111000; // iC= 1976 
// vC = 14'b0000001100001110; // vC=  782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101001; // iC= 1769 
// vC = 14'b0000001001111101; // vC=  637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b0000001011001010; // vC=  714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111110; // iC= 1918 
// vC = 14'b0000001000100100; // vC=  548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011111; // iC= 1759 
// vC = 14'b0000001001100110; // vC=  614 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b0000001011011100; // vC=  732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010001; // iC= 1809 
// vC = 14'b0000001010110110; // vC=  694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b0000001100011001; // vC=  793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b0000001100101100; // vC=  812 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111101; // iC= 1725 
// vC = 14'b0000001001100101; // vC=  613 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101001; // iC= 1833 
// vC = 14'b0000001010101010; // vC=  682 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111001; // iC= 1785 
// vC = 14'b0000001110010000; // vC=  912 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000100; // iC= 1860 
// vC = 14'b0000001010100111; // vC=  679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001110; // iC= 1678 
// vC = 14'b0000001110100011; // vC=  931 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b0000001101000111; // vC=  839 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100010; // iC= 1954 
// vC = 14'b0000001100010110; // vC=  790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100011; // iC= 1699 
// vC = 14'b0000001011011011; // vC=  731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b0000001011011101; // vC=  733 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101110; // iC= 1838 
// vC = 14'b0000001010111100; // vC=  700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b0000001110000100; // vC=  900 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000001; // iC= 1665 
// vC = 14'b0000001110010000; // vC=  912 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010100; // iC= 1876 
// vC = 14'b0000001011111011; // vC=  763 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011000; // iC= 1752 
// vC = 14'b0000001110010010; // vC=  914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001001; // iC= 1801 
// vC = 14'b0000001111010011; // vC=  979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b0000001100111110; // vC=  830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b0000001011010110; // vC=  726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011101; // iC= 1693 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111011; // iC= 1659 
// vC = 14'b0000001110101011; // vC=  939 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011000; // iC= 1688 
// vC = 14'b0000001100111010; // vC=  826 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011100; // iC= 1884 
// vC = 14'b0000001101000110; // vC=  838 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110011; // iC= 1907 
// vC = 14'b0000001011101101; // vC=  749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010011; // iC= 1747 
// vC = 14'b0000001011111101; // vC=  765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010001; // iC= 1617 
// vC = 14'b0000001101000000; // vC=  832 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110101; // iC= 1653 
// vC = 14'b0000001110101010; // vC=  938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011000; // iC= 1880 
// vC = 14'b0000001100011011; // vC=  795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111010; // iC= 1594 
// vC = 14'b0000001110010000; // vC=  912 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100001; // iC= 1825 
// vC = 14'b0000001111010010; // vC=  978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011100; // iC= 1756 
// vC = 14'b0000010000110000; // vC= 1072 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100000; // iC= 1824 
// vC = 14'b0000001100100110; // vC=  806 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101110; // iC= 1838 
// vC = 14'b0000001110111010; // vC=  954 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101001; // iC= 1833 
// vC = 14'b0000001111100101; // vC=  997 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101001; // iC= 1577 
// vC = 14'b0000001111111111; // vC= 1023 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101001; // iC= 1641 
// vC = 14'b0000010000001110; // vC= 1038 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001011; // iC= 1867 
// vC = 14'b0000010001100101; // vC= 1125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011101; // iC= 1565 
// vC = 14'b0000001111011001; // vC=  985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100110; // iC= 1574 
// vC = 14'b0000001111101010; // vC= 1002 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001010; // iC= 1866 
// vC = 14'b0000001110110000; // vC=  944 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100000; // iC= 1824 
// vC = 14'b0000001111011010; // vC=  986 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011100; // iC= 1756 
// vC = 14'b0000001111010001; // vC=  977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111011; // iC= 1723 
// vC = 14'b0000010001110110; // vC= 1142 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110011; // iC= 1587 
// vC = 14'b0000001101111110; // vC=  894 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110010; // iC= 1522 
// vC = 14'b0000010010000000; // vC= 1152 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000011; // iC= 1731 
// vC = 14'b0000001110010010; // vC=  914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101001; // iC= 1705 
// vC = 14'b0000010001000111; // vC= 1095 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100100; // iC= 1764 
// vC = 14'b0000001111000000; // vC=  960 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101000; // iC= 1576 
// vC = 14'b0000001110101001; // vC=  937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101010; // iC= 1642 
// vC = 14'b0000010001010010; // vC= 1106 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111011; // iC= 1787 
// vC = 14'b0000010000110101; // vC= 1077 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010110; // iC= 1558 
// vC = 14'b0000010010100100; // vC= 1188 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001101; // iC= 1677 
// vC = 14'b0000010001101001; // vC= 1129 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000101; // iC= 1669 
// vC = 14'b0000010001011001; // vC= 1113 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110100; // iC= 1524 
// vC = 14'b0000010010010100; // vC= 1172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011110; // iC= 1630 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110010; // iC= 1714 
// vC = 14'b0000010100001110; // vC= 1294 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100001; // iC= 1697 
// vC = 14'b0000001111111010; // vC= 1018 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111100; // iC= 1596 
// vC = 14'b0000010011100111; // vC= 1255 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010000; // iC= 1616 
// vC = 14'b0000010010000000; // vC= 1152 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100001; // iC= 1697 
// vC = 14'b0000010000000010; // vC= 1026 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000101; // iC= 1669 
// vC = 14'b0000010100000011; // vC= 1283 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110000; // iC= 1584 
// vC = 14'b0000010011000011; // vC= 1219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001000; // iC= 1480 
// vC = 14'b0000010000101010; // vC= 1066 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011111; // iC= 1503 
// vC = 14'b0000010010101101; // vC= 1197 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100101; // iC= 1701 
// vC = 14'b0000010010001101; // vC= 1165 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111011; // iC= 1467 
// vC = 14'b0000010001101111; // vC= 1135 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100000; // iC= 1568 
// vC = 14'b0000010000100001; // vC= 1057 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010110; // iC= 1622 
// vC = 14'b0000010011101101; // vC= 1261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000010; // iC= 1538 
// vC = 14'b0000010100010001; // vC= 1297 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010111; // iC= 1431 
// vC = 14'b0000010011000001; // vC= 1217 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110111; // iC= 1527 
// vC = 14'b0000010100111111; // vC= 1343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101001; // iC= 1577 
// vC = 14'b0000010010010011; // vC= 1171 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010100; // iC= 1620 
// vC = 14'b0000010001011001; // vC= 1113 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010101; // iC= 1685 
// vC = 14'b0000010001101101; // vC= 1133 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110000; // iC= 1456 
// vC = 14'b0000010011001100; // vC= 1228 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010001; // iC= 1617 
// vC = 14'b0000010011011011; // vC= 1243 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011001; // iC= 1689 
// vC = 14'b0000010001100000; // vC= 1120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000100; // iC= 1604 
// vC = 14'b0000010010101110; // vC= 1198 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011011; // iC= 1371 
// vC = 14'b0000010011001011; // vC= 1227 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111000; // iC= 1528 
// vC = 14'b0000010010100100; // vC= 1188 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001111; // iC= 1615 
// vC = 14'b0000010101101010; // vC= 1386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001100; // iC= 1676 
// vC = 14'b0000010011011001; // vC= 1241 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110001; // iC= 1457 
// vC = 14'b0000010010011001; // vC= 1177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101010; // iC= 1578 
// vC = 14'b0000010100101000; // vC= 1320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001011; // iC= 1355 
// vC = 14'b0000010110011000; // vC= 1432 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110001; // iC= 1521 
// vC = 14'b0000010110010110; // vC= 1430 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100111; // iC= 1447 
// vC = 14'b0000010011111000; // vC= 1272 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000001; // iC= 1473 
// vC = 14'b0000010011100111; // vC= 1255 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101010; // iC= 1514 
// vC = 14'b0000010110110001; // vC= 1457 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011101; // iC= 1373 
// vC = 14'b0000010111001100; // vC= 1484 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010101; // iC= 1365 
// vC = 14'b0000010110100011; // vC= 1443 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101001; // iC= 1513 
// vC = 14'b0000010011111010; // vC= 1274 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011011; // iC= 1499 
// vC = 14'b0000010100110011; // vC= 1331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010010; // iC= 1426 
// vC = 14'b0000010101101010; // vC= 1386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010111; // iC= 1495 
// vC = 14'b0000011000001111; // vC= 1551 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111110; // iC= 1534 
// vC = 14'b0000010100100101; // vC= 1317 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101110; // iC= 1582 
// vC = 14'b0000010101101100; // vC= 1388 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101101; // iC= 1581 
// vC = 14'b0000010111111011; // vC= 1531 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010010; // iC= 1426 
// vC = 14'b0000010011101001; // vC= 1257 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000011; // iC= 1475 
// vC = 14'b0000011000101110; // vC= 1582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100011; // iC= 1315 
// vC = 14'b0000010101011011; // vC= 1371 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111001; // iC= 1465 
// vC = 14'b0000010100100101; // vC= 1317 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001010; // iC= 1546 
// vC = 14'b0000011000110101; // vC= 1589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b0000010110001100; // vC= 1420 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010001; // iC= 1233 
// vC = 14'b0000011000100000; // vC= 1568 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111111; // iC= 1279 
// vC = 14'b0000010101110110; // vC= 1398 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010110; // iC= 1238 
// vC = 14'b0000010100101001; // vC= 1321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110001; // iC= 1265 
// vC = 14'b0000010101101110; // vC= 1390 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011010; // iC= 1306 
// vC = 14'b0000010101110100; // vC= 1396 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111110; // iC= 1214 
// vC = 14'b0000010110010000; // vC= 1424 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010000; // iC= 1424 
// vC = 14'b0000011001000010; // vC= 1602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101001; // iC= 1385 
// vC = 14'b0000011000110010; // vC= 1586 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011110; // iC= 1438 
// vC = 14'b0000010101111000; // vC= 1400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000110; // iC= 1286 
// vC = 14'b0000011001001011; // vC= 1611 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001000; // iC= 1416 
// vC = 14'b0000010111101110; // vC= 1518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001111; // iC= 1295 
// vC = 14'b0000011001111101; // vC= 1661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100100; // iC= 1252 
// vC = 14'b0000011001000101; // vC= 1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101000; // iC= 1192 
// vC = 14'b0000010111010001; // vC= 1489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101100; // iC= 1388 
// vC = 14'b0000011010001000; // vC= 1672 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010110; // iC= 1238 
// vC = 14'b0000010110100001; // vC= 1441 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101101; // iC= 1325 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100100; // iC= 1316 
// vC = 14'b0000010101110100; // vC= 1396 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000111; // iC= 1159 
// vC = 14'b0000011010100110; // vC= 1702 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111001; // iC= 1209 
// vC = 14'b0000011001001000; // vC= 1608 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001000; // iC= 1224 
// vC = 14'b0000010111001000; // vC= 1480 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100000; // iC= 1312 
// vC = 14'b0000011000010111; // vC= 1559 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010010; // iC= 1298 
// vC = 14'b0000011001110111; // vC= 1655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110100; // iC= 1396 
// vC = 14'b0000011000011000; // vC= 1560 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101110; // iC= 1134 
// vC = 14'b0000010110110100; // vC= 1460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101010; // iC= 1322 
// vC = 14'b0000011010010100; // vC= 1684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010111; // iC= 1303 
// vC = 14'b0000010111111010; // vC= 1530 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100001; // iC= 1249 
// vC = 14'b0000011000100010; // vC= 1570 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001000; // iC= 1288 
// vC = 14'b0000011011010111; // vC= 1751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101101; // iC= 1133 
// vC = 14'b0000010111011000; // vC= 1496 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001110; // iC= 1358 
// vC = 14'b0000011001111111; // vC= 1663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101101; // iC= 1261 
// vC = 14'b0000010111100101; // vC= 1509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110110; // iC= 1142 
// vC = 14'b0000011000110100; // vC= 1588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001000; // iC= 1224 
// vC = 14'b0000011010011100; // vC= 1692 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011010; // iC= 1178 
// vC = 14'b0000011011101110; // vC= 1774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001110; // iC= 1102 
// vC = 14'b0000011010010110; // vC= 1686 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101101; // iC= 1133 
// vC = 14'b0000011011000110; // vC= 1734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000111; // iC= 1031 
// vC = 14'b0000011000100100; // vC= 1572 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111111; // iC= 1343 
// vC = 14'b0000011001010010; // vC= 1618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001111; // iC= 1231 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001011; // iC= 1163 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001111; // iC= 1167 
// vC = 14'b0000011000100100; // vC= 1572 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011111; // iC= 1183 
// vC = 14'b0000011010010011; // vC= 1683 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110110; // iC= 1270 
// vC = 14'b0000011000001001; // vC= 1545 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111100; // iC= 1084 
// vC = 14'b0000011011000110; // vC= 1734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111001; // iC= 1017 
// vC = 14'b0000011011100010; // vC= 1762 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000010; // iC= 1026 
// vC = 14'b0000010111111111; // vC= 1535 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100101; // iC=  997 
// vC = 14'b0000011000000011; // vC= 1539 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001000; // iC= 1160 
// vC = 14'b0000011000110001; // vC= 1585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100011; // iC= 1123 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101011; // iC= 1131 
// vC = 14'b0000011001111111; // vC= 1663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010100; // iC=  980 
// vC = 14'b0000011001000101; // vC= 1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011100; // iC= 1052 
// vC = 14'b0000011101000101; // vC= 1861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100100; // iC=  996 
// vC = 14'b0000011100111100; // vC= 1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110000; // iC= 1200 
// vC = 14'b0000011001011111; // vC= 1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001000; // iC= 1160 
// vC = 14'b0000011001101100; // vC= 1644 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001110; // iC=  974 
// vC = 14'b0000011001000011; // vC= 1603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011101; // iC= 1053 
// vC = 14'b0000011010100010; // vC= 1698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001010; // iC= 1162 
// vC = 14'b0000011001101001; // vC= 1641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010010; // iC= 1042 
// vC = 14'b0000011011001100; // vC= 1740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100001; // iC=  993 
// vC = 14'b0000011001001110; // vC= 1614 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000000; // iC= 1152 
// vC = 14'b0000011001110001; // vC= 1649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100011; // iC=  931 
// vC = 14'b0000011100111001; // vC= 1849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110000; // iC=  944 
// vC = 14'b0000011010011010; // vC= 1690 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110110; // iC=  886 
// vC = 14'b0000011010001111; // vC= 1679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110010; // iC=  882 
// vC = 14'b0000011010111011; // vC= 1723 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101110; // iC= 1070 
// vC = 14'b0000011100001101; // vC= 1805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101100; // iC= 1132 
// vC = 14'b0000011110000010; // vC= 1922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101011; // iC=  939 
// vC = 14'b0000011100111010; // vC= 1850 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101001; // iC=  873 
// vC = 14'b0000011011001110; // vC= 1742 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011011; // iC=  923 
// vC = 14'b0000011101111111; // vC= 1919 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101001; // iC=  873 
// vC = 14'b0000011101101001; // vC= 1897 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000100; // iC=  964 
// vC = 14'b0000011100111010; // vC= 1850 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011100; // iC=  988 
// vC = 14'b0000011100110111; // vC= 1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101000; // iC=  936 
// vC = 14'b0000011101110010; // vC= 1906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010100; // iC= 1108 
// vC = 14'b0000011110100001; // vC= 1953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100010; // iC=  930 
// vC = 14'b0000011100010111; // vC= 1815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011000; // iC=  792 
// vC = 14'b0000011010111011; // vC= 1723 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011011; // iC=  795 
// vC = 14'b0000011110010100; // vC= 1940 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010111; // iC=  791 
// vC = 14'b0000011011100101; // vC= 1765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110101; // iC=  949 
// vC = 14'b0000011101011100; // vC= 1884 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011111; // iC=  799 
// vC = 14'b0000011011111011; // vC= 1787 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100101; // iC= 1061 
// vC = 14'b0000011011100011; // vC= 1763 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110000; // iC=  816 
// vC = 14'b0000011010100011; // vC= 1699 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111100; // iC=  892 
// vC = 14'b0000011011010101; // vC= 1749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010000; // iC=  912 
// vC = 14'b0000011100111001; // vC= 1849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110101; // iC=  885 
// vC = 14'b0000011011011101; // vC= 1757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001101; // iC=  845 
// vC = 14'b0000011100011000; // vC= 1816 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010000; // iC=  912 
// vC = 14'b0000011101001001; // vC= 1865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000001; // iC=  833 
// vC = 14'b0000011100111101; // vC= 1853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111001; // iC= 1017 
// vC = 14'b0000011101110011; // vC= 1907 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100000; // iC=  928 
// vC = 14'b0000011101101100; // vC= 1900 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101011; // iC=  747 
// vC = 14'b0000011100101000; // vC= 1832 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111100; // iC=  956 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001111; // iC=  911 
// vC = 14'b0000011010111111; // vC= 1727 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010011; // iC=  915 
// vC = 14'b0000011011001010; // vC= 1738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100111; // iC=  935 
// vC = 14'b0000011111001011; // vC= 1995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011100; // iC=  796 
// vC = 14'b0000011100100011; // vC= 1827 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000000; // iC=  832 
// vC = 14'b0000011100101111; // vC= 1839 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100111; // iC=  679 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110011; // iC=  947 
// vC = 14'b0000011011001001; // vC= 1737 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010001; // iC=  657 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111100; // iC=  892 
// vC = 14'b0000011111111000; // vC= 2040 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010001; // iC=  721 
// vC = 14'b0000011110111010; // vC= 1978 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111011; // iC=  891 
// vC = 14'b0000011011101110; // vC= 1774 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011110; // iC=  798 
// vC = 14'b0000011110110100; // vC= 1972 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011110; // iC=  926 
// vC = 14'b0000011101110111; // vC= 1911 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010011; // iC=  595 
// vC = 14'b0000011100111010; // vC= 1850 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001001; // iC=  841 
// vC = 14'b0000011111101010; // vC= 2026 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000100; // iC=  772 
// vC = 14'b0000011011110111; // vC= 1783 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100010; // iC=  674 
// vC = 14'b0000011100000100; // vC= 1796 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010000; // iC=  784 
// vC = 14'b0000011101011001; // vC= 1881 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000111; // iC=  647 
// vC = 14'b0000011101001001; // vC= 1865 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101111; // iC=  623 
// vC = 14'b0000011101000010; // vC= 1858 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011011; // iC=  603 
// vC = 14'b0000011100101110; // vC= 1838 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001001; // iC=  585 
// vC = 14'b0000011100000001; // vC= 1793 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111101; // iC=  701 
// vC = 14'b0000011111101111; // vC= 2031 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110001; // iC=  561 
// vC = 14'b0000011100101111; // vC= 1839 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101100; // iC=  812 
// vC = 14'b0000011110100111; // vC= 1959 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000001; // iC=  769 
// vC = 14'b0000011101001111; // vC= 1871 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111001; // iC=  825 
// vC = 14'b0000100000010000; // vC= 2064 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110111; // iC=  759 
// vC = 14'b0000011111010010; // vC= 2002 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010100; // iC=  660 
// vC = 14'b0000011111100001; // vC= 2017 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010010; // iC=  658 
// vC = 14'b0000011111000011; // vC= 1987 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001011; // iC=  715 
// vC = 14'b0000011100101010; // vC= 1834 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100011; // iC=  675 
// vC = 14'b0000011101001110; // vC= 1870 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101110; // iC=  494 
// vC = 14'b0000011101110100; // vC= 1908 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011110; // iC=  606 
// vC = 14'b0000100000001010; // vC= 2058 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011101; // iC=  605 
// vC = 14'b0000100000001100; // vC= 2060 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100100; // iC=  676 
// vC = 14'b0000100001000010; // vC= 2114 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001001; // iC=  521 
// vC = 14'b0000011111001111; // vC= 1999 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010100; // iC=  660 
// vC = 14'b0000011110111000; // vC= 1976 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001000; // iC=  520 
// vC = 14'b0000011101111101; // vC= 1917 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111011; // iC=  443 
// vC = 14'b0000011110000001; // vC= 1921 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000001; // iC=  449 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001001; // iC=  329 
// vC = 14'b0000011101011010; // vC= 1882 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011111; // iC=  607 
// vC = 14'b0000011111111011; // vC= 2043 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010000; // iC=  400 
// vC = 14'b0000011110001110; // vC= 1934 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010000; // iC=  400 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000110; // iC=  262 
// vC = 14'b0000100001011010; // vC= 2138 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010000; // iC=  528 
// vC = 14'b0000011111110001; // vC= 2033 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011110; // iC=  350 
// vC = 14'b0000100000010101; // vC= 2069 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001000; // iC=  456 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001101; // iC=  269 
// vC = 14'b0000011111100110; // vC= 2022 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011010; // iC=  410 
// vC = 14'b0000011110010010; // vC= 1938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100001; // iC=  161 
// vC = 14'b0000011111100001; // vC= 2017 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010101; // iC=  149 
// vC = 14'b0000100000010000; // vC= 2064 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000111; // iC=  327 
// vC = 14'b0000100001101111; // vC= 2159 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101100; // iC=  428 
// vC = 14'b0000100001001011; // vC= 2123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011110; // iC=  414 
// vC = 14'b0000100001010001; // vC= 2129 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110011; // iC=  371 
// vC = 14'b0000011110011011; // vC= 1947 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001101; // iC=   77 
// vC = 14'b0000011110101101; // vC= 1965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100010; // iC=  226 
// vC = 14'b0000100001010101; // vC= 2133 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000010; // iC=  194 
// vC = 14'b0000011100111111; // vC= 1855 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101011; // iC=   43 
// vC = 14'b0000011110000100; // vC= 1924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110100; // iC=  244 
// vC = 14'b0000100001001010; // vC= 2122 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100010; // iC=   98 
// vC = 14'b0000100001100010; // vC= 2146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000011; // iC=  195 
// vC = 14'b0000100000100110; // vC= 2086 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100110; // iC=  230 
// vC = 14'b0000011101010011; // vC= 1875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100101; // iC=  101 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100101; // iC=  101 
// vC = 14'b0000100001101100; // vC= 2156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000000; // iC=    0 
// vC = 14'b0000011101111101; // vC= 1917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001000; // iC= -120 
// vC = 14'b0000011111110010; // vC= 2034 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011011; // iC=  155 
// vC = 14'b0000011101110011; // vC= 1907 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100100; // iC=  -28 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111101; // iC=   -3 
// vC = 14'b0000011110111011; // vC= 1979 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011010; // iC=   26 
// vC = 14'b0000100000010011; // vC= 2067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110010; // iC= -206 
// vC = 14'b0000100001100010; // vC= 2146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010100; // iC=  -44 
// vC = 14'b0000011111000001; // vC= 1985 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100011; // iC=  -29 
// vC = 14'b0000011101101010; // vC= 1898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111000; // iC= -200 
// vC = 14'b0000100000000110; // vC= 2054 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010011; // iC= -109 
// vC = 14'b0000100000100010; // vC= 2082 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100111; // iC= -153 
// vC = 14'b0000011101110011; // vC= 1907 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011001; // iC= -231 
// vC = 14'b0000011110111010; // vC= 1978 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110000; // iC= -208 
// vC = 14'b0000011111111000; // vC= 2040 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110111; // iC= -329 
// vC = 14'b0000011101111111; // vC= 1919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011110101; // iC= -267 
// vC = 14'b0000011110010001; // vC= 1937 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011101; // iC= -355 
// vC = 14'b0000011110100100; // vC= 1956 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101000; // iC= -280 
// vC = 14'b0000011111001001; // vC= 1993 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111100; // iC= -196 
// vC = 14'b0000100000101011; // vC= 2091 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000101; // iC= -315 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100000; // iC= -544 
// vC = 14'b0000100000010011; // vC= 2067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001011; // iC= -565 
// vC = 14'b0000011111100100; // vC= 2020 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110100; // iC= -588 
// vC = 14'b0000011101001000; // vC= 1864 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100111; // iC= -601 
// vC = 14'b0000011111110101; // vC= 2037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011111; // iC= -353 
// vC = 14'b0000011110101100; // vC= 1964 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001110; // iC= -626 
// vC = 14'b0000100001000011; // vC= 2115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000000; // iC= -448 
// vC = 14'b0000100001010011; // vC= 2131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101001; // iC= -663 
// vC = 14'b0000011100101111; // vC= 1839 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001110; // iC= -498 
// vC = 14'b0000011110000001; // vC= 1921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100010; // iC= -670 
// vC = 14'b0000011110100110; // vC= 1958 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100001; // iC= -543 
// vC = 14'b0000011111111011; // vC= 2043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011101; // iC= -547 
// vC = 14'b0000011110100001; // vC= 1953 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101111; // iC= -721 
// vC = 14'b0000011101100111; // vC= 1895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010011; // iC= -621 
// vC = 14'b0000011111110011; // vC= 2035 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011101; // iC= -803 
// vC = 14'b0000011100110001; // vC= 1841 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001111; // iC= -817 
// vC = 14'b0000011101000100; // vC= 1860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010010; // iC= -750 
// vC = 14'b0000011110111000; // vC= 1976 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111110; // iC= -962 
// vC = 14'b0000100000101110; // vC= 2094 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110011; // iC= -845 
// vC = 14'b0000011111100001; // vC= 2017 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011010; // iC= -998 
// vC = 14'b0000011111110000; // vC= 2032 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001010; // iC= -822 
// vC = 14'b0000011100100010; // vC= 1826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110101; // iC= -843 
// vC = 14'b0000011011100100; // vC= 1764 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110010; // iC= -846 
// vC = 14'b0000011110111010; // vC= 1978 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b0000011011101011; // vC= 1771 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100011; // iC= -989 
// vC = 14'b0000011101001010; // vC= 1866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100111; // iC= -921 
// vC = 14'b0000011011110100; // vC= 1780 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101000; // iC= -920 
// vC = 14'b0000011011100001; // vC= 1761 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111101; // iC=-1091 
// vC = 14'b0000011100111011; // vC= 1851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111101; // iC=-1027 
// vC = 14'b0000011100110110; // vC= 1846 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111111; // iC=-1153 
// vC = 14'b0000011011111011; // vC= 1787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001010; // iC=-1078 
// vC = 14'b0000011111001110; // vC= 1998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011000; // iC=-1192 
// vC = 14'b0000011011101010; // vC= 1770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011101; // iC=-1187 
// vC = 14'b0000011101001111; // vC= 1871 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111011; // iC=-1029 
// vC = 14'b0000011010100110; // vC= 1702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001000; // iC=-1144 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110001; // iC=-1039 
// vC = 14'b0000011010100100; // vC= 1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011101; // iC=-1315 
// vC = 14'b0000011011111000; // vC= 1784 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000110; // iC=-1082 
// vC = 14'b0000011011000011; // vC= 1731 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110010; // iC=-1102 
// vC = 14'b0000011100010000; // vC= 1808 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111110; // iC=-1154 
// vC = 14'b0000011101111111; // vC= 1919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011110; // iC=-1186 
// vC = 14'b0000011010101101; // vC= 1709 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100011; // iC=-1245 
// vC = 14'b0000011110110100; // vC= 1972 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001011; // iC=-1333 
// vC = 14'b0000011011100111; // vC= 1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110111; // iC=-1225 
// vC = 14'b0000011011001111; // vC= 1743 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100101; // iC=-1371 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111000; // iC=-1416 
// vC = 14'b0000011011100110; // vC= 1766 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010010; // iC=-1454 
// vC = 14'b0000011010011000; // vC= 1688 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001000; // iC=-1400 
// vC = 14'b0000011001010111; // vC= 1623 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010011; // iC=-1325 
// vC = 14'b0000011101011100; // vC= 1884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010110; // iC=-1386 
// vC = 14'b0000011100001110; // vC= 1806 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000000; // iC=-1536 
// vC = 14'b0000011010111111; // vC= 1727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000000; // iC=-1408 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010111; // iC=-1641 
// vC = 14'b0000011100101001; // vC= 1833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101010; // iC=-1494 
// vC = 14'b0000011100110100; // vC= 1844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010010; // iC=-1454 
// vC = 14'b0000011001011010; // vC= 1626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011010; // iC=-1382 
// vC = 14'b0000011001110101; // vC= 1653 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111010; // iC=-1478 
// vC = 14'b0000011001101101; // vC= 1645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100010; // iC=-1438 
// vC = 14'b0000011101010011; // vC= 1875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011101; // iC=-1507 
// vC = 14'b0000011100011101; // vC= 1821 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101110; // iC=-1426 
// vC = 14'b0000011100001010; // vC= 1802 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010011; // iC=-1581 
// vC = 14'b0000011010000100; // vC= 1668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010110; // iC=-1770 
// vC = 14'b0000011010011100; // vC= 1692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010110; // iC=-1642 
// vC = 14'b0000011001101101; // vC= 1645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101101; // iC=-1619 
// vC = 14'b0000011001011010; // vC= 1626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b0000011000111000; // vC= 1592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011011; // iC=-1509 
// vC = 14'b0000011000110100; // vC= 1588 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101011; // iC=-1749 
// vC = 14'b0000011000010101; // vC= 1557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b0000011000000011; // vC= 1539 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110001; // iC=-1743 
// vC = 14'b0000011000110011; // vC= 1587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001001; // iC=-1591 
// vC = 14'b0000011000000100; // vC= 1540 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101100; // iC=-1684 
// vC = 14'b0000011011100010; // vC= 1762 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101110; // iC=-1682 
// vC = 14'b0000011001001001; // vC= 1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001101; // iC=-1907 
// vC = 14'b0000010110110111; // vC= 1463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001110; // iC=-1714 
// vC = 14'b0000011001101100; // vC= 1644 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110101; // iC=-1675 
// vC = 14'b0000010111110101; // vC= 1525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b0000011000101010; // vC= 1578 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b0000011010001001; // vC= 1673 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110000; // iC=-1936 
// vC = 14'b0000011010100100; // vC= 1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001101; // iC=-1651 
// vC = 14'b0000011010011011; // vC= 1691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101000; // iC=-1816 
// vC = 14'b0000010110110111; // vC= 1463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000011; // iC=-1725 
// vC = 14'b0000010110010000; // vC= 1424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010101; // iC=-1771 
// vC = 14'b0000011001010110; // vC= 1622 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001110; // iC=-1714 
// vC = 14'b0000011000011011; // vC= 1563 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000100; // iC=-1980 
// vC = 14'b0000011000011110; // vC= 1566 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b0000010101001111; // vC= 1359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b0000011000100010; // vC= 1570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b0000010101100100; // vC= 1380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b0000010100101111; // vC= 1327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b0000010101111000; // vC= 1400 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000011001010100; // vC= 1620 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110011; // iC=-1869 
// vC = 14'b0000010110011110; // vC= 1438 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b0000010110000010; // vC= 1410 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b0000011000010000; // vC= 1552 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101111; // iC=-1873 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b0000011000100010; // vC= 1570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010000; // iC=-2096 
// vC = 14'b0000010101001011; // vC= 1355 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b0000010011100010; // vC= 1250 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011101; // iC=-1827 
// vC = 14'b0000010111100110; // vC= 1510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b0000010101010110; // vC= 1366 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b0000010101100101; // vC= 1381 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111110; // iC=-1922 
// vC = 14'b0000010101101000; // vC= 1384 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000010100100000; // vC= 1312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010110; // iC=-1834 
// vC = 14'b0000010110011000; // vC= 1432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100011; // iC=-1949 
// vC = 14'b0000010101101001; // vC= 1385 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b0000010011010011; // vC= 1235 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000010011011011; // vC= 1243 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b0000010101100100; // vC= 1380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b0000010100001100; // vC= 1292 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b0000010100101011; // vC= 1323 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011100; // iC=-1892 
// vC = 14'b0000010101110000; // vC= 1392 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b0000010100101010; // vC= 1322 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b0000010101111111; // vC= 1407 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010111; // iC=-2153 
// vC = 14'b0000010010001010; // vC= 1162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010011; // iC=-2093 
// vC = 14'b0000010010100011; // vC= 1187 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b0000010101101110; // vC= 1390 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111001; // iC=-1991 
// vC = 14'b0000010010100000; // vC= 1184 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b0000010100000110; // vC= 1286 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010000; // iC=-1968 
// vC = 14'b0000010101001110; // vC= 1358 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b0000010011001000; // vC= 1224 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b0000010100110111; // vC= 1335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b0000010010010100; // vC= 1172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010101; // iC=-2155 
// vC = 14'b0000010010101100; // vC= 1196 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b0000010100100101; // vC= 1317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b0000010011100100; // vC= 1252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000100; // iC=-1916 
// vC = 14'b0000010011111100; // vC= 1276 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001011; // iC=-2165 
// vC = 14'b0000010100011000; // vC= 1304 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101101; // iC=-2195 
// vC = 14'b0000001111010111; // vC=  983 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000110; // iC=-1978 
// vC = 14'b0000010000010111; // vC= 1047 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010001; // iC=-2031 
// vC = 14'b0000010010010001; // vC= 1169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b0000010010010111; // vC= 1175 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b0000001111001001; // vC=  969 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000010010000011; // vC= 1155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101100; // iC=-2068 
// vC = 14'b0000001111000000; // vC=  960 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111011; // iC=-2117 
// vC = 14'b0000010010010110; // vC= 1174 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b0000010010100111; // vC= 1191 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111111; // iC=-2113 
// vC = 14'b0000010000001111; // vC= 1039 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b0000010010110100; // vC= 1204 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010010; // iC=-2094 
// vC = 14'b0000001111110000; // vC= 1008 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b0000010000001011; // vC= 1035 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000010001100001; // vC= 1121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011111; // iC=-2081 
// vC = 14'b0000001111011011; // vC=  987 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b0000001111010110; // vC=  982 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000010001100011; // vC= 1123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b0000010000110011; // vC= 1075 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b0000001110010110; // vC=  918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011100; // iC=-2148 
// vC = 14'b0000001110111001; // vC=  953 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000001111001111; // vC=  975 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001110; // iC=-2162 
// vC = 14'b0000001100101010; // vC=  810 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110010; // iC=-2190 
// vC = 14'b0000001100001011; // vC=  779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111101; // iC=-2179 
// vC = 14'b0000001111000111; // vC=  967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000001110101101; // vC=  941 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110000; // iC=-1936 
// vC = 14'b0000001100011100; // vC=  796 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011010; // iC=-2214 
// vC = 14'b0000001111000101; // vC=  965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b0000001110101010; // vC=  938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111111; // iC=-2177 
// vC = 14'b0000001110111111; // vC=  959 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000001101000010; // vC=  834 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b0000001111011111; // vC=  991 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000001; // iC=-2239 
// vC = 14'b0000001100111011; // vC=  827 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000010; // iC=-1918 
// vC = 14'b0000001010111100; // vC=  700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010111; // iC=-2153 
// vC = 14'b0000001011011000; // vC=  728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001101; // iC=-2163 
// vC = 14'b0000001011000100; // vC=  708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011101; // iC=-2211 
// vC = 14'b0000001110011100; // vC=  924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010011; // iC=-2157 
// vC = 14'b0000001011001000; // vC=  712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111000; // iC=-2120 
// vC = 14'b0000001100100101; // vC=  805 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001110; // iC=-2226 
// vC = 14'b0000001011001000; // vC=  712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000110; // iC=-1978 
// vC = 14'b0000001010000110; // vC=  646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000001010011111; // vC=  671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000110; // iC=-2170 
// vC = 14'b0000001001100000; // vC=  608 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b0000001100001110; // vC=  782 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110101; // iC=-2187 
// vC = 14'b0000001101101101; // vC=  877 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011110; // iC=-2082 
// vC = 14'b0000001010010100; // vC=  660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001101; // iC=-2035 
// vC = 14'b0000001011010001; // vC=  721 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000001101010010; // vC=  850 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000001010110100; // vC=  692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100110; // iC=-2138 
// vC = 14'b0000001010000100; // vC=  644 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100100; // iC=-2140 
// vC = 14'b0000001100011000; // vC=  792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100101; // iC=-2139 
// vC = 14'b0000001100011000; // vC=  792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100011; // iC=-2141 
// vC = 14'b0000001100110000; // vC=  816 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010010; // iC=-1966 
// vC = 14'b0000001000101001; // vC=  553 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101110; // iC=-2194 
// vC = 14'b0000001011010000; // vC=  720 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000010; // iC=-2238 
// vC = 14'b0000001010001110; // vC=  654 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010001; // iC=-2223 
// vC = 14'b0000000111100101; // vC=  485 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001001; // iC=-2103 
// vC = 14'b0000001011010011; // vC=  723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011001; // iC=-2215 
// vC = 14'b0000001000111110; // vC=  574 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b0000001000101100; // vC=  556 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b0000001000000010; // vC=  514 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100111; // iC=-2073 
// vC = 14'b0000001001000101; // vC=  581 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b0000001001100010; // vC=  610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100110; // iC=-2202 
// vC = 14'b0000000110111111; // vC=  447 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000001001000110; // vC=  582 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101100; // iC=-2132 
// vC = 14'b0000001000011111; // vC=  543 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b0000000110101100; // vC=  428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000001001111010; // vC=  634 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100010; // iC=-2206 
// vC = 14'b0000001001001101; // vC=  589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b0000000111110010; // vC=  498 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101010; // iC=-2070 
// vC = 14'b0000000101111010; // vC=  378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000000110011111; // vC=  415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100100; // iC=-1948 
// vC = 14'b0000000111000011; // vC=  451 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000001; // iC=-2175 
// vC = 14'b0000001001101001; // vC=  617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001001; // iC=-2231 
// vC = 14'b0000000101001011; // vC=  331 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b0000001001011100; // vC=  604 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100101; // iC=-2075 
// vC = 14'b0000001000000110; // vC=  518 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100110; // iC=-2074 
// vC = 14'b0000000111100011; // vC=  483 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011110; // iC=-2210 
// vC = 14'b0000001000001000; // vC=  520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110000; // iC=-2256 
// vC = 14'b0000000111101111; // vC=  495 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000000011101110; // vC=  238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110011; // iC=-2125 
// vC = 14'b0000000011100100; // vC=  228 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000001000001011; // vC=  523 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110011; // iC=-2253 
// vC = 14'b0000000110001110; // vC=  398 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b0000000101001110; // vC=  334 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000100; // iC=-2236 
// vC = 14'b0000000110100001; // vC=  417 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110110; // iC=-2122 
// vC = 14'b0000000100001000; // vC=  264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b0000000011001001; // vC=  201 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b0000000011011001; // vC=  217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101000; // iC=-2136 
// vC = 14'b0000000101000100; // vC=  324 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100111; // iC=-2137 
// vC = 14'b0000000111000110; // vC=  454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b0000000010011101; // vC=  157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111110; // iC=-2242 
// vC = 14'b0000000011100100; // vC=  228 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b0000000110100101; // vC=  421 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011100; // iC=-2212 
// vC = 14'b0000000011110101; // vC=  245 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010111; // iC=-2089 
// vC = 14'b0000000001110100; // vC=  116 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b0000000101011010; // vC=  346 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111111; // iC=-2241 
// vC = 14'b0000000011010001; // vC=  209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b0000000001001111; // vC=   79 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000000; // iC=-2240 
// vC = 14'b0000000101011000; // vC=  344 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100110; // iC=-2202 
// vC = 14'b0000000100010110; // vC=  278 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111111; // iC=-2113 
// vC = 14'b0000000001111101; // vC=  125 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100000; // iC=-2208 
// vC = 14'b0000000011011001; // vC=  217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011111; // iC=-2209 
// vC = 14'b0000000100100010; // vC=  290 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b0000000101011010; // vC=  346 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b0000000010100001; // vC=  161 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110010; // iC=-2190 
// vC = 14'b0000000100001010; // vC=  266 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010110; // iC=-2218 
// vC = 14'b0000000011100110; // vC=  230 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110110; // iC=-2122 
// vC = 14'b0000000001100101; // vC=  101 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000100; // iC=-2172 
// vC = 14'b0000000100100111; // vC=  295 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000011; // iC=-1981 
// vC = 14'b1111111111111010; // vC=   -6 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110111; // iC=-2185 
// vC = 14'b0000000010100110; // vC=  166 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110001; // iC=-2127 
// vC = 14'b0000000000001010; // vC=   10 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b1111111111010110; // vC=  -42 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010000; // iC=-2224 
// vC = 14'b0000000010011001; // vC=  153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001101; // iC=-2099 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101100; // iC=-2068 
// vC = 14'b0000000000011000; // vC=   24 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001100; // iC=-2164 
// vC = 14'b0000000000100011; // vC=   35 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110101; // iC=-2123 
// vC = 14'b1111111110100011; // vC=  -93 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b0000000011001001; // vC=  201 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001010; // iC=-2166 
// vC = 14'b0000000011000100; // vC=  196 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b1111111110100111; // vC=  -89 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b1111111110111011; // vC=  -69 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110100; // iC=-2188 
// vC = 14'b1111111101111001; // vC= -135 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b1111111111100101; // vC=  -27 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000000001111111; // vC=  127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000101; // iC=-2171 
// vC = 14'b1111111111101101; // vC=  -19 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100011; // iC=-2141 
// vC = 14'b1111111110100100; // vC=  -92 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010111; // iC=-2025 
// vC = 14'b1111111110111010; // vC=  -70 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100000; // iC=-2016 
// vC = 14'b1111111111100011; // vC=  -29 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b0000000001011011; // vC=   91 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000111; // iC=-2105 
// vC = 14'b1111111111011100; // vC=  -36 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100010; // iC=-2014 
// vC = 14'b1111111101000111; // vC= -185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b1111111101101101; // vC= -147 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b1111111101100001; // vC= -159 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011010; // iC=-2150 
// vC = 14'b1111111111001110; // vC=  -50 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101001; // iC=-2135 
// vC = 14'b1111111100010111; // vC= -233 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010000; // iC=-2160 
// vC = 14'b1111111111010100; // vC=  -44 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b1111111111001011; // vC=  -53 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000101; // iC=-2043 
// vC = 14'b1111111111100000; // vC=  -32 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b1111111111110100; // vC=  -12 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b1111111100111111; // vC= -193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b1111111100011111; // vC= -225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001111; // iC=-2161 
// vC = 14'b1111111100001111; // vC= -241 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b1111111110001001; // vC= -119 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b1111111101110111; // vC= -137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101110; // iC=-1874 
// vC = 14'b1111111101010101; // vC= -171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111110; // iC=-2050 
// vC = 14'b1111111101011001; // vC= -167 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b1111111100011110; // vC= -226 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010011; // iC=-2157 
// vC = 14'b1111111100111101; // vC= -195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000010; // iC=-2174 
// vC = 14'b1111111100111110; // vC= -194 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101011; // iC=-2133 
// vC = 14'b1111111010111101; // vC= -323 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b1111111010110101; // vC= -331 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010110; // iC=-1898 
// vC = 14'b1111111100110010; // vC= -206 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001000; // iC=-2040 
// vC = 14'b1111111101011101; // vC= -163 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000100; // iC=-1852 
// vC = 14'b1111111010100001; // vC= -351 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b1111111010110101; // vC= -331 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b1111111010100011; // vC= -349 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110100; // iC=-1932 
// vC = 14'b1111111001110110; // vC= -394 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b1111111101110001; // vC= -143 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b1111111101101000; // vC= -152 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001101; // iC=-1907 
// vC = 14'b1111111101100101; // vC= -155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000100; // iC=-1852 
// vC = 14'b1111111000110001; // vC= -463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b1111111010110111; // vC= -329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b1111111010100111; // vC= -345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000100; // iC=-2108 
// vC = 14'b1111111000000000; // vC= -512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011110; // iC=-1826 
// vC = 14'b1111111001010101; // vC= -427 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b1111111001111110; // vC= -386 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b1111111001100101; // vC= -411 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010111; // iC=-1833 
// vC = 14'b1111111011010010; // vC= -302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111110111100100; // vC= -540 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110010; // iC=-1934 
// vC = 14'b1111111010001001; // vC= -375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111100; // iC=-1924 
// vC = 14'b1111111001011100; // vC= -420 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000111; // iC=-2105 
// vC = 14'b1111110111001101; // vC= -563 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010101; // iC=-1835 
// vC = 14'b1111111011100010; // vC= -286 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110100; // iC=-1804 
// vC = 14'b1111110111011001; // vC= -551 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b1111111011010001; // vC= -303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100010; // iC=-1886 
// vC = 14'b1111111010110111; // vC= -329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b1111111000000101; // vC= -507 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b1111111001100101; // vC= -411 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b1111111010111001; // vC= -327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001010; // iC=-1846 
// vC = 14'b1111111001101110; // vC= -402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111001; // iC=-1799 
// vC = 14'b1111111001101100; // vC= -404 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100010; // iC=-2014 
// vC = 14'b1111111001001100; // vC= -436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111111; // iC=-2049 
// vC = 14'b1111111001010101; // vC= -427 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b1111111001000111; // vC= -441 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b1111110101101011; // vC= -661 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100011; // iC=-2077 
// vC = 14'b1111110111011011; // vC= -549 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101111; // iC=-2001 
// vC = 14'b1111110111001101; // vC= -563 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111111; // iC=-2049 
// vC = 14'b1111111000111100; // vC= -452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011001; // iC=-1767 
// vC = 14'b1111110110000010; // vC= -638 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010010; // iC=-1774 
// vC = 14'b1111110111101101; // vC= -531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b1111111000010001; // vC= -495 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b1111110110001001; // vC= -631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b1111110110101101; // vC= -595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100001; // iC=-1759 
// vC = 14'b1111111000011100; // vC= -484 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001101; // iC=-1907 
// vC = 14'b1111110110001010; // vC= -630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010001; // iC=-1775 
// vC = 14'b1111111000110111; // vC= -457 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110101; // iC=-1739 
// vC = 14'b1111111000010110; // vC= -490 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010001; // iC=-2031 
// vC = 14'b1111110110100110; // vC= -602 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100011; // iC=-1821 
// vC = 14'b1111110100001111; // vC= -753 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111011; // iC=-1733 
// vC = 14'b1111110111100110; // vC= -538 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b1111110110111111; // vC= -577 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b1111110111001001; // vC= -567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b1111111000000010; // vC= -510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001000; // iC=-2040 
// vC = 14'b1111110111110110; // vC= -522 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101111; // iC=-1809 
// vC = 14'b1111110111100101; // vC= -539 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b1111110011100110; // vC= -794 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000111; // iC=-1785 
// vC = 14'b1111110110101110; // vC= -594 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100011; // iC=-1821 
// vC = 14'b1111110010111010; // vC= -838 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000000; // iC=-1728 
// vC = 14'b1111110110011110; // vC= -610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110010; // iC=-1870 
// vC = 14'b1111110101111001; // vC= -647 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b1111110101001010; // vC= -694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001100; // iC=-1716 
// vC = 14'b1111110101100100; // vC= -668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001001; // iC=-1783 
// vC = 14'b1111110011100111; // vC= -793 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b1111110010011110; // vC= -866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100000; // iC=-1760 
// vC = 14'b1111110001100111; // vC= -921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000110; // iC=-1850 
// vC = 14'b1111110100100001; // vC= -735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b1111110100100100; // vC= -732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b1111110001110001; // vC= -911 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001110; // iC=-1714 
// vC = 14'b1111110100111111; // vC= -705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010001; // iC=-1839 
// vC = 14'b1111110101110000; // vC= -656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b1111110000111101; // vC= -963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001101; // iC=-1907 
// vC = 14'b1111110101100101; // vC= -667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111111; // iC=-1921 
// vC = 14'b1111110001110001; // vC= -911 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110110; // iC=-1674 
// vC = 14'b1111110001000001; // vC= -959 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b1111110011000011; // vC= -829 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b1111110100010000; // vC= -752 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001001; // iC=-1719 
// vC = 14'b1111110000100101; // vC= -987 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001010; // iC=-1718 
// vC = 14'b1111110011000000; // vC= -832 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b1111110001011100; // vC= -932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111111; // iC=-1729 
// vC = 14'b1111110011010111; // vC= -809 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100111; // iC=-1817 
// vC = 14'b1111110010001001; // vC= -887 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011011; // iC=-1829 
// vC = 14'b1111110011011011; // vC= -805 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111111; // iC=-1793 
// vC = 14'b1111110010111111; // vC= -833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001000; // iC=-1720 
// vC = 14'b1111110000101100; // vC= -980 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b1111110010010000; // vC= -880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001100; // iC=-1780 
// vC = 14'b1111110000111011; // vC= -965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010110; // iC=-1642 
// vC = 14'b1111110000101010; // vC= -982 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001101; // iC=-1651 
// vC = 14'b1111110011100101; // vC= -795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100101; // iC=-1755 
// vC = 14'b1111110011001101; // vC= -819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001010; // iC=-1782 
// vC = 14'b1111110010010000; // vC= -880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111101; // iC=-1667 
// vC = 14'b1111110010011110; // vC= -866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111011; // iC=-1605 
// vC = 14'b1111110000100101; // vC= -987 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b1111101111000010; // vC=-1086 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010000; // iC=-1648 
// vC = 14'b1111101110011100; // vC=-1124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011011; // iC=-1573 
// vC = 14'b1111110001100101; // vC= -923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111010; // iC=-1670 
// vC = 14'b1111110000010101; // vC=-1003 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110001; // iC=-1679 
// vC = 14'b1111101111100101; // vC=-1051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b1111101111001011; // vC=-1077 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010100; // iC=-1580 
// vC = 14'b1111101111011111; // vC=-1057 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011001; // iC=-1575 
// vC = 14'b1111110001010110; // vC= -938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011100; // iC=-1700 
// vC = 14'b1111110000111101; // vC= -963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000110; // iC=-1594 
// vC = 14'b1111110010001001; // vC= -887 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101000; // iC=-1624 
// vC = 14'b1111101111100101; // vC=-1051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000101; // iC=-1595 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110111; // iC=-1673 
// vC = 14'b1111110001010110; // vC= -938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010100; // iC=-1772 
// vC = 14'b1111110001001110; // vC= -946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100101; // iC=-1819 
// vC = 14'b1111101100101110; // vC=-1234 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100110; // iC=-1626 
// vC = 14'b1111101100101011; // vC=-1237 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010101; // iC=-1643 
// vC = 14'b1111110001010110; // vC= -938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110010; // iC=-1678 
// vC = 14'b1111101110011100; // vC=-1124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000010; // iC=-1598 
// vC = 14'b1111101100011100; // vC=-1252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010111; // iC=-1769 
// vC = 14'b1111101110001011; // vC=-1141 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b1111101100000011; // vC=-1277 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010011; // iC=-1581 
// vC = 14'b1111101100000000; // vC=-1280 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010011; // iC=-1773 
// vC = 14'b1111101110111010; // vC=-1094 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111100; // iC=-1796 
// vC = 14'b1111101101001100; // vC=-1204 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111110; // iC=-1666 
// vC = 14'b1111101101101101; // vC=-1171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110000; // iC=-1488 
// vC = 14'b1111101110011110; // vC=-1122 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110111; // iC=-1545 
// vC = 14'b1111101111011110; // vC=-1058 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110001; // iC=-1551 
// vC = 14'b1111101100101010; // vC=-1238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010110; // iC=-1642 
// vC = 14'b1111101110101111; // vC=-1105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000010; // iC=-1726 
// vC = 14'b1111101101111101; // vC=-1155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011001; // iC=-1639 
// vC = 14'b1111101101001011; // vC=-1205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011111; // iC=-1505 
// vC = 14'b1111101111010101; // vC=-1067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101111; // iC=-1745 
// vC = 14'b1111101101011100; // vC=-1188 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111111; // iC=-1473 
// vC = 14'b1111101010100101; // vC=-1371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110000; // iC=-1552 
// vC = 14'b1111101100001111; // vC=-1265 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111010; // iC=-1734 
// vC = 14'b1111101100011110; // vC=-1250 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101010; // iC=-1558 
// vC = 14'b1111101110001001; // vC=-1143 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100100; // iC=-1692 
// vC = 14'b1111101110110011; // vC=-1101 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111011; // iC=-1413 
// vC = 14'b1111101011111100; // vC=-1284 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101010; // iC=-1558 
// vC = 14'b1111101110001001; // vC=-1143 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100011; // iC=-1629 
// vC = 14'b1111101001110111; // vC=-1417 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010100; // iC=-1644 
// vC = 14'b1111101010100111; // vC=-1369 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111111; // iC=-1665 
// vC = 14'b1111101010101011; // vC=-1365 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011110; // iC=-1506 
// vC = 14'b1111101100000010; // vC=-1278 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011000; // iC=-1640 
// vC = 14'b1111101110100000; // vC=-1120 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001011; // iC=-1397 
// vC = 14'b1111101101111100; // vC=-1156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000011; // iC=-1661 
// vC = 14'b1111101100000100; // vC=-1276 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100100; // iC=-1500 
// vC = 14'b1111101101001011; // vC=-1205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010010; // iC=-1518 
// vC = 14'b1111101100010000; // vC=-1264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101111; // iC=-1425 
// vC = 14'b1111101001010100; // vC=-1452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010111; // iC=-1577 
// vC = 14'b1111101101001100; // vC=-1204 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111110; // iC=-1602 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000011; // iC=-1405 
// vC = 14'b1111101000111001; // vC=-1479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000000; // iC=-1536 
// vC = 14'b1111101001100010; // vC=-1438 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011001; // iC=-1447 
// vC = 14'b1111101010100001; // vC=-1375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110111; // iC=-1545 
// vC = 14'b1111101011111100; // vC=-1284 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100101; // iC=-1499 
// vC = 14'b1111101010000111; // vC=-1401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011100; // iC=-1508 
// vC = 14'b1111101011100111; // vC=-1305 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111000; // iC=-1352 
// vC = 14'b1111101001110100; // vC=-1420 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011110; // iC=-1570 
// vC = 14'b1111101010100011; // vC=-1373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101101; // iC=-1555 
// vC = 14'b1111101001010000; // vC=-1456 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100010; // iC=-1566 
// vC = 14'b1111101000000010; // vC=-1534 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100100; // iC=-1500 
// vC = 14'b1111101010110010; // vC=-1358 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100011; // iC=-1565 
// vC = 14'b1111101000111001; // vC=-1479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110111; // iC=-1545 
// vC = 14'b1111101011011101; // vC=-1315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001001; // iC=-1399 
// vC = 14'b1111101010101100; // vC=-1364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011100; // iC=-1572 
// vC = 14'b1111101010011011; // vC=-1381 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000010; // iC=-1534 
// vC = 14'b1111101010000111; // vC=-1401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001100; // iC=-1524 
// vC = 14'b1111101011000001; // vC=-1343 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000100; // iC=-1404 
// vC = 14'b1111101000000110; // vC=-1530 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101100; // iC=-1492 
// vC = 14'b1111101001100001; // vC=-1439 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100110; // iC=-1306 
// vC = 14'b1111101001101010; // vC=-1430 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111100; // iC=-1476 
// vC = 14'b1111101000001111; // vC=-1521 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100100; // iC=-1308 
// vC = 14'b1111100111110101; // vC=-1547 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111001; // iC=-1543 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010110; // iC=-1450 
// vC = 14'b1111101011001011; // vC=-1333 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001000; // iC=-1464 
// vC = 14'b1111101010001100; // vC=-1396 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011110; // iC=-1378 
// vC = 14'b1111101001000010; // vC=-1470 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111011; // iC=-1285 
// vC = 14'b1111101010110110; // vC=-1354 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111100; // iC=-1348 
// vC = 14'b1111101011000100; // vC=-1340 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101111; // iC=-1489 
// vC = 14'b1111101000110011; // vC=-1485 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011100; // iC=-1508 
// vC = 14'b1111100110011111; // vC=-1633 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010001; // iC=-1199 
// vC = 14'b1111100111000100; // vC=-1596 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000111; // iC=-1209 
// vC = 14'b1111100111011111; // vC=-1569 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000011; // iC=-1405 
// vC = 14'b1111101000111100; // vC=-1476 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101111; // iC=-1233 
// vC = 14'b1111101010011101; // vC=-1379 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010111; // iC=-1257 
// vC = 14'b1111101001001001; // vC=-1463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100001; // iC=-1247 
// vC = 14'b1111100110010110; // vC=-1642 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011100; // iC=-1316 
// vC = 14'b1111101010010101; // vC=-1387 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001000; // iC=-1272 
// vC = 14'b1111100111101111; // vC=-1553 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010101; // iC=-1451 
// vC = 14'b1111101001100011; // vC=-1437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010001; // iC=-1455 
// vC = 14'b1111100111101110; // vC=-1554 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000101; // iC=-1403 
// vC = 14'b1111100111011011; // vC=-1573 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001000; // iC=-1336 
// vC = 14'b1111100111010001; // vC=-1583 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010100; // iC=-1132 
// vC = 14'b1111100110000010; // vC=-1662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011011; // iC=-1253 
// vC = 14'b1111100101010100; // vC=-1708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000100; // iC=-1276 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001001; // iC=-1335 
// vC = 14'b1111101000000001; // vC=-1535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110000; // iC=-1360 
// vC = 14'b1111100101111101; // vC=-1667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101001; // iC=-1239 
// vC = 14'b1111100110100001; // vC=-1631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000100; // iC=-1404 
// vC = 14'b1111100111011010; // vC=-1574 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000110; // iC=-1210 
// vC = 14'b1111100111011110; // vC=-1570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110111; // iC=-1289 
// vC = 14'b1111101000100100; // vC=-1500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101011; // iC=-1365 
// vC = 14'b1111100110000111; // vC=-1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011101; // iC=-1315 
// vC = 14'b1111100110111000; // vC=-1608 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101111; // iC=-1169 
// vC = 14'b1111100101000110; // vC=-1722 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100101; // iC=-1179 
// vC = 14'b1111100100110101; // vC=-1739 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011101; // iC=-1187 
// vC = 14'b1111100100111110; // vC=-1730 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001011; // iC=-1141 
// vC = 14'b1111101000011111; // vC=-1505 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101001; // iC=-1111 
// vC = 14'b1111100110010011; // vC=-1645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110010; // iC=-1166 
// vC = 14'b1111100111001011; // vC=-1589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101000; // iC=-1304 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010010; // iC=-1070 
// vC = 14'b1111100011110100; // vC=-1804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110011; // iC=-1293 
// vC = 14'b1111101000000010; // vC=-1534 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010001; // iC=-1135 
// vC = 14'b1111100101010110; // vC=-1706 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110011; // iC=-1101 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010101; // iC=-1259 
// vC = 14'b1111100101010110; // vC=-1706 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b1111100111100111; // vC=-1561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111111; // iC=-1217 
// vC = 14'b1111100100010001; // vC=-1775 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010101; // iC=-1131 
// vC = 14'b1111100011100100; // vC=-1820 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000001; // iC=-1151 
// vC = 14'b1111100101011001; // vC=-1703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011101; // iC=-1123 
// vC = 14'b1111100101011011; // vC=-1701 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111000; // iC=-1096 
// vC = 14'b1111100111001110; // vC=-1586 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111100; // iC=-1156 
// vC = 14'b1111100010111010; // vC=-1862 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111010; // iC= -966 
// vC = 14'b1111100110011101; // vC=-1635 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000000; // iC=-1024 
// vC = 14'b1111100110001011; // vC=-1653 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010011; // iC=-1197 
// vC = 14'b1111100111000110; // vC=-1594 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110111; // iC= -969 
// vC = 14'b1111100011001110; // vC=-1842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111011; // iC=-1221 
// vC = 14'b1111100010110001; // vC=-1871 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000001; // iC=-1087 
// vC = 14'b1111100111001001; // vC=-1591 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110111; // iC=-1097 
// vC = 14'b1111100011010000; // vC=-1840 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101001; // iC=-1047 
// vC = 14'b1111100110011101; // vC=-1635 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001111; // iC=-1073 
// vC = 14'b1111100011110001; // vC=-1807 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110010; // iC=-1038 
// vC = 14'b1111100011111110; // vC=-1794 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010001; // iC=-1007 
// vC = 14'b1111100100101110; // vC=-1746 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101001; // iC= -919 
// vC = 14'b1111100101000000; // vC=-1728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010101; // iC=-1195 
// vC = 14'b1111100101010010; // vC=-1710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001001; // iC= -951 
// vC = 14'b1111100101111011; // vC=-1669 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001100; // iC=-1076 
// vC = 14'b1111100101100010; // vC=-1694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011010; // iC= -934 
// vC = 14'b1111100011011010; // vC=-1830 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000001; // iC= -895 
// vC = 14'b1111100100000000; // vC=-1792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011011; // iC= -869 
// vC = 14'b1111100010011100; // vC=-1892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000100; // iC=-1020 
// vC = 14'b1111100101000100; // vC=-1724 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110000; // iC= -976 
// vC = 14'b1111100011110000; // vC=-1808 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011100; // iC=-1060 
// vC = 14'b1111100100110010; // vC=-1742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010111; // iC=-1001 
// vC = 14'b1111100010101010; // vC=-1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011000; // iC=-1000 
// vC = 14'b1111100100011110; // vC=-1762 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101001; // iC= -855 
// vC = 14'b1111100010011100; // vC=-1892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011011; // iC= -933 
// vC = 14'b1111100101110100; // vC=-1676 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111000; // iC= -904 
// vC = 14'b1111100011010100; // vC=-1836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101110; // iC= -786 
// vC = 14'b1111100001100100; // vC=-1948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110001; // iC= -975 
// vC = 14'b1111100000111011; // vC=-1989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000010; // iC= -894 
// vC = 14'b1111100101101001; // vC=-1687 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100101; // iC=-1051 
// vC = 14'b1111100101010010; // vC=-1710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000100; // iC= -828 
// vC = 14'b1111100011101000; // vC=-1816 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010111; // iC=-1001 
// vC = 14'b1111100000110010; // vC=-1998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011000; // iC= -808 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101100; // iC= -916 
// vC = 14'b1111100010011101; // vC=-1891 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110011; // iC= -845 
// vC = 14'b1111100010000001; // vC=-1919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111010; // iC= -838 
// vC = 14'b1111100101100001; // vC=-1695 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110101; // iC=-1035 
// vC = 14'b1111100100101110; // vC=-1746 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000111; // iC= -889 
// vC = 14'b1111100101010000; // vC=-1712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111100; // iC= -836 
// vC = 14'b1111100100110101; // vC=-1739 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101011; // iC= -725 
// vC = 14'b1111100010000100; // vC=-1916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100001; // iC= -863 
// vC = 14'b1111100010100000; // vC=-1888 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000000; // iC= -768 
// vC = 14'b1111100000111100; // vC=-1988 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001000; // iC= -696 
// vC = 14'b1111100100101010; // vC=-1750 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b1111100011011010; // vC=-1830 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101010; // iC= -790 
// vC = 14'b1111100000111111; // vC=-1985 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101000; // iC= -984 
// vC = 14'b1111100001101100; // vC=-1940 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101101; // iC= -979 
// vC = 14'b1111100100101110; // vC=-1746 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000110; // iC= -954 
// vC = 14'b1111100001110111; // vC=-1929 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111010; // iC= -646 
// vC = 14'b1111100000110101; // vC=-1995 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101001; // iC= -855 
// vC = 14'b1111100001010000; // vC=-1968 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011011; // iC= -741 
// vC = 14'b1111100000001110; // vC=-2034 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011101; // iC= -675 
// vC = 14'b1111100011001110; // vC=-1842 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111000; // iC= -648 
// vC = 14'b1111100100100111; // vC=-1753 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110110; // iC= -906 
// vC = 14'b1111100001011110; // vC=-1954 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101111; // iC= -785 
// vC = 14'b1111100100010011; // vC=-1773 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100101; // iC= -731 
// vC = 14'b1111100011000110; // vC=-1850 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010101; // iC= -619 
// vC = 14'b1111100011100001; // vC=-1823 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111000; // iC= -712 
// vC = 14'b1111100001110111; // vC=-1929 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101111; // iC= -785 
// vC = 14'b1111100011100011; // vC=-1821 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100010; // iC= -606 
// vC = 14'b1111100100000000; // vC=-1792 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110000; // iC= -656 
// vC = 14'b1111100010000101; // vC=-1915 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001101; // iC= -691 
// vC = 14'b1111100010010111; // vC=-1897 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111011; // iC= -581 
// vC = 14'b1111100001100010; // vC=-1950 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000101; // iC= -763 
// vC = 14'b1111100001101000; // vC=-1944 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111001; // iC= -711 
// vC = 14'b1111100010111010; // vC=-1862 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101110; // iC= -594 
// vC = 14'b1111100000111001; // vC=-1991 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111010; // iC= -582 
// vC = 14'b1111100000100000; // vC=-2016 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111001; // iC= -519 
// vC = 14'b1111100001101111; // vC=-1937 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101101; // iC= -659 
// vC = 14'b1111011111100100; // vC=-2076 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100000; // iC= -608 
// vC = 14'b1111011111000101; // vC=-2107 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101010; // iC= -662 
// vC = 14'b1111100010100001; // vC=-1887 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001011; // iC= -693 
// vC = 14'b1111100000011110; // vC=-2018 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001011; // iC= -693 
// vC = 14'b1111011110111011; // vC=-2117 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000100; // iC= -444 
// vC = 14'b1111100011101000; // vC=-1816 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100100; // iC= -668 
// vC = 14'b1111011111010010; // vC=-2094 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010101; // iC= -491 
// vC = 14'b1111100001101001; // vC=-1943 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010000; // iC= -496 
// vC = 14'b1111011111110010; // vC=-2062 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111110011; // iC= -525 
// vC = 14'b1111011111111000; // vC=-2056 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111101; // iC= -515 
// vC = 14'b1111100001000101; // vC=-1979 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101111; // iC= -401 
// vC = 14'b1111011110111011; // vC=-2117 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101100; // iC= -532 
// vC = 14'b1111011111111011; // vC=-2053 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101101; // iC= -595 
// vC = 14'b1111100010001110; // vC=-1906 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100010; // iC= -350 
// vC = 14'b1111100000010000; // vC=-2032 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000101; // iC= -379 
// vC = 14'b1111100000011101; // vC=-2019 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110010; // iC= -590 
// vC = 14'b1111100011010101; // vC=-1835 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111110; // iC= -450 
// vC = 14'b1111100010010000; // vC=-1904 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111100; // iC= -324 
// vC = 14'b1111100010011110; // vC=-1890 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010011; // iC= -493 
// vC = 14'b1111011111010100; // vC=-2092 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001101; // iC= -307 
// vC = 14'b1111011111111011; // vC=-2053 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001010; // iC= -374 
// vC = 14'b1111011111010111; // vC=-2089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011110; // iC= -354 
// vC = 14'b1111011111011101; // vC=-2083 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111000; // iC= -456 
// vC = 14'b1111011110110101; // vC=-2123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010000; // iC= -240 
// vC = 14'b1111011110111000; // vC=-2120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110110; // iC= -394 
// vC = 14'b1111100010100010; // vC=-1886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000011; // iC= -189 
// vC = 14'b1111100011000101; // vC=-1851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010111; // iC= -233 
// vC = 14'b1111100001001111; // vC=-1969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001110; // iC= -114 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110101; // iC= -203 
// vC = 14'b1111011111010110; // vC=-2090 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110100; // iC= -396 
// vC = 14'b1111100010001110; // vC=-1906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001101; // iC= -243 
// vC = 14'b1111100001011000; // vC=-1960 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101111; // iC= -209 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000100; // iC= -188 
// vC = 14'b1111011111000001; // vC=-2111 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100100; // iC=  -92 
// vC = 14'b1111100010111110; // vC=-1858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110101010; // iC=  -86 
// vC = 14'b1111100011001001; // vC=-1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111011000; // iC=  -40 
// vC = 14'b1111100000110101; // vC=-1995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000001; // iC= -255 
// vC = 14'b1111100000010010; // vC=-2030 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001000; // iC=  -56 
// vC = 14'b1111011111001000; // vC=-2104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111110111; // iC=   -9 
// vC = 14'b1111011111100000; // vC=-2080 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001100; // iC=   12 
// vC = 14'b1111011111100011; // vC=-2077 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111101; // iC=  -67 
// vC = 14'b1111100001001110; // vC=-1970 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001011; // iC=   75 
// vC = 14'b1111100000101010; // vC=-2006 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000110; // iC= -122 
// vC = 14'b1111100000100101; // vC=-2011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110101111; // iC=  -81 
// vC = 14'b1111011110001111; // vC=-2161 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111001; // iC=   -7 
// vC = 14'b1111100000011110; // vC=-2018 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010011; // iC=  -45 
// vC = 14'b1111100000000111; // vC=-2041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111000; // iC=  120 
// vC = 14'b1111100000111101; // vC=-1987 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111000; // iC=  184 
// vC = 14'b1111100001101111; // vC=-1937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101001; // iC=   41 
// vC = 14'b1111011111101010; // vC=-2070 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011010; // iC=  154 
// vC = 14'b1111100000100010; // vC=-2014 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010100; // iC=   84 
// vC = 14'b1111011110110101; // vC=-2123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110110; // iC=  310 
// vC = 14'b1111100010110100; // vC=-1868 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001010; // iC=  202 
// vC = 14'b1111100001101110; // vC=-1938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001010; // iC=  394 
// vC = 14'b1111011111110010; // vC=-2062 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110110; // iC=  118 
// vC = 14'b1111100000011111; // vC=-2017 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110111; // iC=  375 
// vC = 14'b1111011110111100; // vC=-2116 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010110; // iC=  150 
// vC = 14'b1111100010100001; // vC=-1887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011110; // iC=  350 
// vC = 14'b1111100000000100; // vC=-2044 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110000; // iC=  240 
// vC = 14'b1111100010101111; // vC=-1873 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100001; // iC=  289 
// vC = 14'b1111011111011111; // vC=-2081 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001001; // iC=  265 
// vC = 14'b1111100011000101; // vC=-1851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101001; // iC=  425 
// vC = 14'b1111100011001011; // vC=-1845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100101; // iC=  485 
// vC = 14'b1111100011011110; // vC=-1826 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000010; // iC=  450 
// vC = 14'b1111011111110000; // vC=-2064 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010101; // iC=  405 
// vC = 14'b1111100011011110; // vC=-1826 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100011; // iC=  611 
// vC = 14'b1111100000111001; // vC=-1991 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100001; // iC=  545 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100110; // iC=  486 
// vC = 14'b1111011110111001; // vC=-2119 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111011; // iC=  699 
// vC = 14'b1111100000100100; // vC=-2012 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000111; // iC=  455 
// vC = 14'b1111100001110110; // vC=-1930 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101110; // iC=  686 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001010; // iC=  778 
// vC = 14'b1111100001011100; // vC=-1956 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011101; // iC=  733 
// vC = 14'b1111100000101100; // vC=-2004 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110001; // iC=  753 
// vC = 14'b1111100011110000; // vC=-1808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111100; // iC=  636 
// vC = 14'b1111100001111100; // vC=-1924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001010; // iC=  714 
// vC = 14'b1111100011011111; // vC=-1825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000101; // iC=  709 
// vC = 14'b1111100010001110; // vC=-1906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001010; // iC=  778 
// vC = 14'b1111100001011110; // vC=-1954 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000101; // iC=  773 
// vC = 14'b1111011111101010; // vC=-2070 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100101; // iC=  677 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111111; // iC= 1023 
// vC = 14'b1111100000111010; // vC=-1990 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011101; // iC=  797 
// vC = 14'b1111100011001010; // vC=-1846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000001; // iC= 1025 
// vC = 14'b1111011111111100; // vC=-2052 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000101; // iC=  837 
// vC = 14'b1111100001000010; // vC=-1982 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101101; // iC=  813 
// vC = 14'b1111100100001101; // vC=-1779 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011010; // iC=  922 
// vC = 14'b1111100011000110; // vC=-1850 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100101; // iC= 1061 
// vC = 14'b1111100000011010; // vC=-2022 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010001; // iC=  913 
// vC = 14'b1111100100010110; // vC=-1770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000110; // iC= 1158 
// vC = 14'b1111100011010011; // vC=-1837 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111110; // iC= 1022 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010010; // iC= 1170 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111010; // iC= 1018 
// vC = 14'b1111100001110000; // vC=-1936 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111111; // iC= 1087 
// vC = 14'b1111100011110101; // vC=-1803 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010000; // iC= 1168 
// vC = 14'b1111100010000010; // vC=-1918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001101; // iC= 1101 
// vC = 14'b1111100001000010; // vC=-1982 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001001; // iC= 1033 
// vC = 14'b1111100001111011; // vC=-1925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111000; // iC= 1272 
// vC = 14'b1111100011100110; // vC=-1818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010110; // iC= 1238 
// vC = 14'b1111100010111110; // vC=-1858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010011; // iC= 1363 
// vC = 14'b1111100011011011; // vC=-1829 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000010; // iC= 1282 
// vC = 14'b1111100100110100; // vC=-1740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001010; // iC= 1290 
// vC = 14'b1111100101010011; // vC=-1709 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101011; // iC= 1195 
// vC = 14'b1111100100000110; // vC=-1786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000010; // iC= 1346 
// vC = 14'b1111100101000100; // vC=-1724 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111100; // iC= 1340 
// vC = 14'b1111100011001001; // vC=-1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110000; // iC= 1328 
// vC = 14'b1111100010110010; // vC=-1870 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111101; // iC= 1405 
// vC = 14'b1111100011010000; // vC=-1840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011101; // iC= 1309 
// vC = 14'b1111100110011000; // vC=-1640 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100111; // iC= 1383 
// vC = 14'b1111100011010010; // vC=-1838 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001011; // iC= 1355 
// vC = 14'b1111100110010000; // vC=-1648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011001; // iC= 1497 
// vC = 14'b1111100101010010; // vC=-1710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001110; // iC= 1550 
// vC = 14'b1111100101101000; // vC=-1688 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001100; // iC= 1484 
// vC = 14'b1111100110000101; // vC=-1659 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110111; // iC= 1527 
// vC = 14'b1111100010111101; // vC=-1859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110101; // iC= 1653 
// vC = 14'b1111100011100011; // vC=-1821 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110011; // iC= 1459 
// vC = 14'b1111100011100111; // vC=-1817 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100001; // iC= 1633 
// vC = 14'b1111100011000101; // vC=-1851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100100; // iC= 1444 
// vC = 14'b1111100111000101; // vC=-1595 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000010; // iC= 1602 
// vC = 14'b1111100110101111; // vC=-1617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011001; // iC= 1625 
// vC = 14'b1111100101010011; // vC=-1709 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010010; // iC= 1682 
// vC = 14'b1111100101100110; // vC=-1690 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001000; // iC= 1608 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010001; // iC= 1745 
// vC = 14'b1111100011001001; // vC=-1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100110; // iC= 1638 
// vC = 14'b1111100110001111; // vC=-1649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001010; // iC= 1482 
// vC = 14'b1111100011110000; // vC=-1808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110100; // iC= 1652 
// vC = 14'b1111100111010111; // vC=-1577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100100; // iC= 1764 
// vC = 14'b1111100101011111; // vC=-1697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000000; // iC= 1728 
// vC = 14'b1111100101000100; // vC=-1724 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100111; // iC= 1639 
// vC = 14'b1111101000110000; // vC=-1488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111100; // iC= 1788 
// vC = 14'b1111100100111011; // vC=-1733 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011011; // iC= 1755 
// vC = 14'b1111101000010000; // vC=-1520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001001; // iC= 1673 
// vC = 14'b1111100101011001; // vC=-1703 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b1111100100100101; // vC=-1755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011111; // iC= 1759 
// vC = 14'b1111100111111110; // vC=-1538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000111; // iC= 1735 
// vC = 14'b1111101001000100; // vC=-1468 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b1111100100111010; // vC=-1734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010100; // iC= 1684 
// vC = 14'b1111100110001101; // vC=-1651 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101111; // iC= 1711 
// vC = 14'b1111100110110001; // vC=-1615 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010101; // iC= 1877 
// vC = 14'b1111100111101010; // vC=-1558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001001; // iC= 1737 
// vC = 14'b1111100101011001; // vC=-1703 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100001; // iC= 1761 
// vC = 14'b1111101000011100; // vC=-1508 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111100111101100; // vC=-1556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011010; // iC= 1882 
// vC = 14'b1111100110000100; // vC=-1660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b1111100110010000; // vC=-1648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100010; // iC= 1954 
// vC = 14'b1111101000000100; // vC=-1532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010011; // iC= 1811 
// vC = 14'b1111101001011100; // vC=-1444 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001000; // iC= 1928 
// vC = 14'b1111100110101110; // vC=-1618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b1111101010110101; // vC=-1355 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001000; // iC= 1736 
// vC = 14'b1111101001111001; // vC=-1415 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b1111100111000111; // vC=-1593 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110010; // iC= 1906 
// vC = 14'b1111101000000011; // vC=-1533 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010011; // iC= 1875 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110101; // iC= 2037 
// vC = 14'b1111100111110110; // vC=-1546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111101001111011; // vC=-1413 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111101000001111; // vC=-1521 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011101; // iC= 1821 
// vC = 14'b1111101010111111; // vC=-1345 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010100; // iC= 1876 
// vC = 14'b1111101000001000; // vC=-1528 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b1111101001101011; // vC=-1429 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111101010011111; // vC=-1377 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001001; // iC= 2121 
// vC = 14'b1111101010011110; // vC=-1378 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100101; // iC= 1957 
// vC = 14'b1111101000000011; // vC=-1533 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111101010000011; // vC=-1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101110; // iC= 1902 
// vC = 14'b1111101011101100; // vC=-1300 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b1111101010010001; // vC=-1391 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110100; // iC= 1844 
// vC = 14'b1111101011011010; // vC=-1318 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b1111101001111000; // vC=-1416 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b1111101100110010; // vC=-1230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110001; // iC= 1841 
// vC = 14'b1111101010010110; // vC=-1386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011000; // iC= 2136 
// vC = 14'b1111101100011110; // vC=-1250 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111101011111001; // vC=-1287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b1111101011111100; // vC=-1284 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b1111101011000011; // vC=-1341 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110000; // iC= 1968 
// vC = 14'b1111101010111100; // vC=-1348 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b1111101010011101; // vC=-1379 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b1111101100101111; // vC=-1233 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111110; // iC= 2046 
// vC = 14'b1111101011100100; // vC=-1308 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111101010011011; // vC=-1381 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b1111101110011010; // vC=-1126 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111101010101001; // vC=-1367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001001; // iC= 2185 
// vC = 14'b1111101100111000; // vC=-1224 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010010; // iC= 2002 
// vC = 14'b1111101011110001; // vC=-1295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100010; // iC= 2146 
// vC = 14'b1111110000000010; // vC=-1022 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111101110001001; // vC=-1143 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001011; // iC= 2123 
// vC = 14'b1111101111100010; // vC=-1054 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b1111101101111100; // vC=-1156 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b1111101101101111; // vC=-1169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100010; // iC= 1954 
// vC = 14'b1111101111110010; // vC=-1038 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011011; // iC= 2203 
// vC = 14'b1111110000001011; // vC=-1013 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011011; // iC= 2203 
// vC = 14'b1111101101110110; // vC=-1162 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b1111101100100111; // vC=-1241 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001101; // iC= 2189 
// vC = 14'b1111110000111100; // vC= -964 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011000; // iC= 2072 
// vC = 14'b1111101111011111; // vC=-1057 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001110; // iC= 1934 
// vC = 14'b1111101101011100; // vC=-1188 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110110; // iC= 2166 
// vC = 14'b1111101111111001; // vC=-1031 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000011; // iC= 2179 
// vC = 14'b1111101111100010; // vC=-1054 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101100; // iC= 2220 
// vC = 14'b1111101111001101; // vC=-1075 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100000; // iC= 2208 
// vC = 14'b1111110001011011; // vC= -933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100011; // iC= 2083 
// vC = 14'b1111101111110100; // vC=-1036 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011101; // iC= 2205 
// vC = 14'b1111110010001001; // vC= -887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111110000101011; // vC= -981 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111110000100001; // vC= -991 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b1111101111000101; // vC=-1083 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111110000101101; // vC= -979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101110; // iC= 2222 
// vC = 14'b1111101111000010; // vC=-1086 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111110011001110; // vC= -818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101110; // iC= 2222 
// vC = 14'b1111110001100100; // vC= -924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111110001010110; // vC= -938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110111; // iC= 1911 
// vC = 14'b1111101111110111; // vC=-1033 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100000; // iC= 2144 
// vC = 14'b1111101111000100; // vC=-1084 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110000; // iC= 2096 
// vC = 14'b1111110001000011; // vC= -957 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b1111110011011001; // vC= -807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110101; // iC= 2101 
// vC = 14'b1111110011101000; // vC= -792 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100111; // iC= 2087 
// vC = 14'b1111110011010000; // vC= -816 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011111; // iC= 2015 
// vC = 14'b1111110010110001; // vC= -847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000000; // iC= 2240 
// vC = 14'b1111110000110001; // vC= -975 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b1111110011010010; // vC= -814 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001001; // iC= 1993 
// vC = 14'b1111110011001011; // vC= -821 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b1111110101010000; // vC= -688 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100110; // iC= 2214 
// vC = 14'b1111110000100100; // vC= -988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b1111110000110011; // vC= -973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111010; // iC= 2106 
// vC = 14'b1111110011001111; // vC= -817 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110110; // iC= 1974 
// vC = 14'b1111110011001110; // vC= -818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111110011110101; // vC= -779 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001000; // iC= 2184 
// vC = 14'b1111110001110110; // vC= -906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000101; // iC= 2053 
// vC = 14'b1111110010010100; // vC= -876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b1111110101110000; // vC= -656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110000; // iC= 2096 
// vC = 14'b1111110010100111; // vC= -857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101011; // iC= 2219 
// vC = 14'b1111110110011110; // vC= -610 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111110010110110; // vC= -842 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111110010011101; // vC= -867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110010; // iC= 2226 
// vC = 14'b1111110100101000; // vC= -728 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010000; // iC= 2064 
// vC = 14'b1111110101111101; // vC= -643 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110001; // iC= 1969 
// vC = 14'b1111110111001001; // vC= -567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110110; // iC= 2230 
// vC = 14'b1111110100001111; // vC= -753 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111110011000101; // vC= -827 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010100; // iC= 2260 
// vC = 14'b1111110011101010; // vC= -790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111110101101010; // vC= -662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010011; // iC= 2131 
// vC = 14'b1111110111010100; // vC= -556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001111; // iC= 2127 
// vC = 14'b1111110011010110; // vC= -810 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111110100001100; // vC= -756 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001111; // iC= 2191 
// vC = 14'b1111110110010010; // vC= -622 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b1111110101110111; // vC= -649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010011; // iC= 2067 
// vC = 14'b1111110111101000; // vC= -536 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111110101101011; // vC= -661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b1111110101011111; // vC= -673 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110110; // iC= 2102 
// vC = 14'b1111110100111101; // vC= -707 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b1111111000011000; // vC= -488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111110101010000; // vC= -688 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111111000010000; // vC= -496 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b1111111000101010; // vC= -470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111011; // iC= 2171 
// vC = 14'b1111110110000111; // vC= -633 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011000; // iC= 2200 
// vC = 14'b1111110111101101; // vC= -531 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011110; // iC= 2142 
// vC = 14'b1111111001101110; // vC= -402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100110; // iC= 2022 
// vC = 14'b1111111000111000; // vC= -456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000011; // iC= 2179 
// vC = 14'b1111111000011000; // vC= -488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111010; // iC= 2106 
// vC = 14'b1111111001111100; // vC= -388 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011110; // iC= 2014 
// vC = 14'b1111110111111001; // vC= -519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001000; // iC= 2120 
// vC = 14'b1111110110000110; // vC= -634 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000110; // iC= 2182 
// vC = 14'b1111111000111100; // vC= -452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010000; // iC= 2256 
// vC = 14'b1111110111000001; // vC= -575 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b1111110111111001; // vC= -519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100101; // iC= 2149 
// vC = 14'b1111111001111110; // vC= -386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b1111110111100000; // vC= -544 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111111000010001; // vC= -495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b1111110111111110; // vC= -514 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111100; // iC= 2108 
// vC = 14'b1111111000101101; // vC= -467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010000; // iC= 2064 
// vC = 14'b1111111010111000; // vC= -328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000101; // iC= 2245 
// vC = 14'b1111111001011001; // vC= -423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001110; // iC= 2254 
// vC = 14'b1111111011111111; // vC= -257 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010111; // iC= 2263 
// vC = 14'b1111111010101111; // vC= -337 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101101; // iC= 2029 
// vC = 14'b1111111000111110; // vC= -450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111100; // iC= 1980 
// vC = 14'b1111111100100100; // vC= -220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000011; // iC= 2051 
// vC = 14'b1111111000111000; // vC= -456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110011; // iC= 2227 
// vC = 14'b1111111011111110; // vC= -258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b1111111010111011; // vC= -325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100100; // iC= 2148 
// vC = 14'b1111111010101010; // vC= -342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110011; // iC= 2163 
// vC = 14'b1111111001010001; // vC= -431 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b1111111100110110; // vC= -202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111111100010010; // vC= -238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100000; // iC= 2016 
// vC = 14'b1111111001111000; // vC= -392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111111; // iC= 2111 
// vC = 14'b1111111101110111; // vC= -137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011110; // iC= 2014 
// vC = 14'b1111111100100011; // vC= -221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011010; // iC= 2074 
// vC = 14'b1111111010011001; // vC= -359 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101101; // iC= 2157 
// vC = 14'b1111111100001100; // vC= -244 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111111110010101; // vC= -107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b1111111010001000; // vC= -376 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111111011100000; // vC= -288 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b1111111110100011; // vC=  -93 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000100; // iC= 2244 
// vC = 14'b1111111111011010; // vC=  -38 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b1111111100010101; // vC= -235 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110000; // iC= 2032 
// vC = 14'b1111111110100100; // vC=  -92 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000010; // iC= 2050 
// vC = 14'b1111111110010100; // vC= -108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111111100111001; // vC= -199 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b1111111011100100; // vC= -284 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011010; // iC= 2138 
// vC = 14'b1111111110100010; // vC=  -94 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111111111011101; // vC=  -35 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b1111111100001111; // vC= -241 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011001; // iC= 2201 
// vC = 14'b1111111111010100; // vC=  -44 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010001; // iC= 2065 
// vC = 14'b1111111101111011; // vC= -133 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011100; // iC= 2204 
// vC = 14'b1111111110110011; // vC=  -77 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101100; // iC= 2156 
// vC = 14'b0000000000010011; // vC=   19 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111111110011111; // vC=  -97 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111111101110001; // vC= -143 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011111; // iC= 2143 
// vC = 14'b0000000000101110; // vC=   46 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101000; // iC= 2216 
// vC = 14'b1111111110001001; // vC= -119 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110001; // iC= 2033 
// vC = 14'b0000000001100101; // vC=  101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000010; // iC= 2050 
// vC = 14'b1111111111011010; // vC=  -38 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010011; // iC= 2067 
// vC = 14'b0000000000011100; // vC=   28 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100001; // iC= 2209 
// vC = 14'b0000000001000010; // vC=   66 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100101; // iC= 2149 
// vC = 14'b0000000000101000; // vC=   40 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b0000000001010000; // vC=   80 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111111111101111; // vC=  -17 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010010; // iC= 2194 
// vC = 14'b0000000010110010; // vC=  178 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000010; // iC= 1922 
// vC = 14'b1111111110011010; // vC= -102 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111111111111111; // vC=   -1 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000101; // iC= 1925 
// vC = 14'b0000000010111101; // vC=  189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b0000000010110011; // vC=  179 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111000; // iC= 2168 
// vC = 14'b0000000010000111; // vC=  135 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b0000000010011101; // vC=  157 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b0000000010101010; // vC=  170 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110001; // iC= 2161 
// vC = 14'b0000000001110011; // vC=  115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101101; // iC= 2029 
// vC = 14'b0000000000000101; // vC=    5 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101000; // iC= 2024 
// vC = 14'b0000000011110100; // vC=  244 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b0000000010001100; // vC=  140 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011111; // iC= 2207 
// vC = 14'b0000000000001010; // vC=   10 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000110; // iC= 2118 
// vC = 14'b0000000100011001; // vC=  281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b0000000010110101; // vC=  181 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001000; // iC= 1992 
// vC = 14'b0000000010010110; // vC=  150 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b0000000001010100; // vC=   84 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111110; // iC= 2046 
// vC = 14'b0000000000001101; // vC=   13 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b0000000010001101; // vC=  141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b0000000100011101; // vC=  285 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b0000000100000111; // vC=  263 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b0000000101100110; // vC=  358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001011; // iC= 2187 
// vC = 14'b0000000101001110; // vC=  334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001011; // iC= 2123 
// vC = 14'b0000000011011100; // vC=  220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b0000000001001100; // vC=   76 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b0000000101101010; // vC=  362 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110000; // iC= 1904 
// vC = 14'b0000000010011110; // vC=  158 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b0000000101011000; // vC=  344 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110001; // iC= 1969 
// vC = 14'b0000000001110101; // vC=  117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000000; // iC= 1856 
// vC = 14'b0000000110100101; // vC=  421 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b0000000011101111; // vC=  239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110110; // iC= 2166 
// vC = 14'b0000000100111110; // vC=  318 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111100; // iC= 2108 
// vC = 14'b0000000010100111; // vC=  167 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b0000000110101111; // vC=  431 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100001; // iC= 2017 
// vC = 14'b0000000110000000; // vC=  384 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001101; // iC= 2125 
// vC = 14'b0000000011010100; // vC=  212 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b0000000100001101; // vC=  269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011011; // iC= 2075 
// vC = 14'b0000000100010011; // vC=  275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b0000000011111000; // vC=  248 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b0000000100111000; // vC=  312 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001010; // iC= 1866 
// vC = 14'b0000000101011000; // vC=  344 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b0000000111101001; // vC=  489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101000; // iC= 1832 
// vC = 14'b0000000101111010; // vC=  378 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b0000000111000011; // vC=  451 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b0000000111000101; // vC=  453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000000101101101; // vC=  365 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011000; // iC= 1816 
// vC = 14'b0000000100001100; // vC=  268 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b0000000100110100; // vC=  308 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b0000000100111101; // vC=  317 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b0000000111010001; // vC=  465 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000000; // iC= 1920 
// vC = 14'b0000001000001001; // vC=  521 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001001; // iC= 1865 
// vC = 14'b0000001000111101; // vC=  573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b0000000110101011; // vC=  427 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b0000000111010101; // vC=  469 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011100; // iC= 1884 
// vC = 14'b0000000110111101; // vC=  445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100000; // iC= 2080 
// vC = 14'b0000000110101110; // vC=  430 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b0000000101011011; // vC=  347 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b0000000111111011; // vC=  507 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b0000000111011100; // vC=  476 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011110; // iC= 2078 
// vC = 14'b0000000111010101; // vC=  469 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000001001100010; // vC=  610 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b0000001000110100; // vC=  564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110001; // iC= 1777 
// vC = 14'b0000000110000110; // vC=  390 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110010; // iC= 1906 
// vC = 14'b0000001010110111; // vC=  695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b0000001010010010; // vC=  658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001001; // iC= 2057 
// vC = 14'b0000001000110010; // vC=  562 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000001; // iC= 1793 
// vC = 14'b0000001001111011; // vC=  635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b0000001001011101; // vC=  605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000101; // iC= 2053 
// vC = 14'b0000001011110000; // vC=  752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110111; // iC= 2039 
// vC = 14'b0000001001011110; // vC=  606 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b0000001011010100; // vC=  724 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000000; // iC= 1920 
// vC = 14'b0000001001011001; // vC=  601 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010001; // iC= 1937 
// vC = 14'b0000001001011100; // vC=  604 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b0000001001011111; // vC=  607 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101010; // iC= 1834 
// vC = 14'b0000001011100001; // vC=  737 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b0000001011110010; // vC=  754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100111; // iC= 1831 
// vC = 14'b0000001000000110; // vC=  518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110100; // iC= 2036 
// vC = 14'b0000001100101100; // vC=  812 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b0000001100010010; // vC=  786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b0000001011111011; // vC=  763 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000001010110110; // vC=  694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b0000001100101001; // vC=  809 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b0000001001111011; // vC=  635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010111; // iC= 1751 
// vC = 14'b0000001000111100; // vC=  572 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b0000001011111000; // vC=  760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011011; // iC= 1755 
// vC = 14'b0000001011110101; // vC=  757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110010; // iC= 1842 
// vC = 14'b0000001001001100; // vC=  588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001110; // iC= 1870 
// vC = 14'b0000001101010101; // vC=  853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110000; // iC= 1840 
// vC = 14'b0000001101110101; // vC=  885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b0000001101101011; // vC=  875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000000; // iC= 1984 
// vC = 14'b0000001011101110; // vC=  750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101110; // iC= 1838 
// vC = 14'b0000001100011111; // vC=  799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001010; // iC= 1674 
// vC = 14'b0000001101001101; // vC=  845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011111; // iC= 1695 
// vC = 14'b0000001101100111; // vC=  871 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000000; // iC= 1728 
// vC = 14'b0000001100010100; // vC=  788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b0000001110000010; // vC=  898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000100; // iC= 1796 
// vC = 14'b0000001111000111; // vC=  967 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111000; // iC= 1784 
// vC = 14'b0000001111011100; // vC=  988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000011; // iC= 1667 
// vC = 14'b0000001101100110; // vC=  870 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111000; // iC= 1848 
// vC = 14'b0000001011100000; // vC=  736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b0000001101110100; // vC=  884 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100101; // iC= 1765 
// vC = 14'b0000001011011011; // vC=  731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b0000001111011010; // vC=  986 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b0000010000000011; // vC= 1027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100111; // iC= 1895 
// vC = 14'b0000001101111111; // vC=  895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011011; // iC= 1755 
// vC = 14'b0000001110010000; // vC=  912 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100111; // iC= 1703 
// vC = 14'b0000001100101110; // vC=  814 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b0000001101010011; // vC=  851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100001; // iC= 1825 
// vC = 14'b0000001110111100; // vC=  956 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110101; // iC= 1717 
// vC = 14'b0000001011110001; // vC=  753 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b0000001110010110; // vC=  918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111011; // iC= 1723 
// vC = 14'b0000010000000110; // vC= 1030 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101000; // iC= 1640 
// vC = 14'b0000010000110001; // vC= 1073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110011; // iC= 1907 
// vC = 14'b0000010000110011; // vC= 1075 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000110; // iC= 1862 
// vC = 14'b0000001101000110; // vC=  838 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000011; // iC= 1731 
// vC = 14'b0000001101001111; // vC=  847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001110; // iC= 1614 
// vC = 14'b0000001111011001; // vC=  985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010111; // iC= 1815 
// vC = 14'b0000010000101010; // vC= 1066 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101101; // iC= 1645 
// vC = 14'b0000010001010111; // vC= 1111 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000000; // iC= 1728 
// vC = 14'b0000001111000010; // vC=  962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011100; // iC= 1692 
// vC = 14'b0000001111100111; // vC=  999 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011100; // iC= 1692 
// vC = 14'b0000001101100101; // vC=  869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111001; // iC= 1657 
// vC = 14'b0000010001011011; // vC= 1115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010110; // iC= 1558 
// vC = 14'b0000010000000001; // vC= 1025 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010110; // iC= 1750 
// vC = 14'b0000010000011111; // vC= 1055 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100111; // iC= 1575 
// vC = 14'b0000010001011101; // vC= 1117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001111; // iC= 1871 
// vC = 14'b0000001111101100; // vC= 1004 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011011; // iC= 1691 
// vC = 14'b0000010010100000; // vC= 1184 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010011; // iC= 1683 
// vC = 14'b0000001111110110; // vC= 1014 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010000; // iC= 1744 
// vC = 14'b0000010011000101; // vC= 1221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001001; // iC= 1609 
// vC = 14'b0000010000111000; // vC= 1080 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011110; // iC= 1758 
// vC = 14'b0000010011010001; // vC= 1233 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110110; // iC= 1654 
// vC = 14'b0000001110100011; // vC=  931 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010110; // iC= 1686 
// vC = 14'b0000010010111011; // vC= 1211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000101; // iC= 1605 
// vC = 14'b0000010001011111; // vC= 1119 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111011; // iC= 1595 
// vC = 14'b0000010001100100; // vC= 1124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010110; // iC= 1814 
// vC = 14'b0000010010010010; // vC= 1170 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010011; // iC= 1619 
// vC = 14'b0000010000010111; // vC= 1047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011011; // iC= 1819 
// vC = 14'b0000010001110000; // vC= 1136 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011000; // iC= 1752 
// vC = 14'b0000001111010001; // vC=  977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b0000010011100110; // vC= 1254 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001110; // iC= 1550 
// vC = 14'b0000010100000100; // vC= 1284 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000110; // iC= 1670 
// vC = 14'b0000010001010001; // vC= 1105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101001; // iC= 1577 
// vC = 14'b0000010011101000; // vC= 1256 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111100; // iC= 1724 
// vC = 14'b0000010100000110; // vC= 1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101101; // iC= 1645 
// vC = 14'b0000010011011001; // vC= 1241 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111001; // iC= 1721 
// vC = 14'b0000010010100011; // vC= 1187 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101101; // iC= 1709 
// vC = 14'b0000010000000111; // vC= 1031 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101110; // iC= 1774 
// vC = 14'b0000010011100110; // vC= 1254 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010100; // iC= 1556 
// vC = 14'b0000010010100100; // vC= 1188 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111000; // iC= 1656 
// vC = 14'b0000010010110010; // vC= 1202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110011; // iC= 1587 
// vC = 14'b0000010001000000; // vC= 1088 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110111; // iC= 1527 
// vC = 14'b0000010010111001; // vC= 1209 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010111; // iC= 1687 
// vC = 14'b0000010000111001; // vC= 1081 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100011; // iC= 1699 
// vC = 14'b0000010000110110; // vC= 1078 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011101; // iC= 1629 
// vC = 14'b0000010010111110; // vC= 1214 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000001; // iC= 1473 
// vC = 14'b0000010010101011; // vC= 1195 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111111; // iC= 1471 
// vC = 14'b0000010100010101; // vC= 1301 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101010; // iC= 1642 
// vC = 14'b0000010101110001; // vC= 1393 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011101; // iC= 1565 
// vC = 14'b0000010110000100; // vC= 1412 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110110; // iC= 1398 
// vC = 14'b0000010010010111; // vC= 1175 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110100; // iC= 1460 
// vC = 14'b0000010101111011; // vC= 1403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011010; // iC= 1562 
// vC = 14'b0000010001101101; // vC= 1133 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101010; // iC= 1642 
// vC = 14'b0000010101010110; // vC= 1366 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011100; // iC= 1436 
// vC = 14'b0000010101001110; // vC= 1358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100100; // iC= 1508 
// vC = 14'b0000010011011101; // vC= 1245 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110100; // iC= 1524 
// vC = 14'b0000010110011000; // vC= 1432 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011110; // iC= 1374 
// vC = 14'b0000010110110101; // vC= 1461 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101101; // iC= 1645 
// vC = 14'b0000010010011100; // vC= 1180 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100001; // iC= 1441 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000011; // iC= 1603 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011101; // iC= 1565 
// vC = 14'b0000010110011100; // vC= 1436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111101; // iC= 1661 
// vC = 14'b0000010011101000; // vC= 1256 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100100; // iC= 1572 
// vC = 14'b0000010110110101; // vC= 1461 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110000; // iC= 1648 
// vC = 14'b0000010110011110; // vC= 1438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010000; // iC= 1360 
// vC = 14'b0000010100000110; // vC= 1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101001; // iC= 1641 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111100; // iC= 1340 
// vC = 14'b0000010110000100; // vC= 1412 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011011; // iC= 1371 
// vC = 14'b0000010101001101; // vC= 1357 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101101; // iC= 1389 
// vC = 14'b0000010111101100; // vC= 1516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111011; // iC= 1403 
// vC = 14'b0000011000000011; // vC= 1539 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010000; // iC= 1424 
// vC = 14'b0000010100001111; // vC= 1295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111100; // iC= 1532 
// vC = 14'b0000010100000101; // vC= 1285 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111111; // iC= 1279 
// vC = 14'b0000010111111111; // vC= 1535 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100111; // iC= 1511 
// vC = 14'b0000010111001001; // vC= 1481 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000011; // iC= 1539 
// vC = 14'b0000010101110010; // vC= 1394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011010; // iC= 1370 
// vC = 14'b0000010110011000; // vC= 1432 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111110; // iC= 1406 
// vC = 14'b0000010101101010; // vC= 1386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111100; // iC= 1340 
// vC = 14'b0000010111011010; // vC= 1498 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011101; // iC= 1309 
// vC = 14'b0000010101011110; // vC= 1374 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011101; // iC= 1437 
// vC = 14'b0000011001000010; // vC= 1602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010101; // iC= 1429 
// vC = 14'b0000010111101011; // vC= 1515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101101; // iC= 1261 
// vC = 14'b0000011001010110; // vC= 1622 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010110; // iC= 1238 
// vC = 14'b0000010110101010; // vC= 1450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011110; // iC= 1246 
// vC = 14'b0000010111110010; // vC= 1522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100000; // iC= 1440 
// vC = 14'b0000010101010000; // vC= 1360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001100; // iC= 1292 
// vC = 14'b0000011001010110; // vC= 1622 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010010; // iC= 1490 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000011; // iC= 1411 
// vC = 14'b0000010110010101; // vC= 1429 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101111; // iC= 1327 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111010; // iC= 1210 
// vC = 14'b0000010110110010; // vC= 1458 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110010; // iC= 1330 
// vC = 14'b0000010101100010; // vC= 1378 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000011; // iC= 1283 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110000; // iC= 1328 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011001; // iC= 1433 
// vC = 14'b0000011000110001; // vC= 1585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011010; // iC= 1370 
// vC = 14'b0000011001011010; // vC= 1626 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011000; // iC= 1176 
// vC = 14'b0000011001011011; // vC= 1627 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010101; // iC= 1429 
// vC = 14'b0000010110100101; // vC= 1445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101000; // iC= 1448 
// vC = 14'b0000011010010001; // vC= 1681 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101100; // iC= 1260 
// vC = 14'b0000011010000100; // vC= 1668 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010111; // iC= 1175 
// vC = 14'b0000011000101100; // vC= 1580 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110010; // iC= 1330 
// vC = 14'b0000010111111001; // vC= 1529 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111111; // iC= 1215 
// vC = 14'b0000010111101011; // vC= 1515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100010; // iC= 1314 
// vC = 14'b0000011000101101; // vC= 1581 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011111; // iC= 1311 
// vC = 14'b0000011010010011; // vC= 1683 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100101; // iC= 1317 
// vC = 14'b0000011000100101; // vC= 1573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100001; // iC= 1377 
// vC = 14'b0000011010001110; // vC= 1678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000101; // iC= 1349 
// vC = 14'b0000011000110111; // vC= 1591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111010; // iC= 1338 
// vC = 14'b0000011011100000; // vC= 1760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110110; // iC= 1206 
// vC = 14'b0000010111111100; // vC= 1532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101111; // iC= 1391 
// vC = 14'b0000011000111001; // vC= 1593 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011000; // iC= 1240 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111001; // iC= 1273 
// vC = 14'b0000010111001100; // vC= 1484 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011110; // iC= 1374 
// vC = 14'b0000011001000010; // vC= 1602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100100; // iC= 1316 
// vC = 14'b0000011011010100; // vC= 1748 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001000; // iC= 1160 
// vC = 14'b0000011001111000; // vC= 1656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101100; // iC= 1260 
// vC = 14'b0000011011111101; // vC= 1789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000110; // iC= 1350 
// vC = 14'b0000011010110110; // vC= 1718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000011; // iC= 1347 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001010; // iC= 1034 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011100; // iC= 1116 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011000; // iC= 1048 
// vC = 14'b0000011010010100; // vC= 1684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101000; // iC= 1192 
// vC = 14'b0000011011011010; // vC= 1754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010111; // iC= 1047 
// vC = 14'b0000011010100000; // vC= 1696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110110; // iC= 1014 
// vC = 14'b0000011001010001; // vC= 1617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000010; // iC= 1090 
// vC = 14'b0000011010000110; // vC= 1670 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000011; // iC= 1155 
// vC = 14'b0000011001000101; // vC= 1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010110; // iC=  982 
// vC = 14'b0000011000110110; // vC= 1590 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011111; // iC=  991 
// vC = 14'b0000011100101110; // vC= 1838 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101001; // iC= 1129 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110100; // iC= 1076 
// vC = 14'b0000011001011111; // vC= 1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100100; // iC=  996 
// vC = 14'b0000011011111000; // vC= 1784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110100; // iC= 1140 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001001; // iC= 1161 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001010; // iC=  970 
// vC = 14'b0000011010101111; // vC= 1711 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000110; // iC= 1094 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010010; // iC=  978 
// vC = 14'b0000011001001011; // vC= 1611 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010001; // iC= 1105 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111110; // iC= 1214 
// vC = 14'b0000011001001111; // vC= 1615 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110101; // iC= 1013 
// vC = 14'b0000011100010001; // vC= 1809 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011011; // iC= 1115 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111110; // iC= 1214 
// vC = 14'b0000011010000111; // vC= 1671 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100110; // iC= 1062 
// vC = 14'b0000011010110010; // vC= 1714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011011; // iC= 1115 
// vC = 14'b0000011110000010; // vC= 1922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111011; // iC=  891 
// vC = 14'b0000011100110111; // vC= 1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100111; // iC= 1063 
// vC = 14'b0000011010010011; // vC= 1683 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000010; // iC= 1154 
// vC = 14'b0000011010111110; // vC= 1726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101001; // iC= 1129 
// vC = 14'b0000011101000110; // vC= 1862 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011000; // iC=  920 
// vC = 14'b0000011110000100; // vC= 1924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001100; // iC=  908 
// vC = 14'b0000011100101100; // vC= 1836 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000110; // iC= 1094 
// vC = 14'b0000011100000001; // vC= 1793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000110; // iC= 1030 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110110; // iC= 1014 
// vC = 14'b0000011101100110; // vC= 1894 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000100; // iC=  836 
// vC = 14'b0000011010001100; // vC= 1676 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110001; // iC= 1009 
// vC = 14'b0000011010100000; // vC= 1696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011110; // iC= 1054 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001011; // iC= 1099 
// vC = 14'b0000011010000110; // vC= 1670 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011110; // iC=  926 
// vC = 14'b0000011111000010; // vC= 1986 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100110; // iC=  806 
// vC = 14'b0000011110010110; // vC= 1942 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000100; // iC=  900 
// vC = 14'b0000011010011110; // vC= 1694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001100; // iC=  972 
// vC = 14'b0000011011111001; // vC= 1785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100001; // iC=  993 
// vC = 14'b0000011011000001; // vC= 1729 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111110; // iC= 1086 
// vC = 14'b0000011101000001; // vC= 1857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010011; // iC=  915 
// vC = 14'b0000011111001011; // vC= 1995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001100; // iC=  972 
// vC = 14'b0000011010101000; // vC= 1704 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b0000011110010000; // vC= 1936 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010011; // iC=  979 
// vC = 14'b0000011010111100; // vC= 1724 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000100; // iC=  836 
// vC = 14'b0000011110011010; // vC= 1946 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001111; // iC=  975 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101101; // iC= 1005 
// vC = 14'b0000011100001000; // vC= 1800 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011111; // iC=  735 
// vC = 14'b0000011010110001; // vC= 1713 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100101; // iC=  805 
// vC = 14'b0000011111000001; // vC= 1985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010111; // iC=  791 
// vC = 14'b0000011110001010; // vC= 1930 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011111; // iC=  991 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010100; // iC=  724 
// vC = 14'b0000011100011001; // vC= 1817 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011001; // iC=  985 
// vC = 14'b0000011100110110; // vC= 1846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000101; // iC=  965 
// vC = 14'b0000011101011110; // vC= 1886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011111; // iC=  991 
// vC = 14'b0000011101001101; // vC= 1869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001101; // iC=  973 
// vC = 14'b0000011110001101; // vC= 1933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101001; // iC=  745 
// vC = 14'b0000011110100111; // vC= 1959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001010; // iC=  650 
// vC = 14'b0000011110110100; // vC= 1972 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111100; // iC=  892 
// vC = 14'b0000011100010111; // vC= 1815 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011100; // iC=  732 
// vC = 14'b0000011111101101; // vC= 2029 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100110; // iC=  806 
// vC = 14'b0000100000011010; // vC= 2074 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100011; // iC=  803 
// vC = 14'b0000011100111011; // vC= 1851 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111011; // iC=  763 
// vC = 14'b0000011110011001; // vC= 1945 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100110; // iC=  614 
// vC = 14'b0000011110010110; // vC= 1942 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011111; // iC=  607 
// vC = 14'b0000100000011011; // vC= 2075 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110101; // iC=  885 
// vC = 14'b0000011101100000; // vC= 1888 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111011; // iC=  635 
// vC = 14'b0000011100100101; // vC= 1829 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011001; // iC=  665 
// vC = 14'b0000011111110010; // vC= 2034 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000101; // iC=  837 
// vC = 14'b0000011101110000; // vC= 1904 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101000; // iC=  872 
// vC = 14'b0000011111110101; // vC= 2037 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010100; // iC=  596 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110011; // iC=  755 
// vC = 14'b0000011110110000; // vC= 1968 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000001; // iC=  833 
// vC = 14'b0000100000011101; // vC= 2077 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000011; // iC=  579 
// vC = 14'b0000011101111111; // vC= 1919 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001001; // iC=  713 
// vC = 14'b0000011101010011; // vC= 1875 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010000; // iC=  592 
// vC = 14'b0000011111011001; // vC= 2009 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100010; // iC=  802 
// vC = 14'b0000100000010001; // vC= 2065 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011011; // iC=  795 
// vC = 14'b0000011100111101; // vC= 1853 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010001; // iC=  657 
// vC = 14'b0000011110110010; // vC= 1970 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111001; // iC=  761 
// vC = 14'b0000100001000010; // vC= 2114 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010111; // iC=  599 
// vC = 14'b0000011110000111; // vC= 1927 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110011; // iC=  499 
// vC = 14'b0000100000011001; // vC= 2073 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100101; // iC=  613 
// vC = 14'b0000011100100111; // vC= 1831 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101111; // iC=  751 
// vC = 14'b0000100000001100; // vC= 2060 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110101; // iC=  501 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001011; // iC=  523 
// vC = 14'b0000011100100111; // vC= 1831 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110111; // iC=  503 
// vC = 14'b0000011100110000; // vC= 1840 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101100; // iC=  620 
// vC = 14'b0000011101011110; // vC= 1886 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000101; // iC=  389 
// vC = 14'b0000011101000110; // vC= 1862 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001101; // iC=  589 
// vC = 14'b0000011110000100; // vC= 1924 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000110; // iC=  646 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100101; // iC=  485 
// vC = 14'b0000011110100000; // vC= 1952 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001100; // iC=  588 
// vC = 14'b0000011101011110; // vC= 1886 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101010; // iC=  490 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011000; // iC=  600 
// vC = 14'b0000100000110110; // vC= 2102 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101011; // iC=  427 
// vC = 14'b0000011111110110; // vC= 2038 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100101; // iC=  357 
// vC = 14'b0000011110000111; // vC= 1927 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011111; // iC=  351 
// vC = 14'b0000011101011101; // vC= 1885 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001101; // iC=  461 
// vC = 14'b0000011100111111; // vC= 1855 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100101; // iC=  293 
// vC = 14'b0000100000110001; // vC= 2097 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001001; // iC=  201 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000010; // iC=  386 
// vC = 14'b0000011110110100; // vC= 1972 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010110; // iC=  278 
// vC = 14'b0000011111101001; // vC= 2025 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111110; // iC=  190 
// vC = 14'b0000100001000011; // vC= 2115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000000; // iC=  256 
// vC = 14'b0000011100111001; // vC= 1849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100101; // iC=  357 
// vC = 14'b0000011111001100; // vC= 1996 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000110; // iC=  326 
// vC = 14'b0000011111110101; // vC= 2037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111010; // iC=  378 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110001; // iC=  113 
// vC = 14'b0000011101010101; // vC= 1877 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001100; // iC=  332 
// vC = 14'b0000100000101111; // vC= 2095 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100000; // iC=   32 
// vC = 14'b0000100000100010; // vC= 2082 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010110; // iC=  214 
// vC = 14'b0000011111011011; // vC= 2011 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010100; // iC=  212 
// vC = 14'b0000011101011001; // vC= 1881 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110110; // iC=  310 
// vC = 14'b0000011101001001; // vC= 1865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100111; // iC=  103 
// vC = 14'b0000011110000000; // vC= 1920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100000; // iC=   96 
// vC = 14'b0000011101010100; // vC= 1876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110110; // iC=  118 
// vC = 14'b0000011110101011; // vC= 1963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001001; // iC=   73 
// vC = 14'b0000100001110110; // vC= 2166 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111111; // iC=  191 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111110110; // iC=  -10 
// vC = 14'b0000011110010001; // vC= 1937 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100111; // iC=  103 
// vC = 14'b0000100000101111; // vC= 2095 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010101; // iC= -107 
// vC = 14'b0000011101010011; // vC= 1875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000110; // iC=  -58 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101111; // iC=  111 
// vC = 14'b0000100000100000; // vC= 2080 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011110; // iC=  -98 
// vC = 14'b0000100000000011; // vC= 2051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010101; // iC= -171 
// vC = 14'b0000100000000010; // vC= 2050 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101111; // iC= -145 
// vC = 14'b0000100000111011; // vC= 2107 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111011; // iC=   -5 
// vC = 14'b0000011101000101; // vC= 1861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001011; // iC= -181 
// vC = 14'b0000011111001000; // vC= 1992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001111; // iC= -305 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111101; // iC= -323 
// vC = 14'b0000011111001000; // vC= 1992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111110; // iC=  -66 
// vC = 14'b0000011110011010; // vC= 1946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010101101; // iC= -339 
// vC = 14'b0000011101001010; // vC= 1866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010110; // iC= -170 
// vC = 14'b0000011101101101; // vC= 1901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100100; // iC= -220 
// vC = 14'b0000011101010001; // vC= 1873 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100101; // iC= -347 
// vC = 14'b0000100001001111; // vC= 2127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100111; // iC= -409 
// vC = 14'b0000011111111011; // vC= 2043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001010; // iC= -246 
// vC = 14'b0000011100101101; // vC= 1837 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001110; // iC= -498 
// vC = 14'b0000011110111011; // vC= 1979 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011101; // iC= -355 
// vC = 14'b0000100001100100; // vC= 2148 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111011; // iC= -453 
// vC = 14'b0000100000100010; // vC= 2082 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110010; // iC= -398 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101100; // iC= -532 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010011; // iC= -365 
// vC = 14'b0000100000011010; // vC= 2074 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111110; // iC= -514 
// vC = 14'b0000011101011000; // vC= 1880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010100; // iC= -428 
// vC = 14'b0000011111001100; // vC= 1996 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010101; // iC= -491 
// vC = 14'b0000011110111100; // vC= 1980 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011010; // iC= -486 
// vC = 14'b0000011110111000; // vC= 1976 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111000; // iC= -712 
// vC = 14'b0000011101011100; // vC= 1884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001001; // iC= -567 
// vC = 14'b0000011111110001; // vC= 2033 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101110; // iC= -786 
// vC = 14'b0000011100010010; // vC= 1810 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100100; // iC= -668 
// vC = 14'b0000011101110010; // vC= 1906 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111010; // iC= -710 
// vC = 14'b0000011101100010; // vC= 1890 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110101; // iC= -651 
// vC = 14'b0000100001000101; // vC= 2117 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101100; // iC= -788 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111111; // iC= -705 
// vC = 14'b0000100000101111; // vC= 2095 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101101; // iC= -723 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011110; // iC= -930 
// vC = 14'b0000011100001100; // vC= 1804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011101; // iC= -739 
// vC = 14'b0000011110111001; // vC= 1977 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001100; // iC= -820 
// vC = 14'b0000011100110001; // vC= 1841 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010001; // iC= -751 
// vC = 14'b0000011111111010; // vC= 2042 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101010; // iC= -982 
// vC = 14'b0000011100010010; // vC= 1810 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101010; // iC= -854 
// vC = 14'b0000011100011001; // vC= 1817 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111111; // iC=-1025 
// vC = 14'b0000011111101100; // vC= 2028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011011; // iC=-1125 
// vC = 14'b0000011100000000; // vC= 1792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000000; // iC=-1088 
// vC = 14'b0000011111001001; // vC= 1993 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101011; // iC= -853 
// vC = 14'b0000011111100011; // vC= 2019 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100100; // iC=-1180 
// vC = 14'b0000011101100011; // vC= 1891 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010111; // iC= -937 
// vC = 14'b0000011100001111; // vC= 1807 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010111; // iC=-1001 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010110; // iC=-1066 
// vC = 14'b0000011111111011; // vC= 2043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010110; // iC=-1002 
// vC = 14'b0000011111010010; // vC= 2002 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001111; // iC=-1073 
// vC = 14'b0000011101100111; // vC= 1895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011000; // iC=-1192 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000100; // iC=-1148 
// vC = 14'b0000011111011111; // vC= 2015 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000101; // iC=-1147 
// vC = 14'b0000011011010001; // vC= 1745 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111101; // iC=-1347 
// vC = 14'b0000011101111100; // vC= 1916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111000; // iC=-1224 
// vC = 14'b0000011010101000; // vC= 1704 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110000; // iC=-1296 
// vC = 14'b0000011101100000; // vC= 1888 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101011; // iC=-1109 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111100; // iC=-1348 
// vC = 14'b0000011010011010; // vC= 1690 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100000; // iC=-1184 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000110; // iC=-1402 
// vC = 14'b0000011100010110; // vC= 1814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010001; // iC=-1199 
// vC = 14'b0000011101110001; // vC= 1905 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100000; // iC=-1504 
// vC = 14'b0000011010101110; // vC= 1710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111111; // iC=-1537 
// vC = 14'b0000011010100110; // vC= 1702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000010; // iC=-1534 
// vC = 14'b0000011010000001; // vC= 1665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011100; // iC=-1316 
// vC = 14'b0000011100001100; // vC= 1804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111110; // iC=-1282 
// vC = 14'b0000011010100011; // vC= 1699 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101100; // iC=-1492 
// vC = 14'b0000011100110101; // vC= 1845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101010; // iC=-1622 
// vC = 14'b0000011100111010; // vC= 1850 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010111; // iC=-1449 
// vC = 14'b0000011011000000; // vC= 1728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100000; // iC=-1632 
// vC = 14'b0000011011010001; // vC= 1745 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010010; // iC=-1390 
// vC = 14'b0000011101100000; // vC= 1888 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010010; // iC=-1454 
// vC = 14'b0000011001010000; // vC= 1616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111000; // iC=-1544 
// vC = 14'b0000011101000111; // vC= 1863 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001001; // iC=-1591 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100011; // iC=-1437 
// vC = 14'b0000011010011000; // vC= 1688 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111000; // iC=-1608 
// vC = 14'b0000011100101110; // vC= 1838 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111100; // iC=-1540 
// vC = 14'b0000011100111101; // vC= 1853 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101111; // iC=-1489 
// vC = 14'b0000011000110001; // vC= 1585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000110; // iC=-1658 
// vC = 14'b0000011000101011; // vC= 1579 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001000; // iC=-1592 
// vC = 14'b0000011000100011; // vC= 1571 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111111; // iC=-1729 
// vC = 14'b0000011001000000; // vC= 1600 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000110; // iC=-1658 
// vC = 14'b0000011011000001; // vC= 1729 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001101; // iC=-1523 
// vC = 14'b0000010111011010; // vC= 1498 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110001; // iC=-1551 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001010; // iC=-1846 
// vC = 14'b0000011001111110; // vC= 1662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101111; // iC=-1873 
// vC = 14'b0000011010000010; // vC= 1666 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010011; // iC=-1581 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011100; // iC=-1700 
// vC = 14'b0000011001000110; // vC= 1606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100100; // iC=-1692 
// vC = 14'b0000011010011000; // vC= 1688 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110111; // iC=-1609 
// vC = 14'b0000011001000110; // vC= 1606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b0000010111101100; // vC= 1516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001110; // iC=-1778 
// vC = 14'b0000011000001101; // vC= 1549 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011111; // iC=-1953 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011011; // iC=-1765 
// vC = 14'b0000010111010100; // vC= 1492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b0000011010101010; // vC= 1706 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101001; // iC=-1751 
// vC = 14'b0000010110100100; // vC= 1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101011; // iC=-1685 
// vC = 14'b0000010111011001; // vC= 1497 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100100; // iC=-1884 
// vC = 14'b0000010110100101; // vC= 1445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000110; // iC=-1850 
// vC = 14'b0000010101100011; // vC= 1379 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b0000011001010010; // vC= 1618 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010010; // iC=-1966 
// vC = 14'b0000010110010100; // vC= 1428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000011001111011; // vC= 1659 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010111; // iC=-1961 
// vC = 14'b0000010110000111; // vC= 1415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b0000010101000100; // vC= 1348 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000010101011100; // vC= 1372 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101101; // iC=-2067 
// vC = 14'b0000010110010001; // vC= 1425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b0000010110110011; // vC= 1459 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111101; // iC=-1795 
// vC = 14'b0000010100110100; // vC= 1332 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110001; // iC=-1871 
// vC = 14'b0000010100010001; // vC= 1297 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111111; // iC=-1793 
// vC = 14'b0000010100011110; // vC= 1310 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001101; // iC=-1779 
// vC = 14'b0000010110011000; // vC= 1432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100111; // iC=-1945 
// vC = 14'b0000010110111010; // vC= 1466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110000; // iC=-2000 
// vC = 14'b0000010101100100; // vC= 1380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b0000010011101011; // vC= 1259 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b0000010111101001; // vC= 1513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b0000010011101100; // vC= 1260 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000000; // iC=-1856 
// vC = 14'b0000010101110010; // vC= 1394 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101001; // iC=-2007 
// vC = 14'b0000010110010000; // vC= 1424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010000; // iC=-1904 
// vC = 14'b0000010111011001; // vC= 1497 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000010011000010; // vC= 1218 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110111; // iC=-2121 
// vC = 14'b0000010011010110; // vC= 1238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101011; // iC=-2133 
// vC = 14'b0000010110100100; // vC= 1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b0000010010100011; // vC= 1187 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000010101100011; // vC= 1379 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000100; // iC=-1852 
// vC = 14'b0000010011011000; // vC= 1240 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110111; // iC=-2121 
// vC = 14'b0000010011000111; // vC= 1223 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010011; // iC=-2093 
// vC = 14'b0000010010111000; // vC= 1208 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001100; // iC=-1908 
// vC = 14'b0000010001100001; // vC= 1121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100101; // iC=-2139 
// vC = 14'b0000010011100100; // vC= 1252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101100; // iC=-2132 
// vC = 14'b0000010010000001; // vC= 1153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b0000010010000010; // vC= 1154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000010001101010; // vC= 1130 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b0000010011010101; // vC= 1237 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111010; // iC=-2182 
// vC = 14'b0000010100011100; // vC= 1308 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b0000010100110100; // vC= 1332 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001001; // iC=-2167 
// vC = 14'b0000010100111110; // vC= 1342 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111101; // iC=-2115 
// vC = 14'b0000010010010110; // vC= 1174 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b0000010001010001; // vC= 1105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b0000010001110000; // vC= 1136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001100; // iC=-2164 
// vC = 14'b0000010010011010; // vC= 1178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b0000010000011001; // vC= 1049 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011011; // iC=-2149 
// vC = 14'b0000010011100010; // vC= 1250 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b0000010010010001; // vC= 1169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111010; // iC=-2182 
// vC = 14'b0000010001001011; // vC= 1099 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110000; // iC=-1936 
// vC = 14'b0000010010010010; // vC= 1170 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b0000010011011101; // vC= 1245 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100111; // iC=-2009 
// vC = 14'b0000010010011011; // vC= 1179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011000; // iC=-1896 
// vC = 14'b0000010010101011; // vC= 1195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110001; // iC=-1935 
// vC = 14'b0000010001010111; // vC= 1111 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b0000010000010011; // vC= 1043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010110; // iC=-2090 
// vC = 14'b0000001110100100; // vC=  932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000001110000111; // vC=  903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011110; // iC=-2082 
// vC = 14'b0000010001111111; // vC= 1151 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111101; // iC=-2115 
// vC = 14'b0000001101110111; // vC=  887 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b0000001111100010; // vC=  994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b0000001111000110; // vC=  966 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001100; // iC=-2164 
// vC = 14'b0000010010000000; // vC= 1152 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100110; // iC=-2074 
// vC = 14'b0000001110100100; // vC=  932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011010; // iC=-2022 
// vC = 14'b0000001101110100; // vC=  884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000010001100010; // vC= 1122 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100111; // iC=-2009 
// vC = 14'b0000010000011111; // vC= 1055 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000010001101001; // vC= 1129 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001111; // iC=-2097 
// vC = 14'b0000001100111101; // vC=  829 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000001111100000; // vC=  992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b0000001110111100; // vC=  956 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b0000001101110100; // vC=  884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000110; // iC=-2106 
// vC = 14'b0000001110101111; // vC=  943 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000010; // iC=-2174 
// vC = 14'b0000001100001111; // vC=  783 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101000; // iC=-2136 
// vC = 14'b0000001101011000; // vC=  856 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b0000001111110111; // vC= 1015 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100000; // iC=-2208 
// vC = 14'b0000001110010110; // vC=  918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000001111111101; // vC= 1021 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100011; // iC=-2141 
// vC = 14'b0000001011010101; // vC=  725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000001100001100; // vC=  780 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100110; // iC=-2138 
// vC = 14'b0000001011100010; // vC=  738 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b0000001100001000; // vC=  776 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101101; // iC=-2067 
// vC = 14'b0000001101100110; // vC=  870 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000001101011011; // vC=  859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b0000001101011001; // vC=  857 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100111; // iC=-2137 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001001; // iC=-2167 
// vC = 14'b0000001010100100; // vC=  676 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100100; // iC=-2204 
// vC = 14'b0000001100010111; // vC=  791 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010110; // iC=-2218 
// vC = 14'b0000001011110000; // vC=  752 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100100; // iC=-2204 
// vC = 14'b0000001001111101; // vC=  637 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111000; // iC=-2184 
// vC = 14'b0000001101010110; // vC=  854 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110100; // iC=-2252 
// vC = 14'b0000001100011000; // vC=  792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b0000001001100101; // vC=  613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000110; // iC=-2234 
// vC = 14'b0000001010000110; // vC=  646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010111; // iC=-1961 
// vC = 14'b0000001100100010; // vC=  802 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b0000001001111010; // vC=  634 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000100; // iC=-2236 
// vC = 14'b0000001010010011; // vC=  659 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000001010110100; // vC=  692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b0000001011010001; // vC=  721 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101110; // iC=-2258 
// vC = 14'b0000001001101100; // vC=  620 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000111; // iC=-2169 
// vC = 14'b0000001000111000; // vC=  568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b0000001001010111; // vC=  599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000000; // iC=-2176 
// vC = 14'b0000000111110001; // vC=  497 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100010; // iC=-2142 
// vC = 14'b0000001011000011; // vC=  707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010011; // iC=-2093 
// vC = 14'b0000001000111101; // vC=  573 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110110; // iC=-2250 
// vC = 14'b0000001100001110; // vC=  782 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b0000001000100000; // vC=  544 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111111; // iC=-2177 
// vC = 14'b0000001011000101; // vC=  709 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000001011000011; // vC=  707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001110; // iC=-2162 
// vC = 14'b0000001001101000; // vC=  616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b0000000111000010; // vC=  450 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b0000001001101000; // vC=  616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010010; // iC=-2222 
// vC = 14'b0000001010011111; // vC=  671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b0000001000100001; // vC=  545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001001; // iC=-2039 
// vC = 14'b0000001001100100; // vC=  612 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010100; // iC=-2220 
// vC = 14'b0000000111100001; // vC=  481 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001101; // iC=-2035 
// vC = 14'b0000001001011100; // vC=  604 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101101; // iC=-2259 
// vC = 14'b0000001010011011; // vC=  667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000110; // iC=-2170 
// vC = 14'b0000000101101011; // vC=  363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b0000001000010101; // vC=  533 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101010; // iC=-2198 
// vC = 14'b0000000111101100; // vC=  492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000011; // iC=-2173 
// vC = 14'b0000000110011000; // vC=  408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111111; // iC=-2113 
// vC = 14'b0000000101111011; // vC=  379 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100111; // iC=-2009 
// vC = 14'b0000000111100111; // vC=  487 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110111; // iC=-2185 
// vC = 14'b0000000111010000; // vC=  464 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000100; // iC=-2172 
// vC = 14'b0000000110101001; // vC=  425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111010; // iC=-2182 
// vC = 14'b0000000110111010; // vC=  442 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110001; // iC=-2063 
// vC = 14'b0000000101001000; // vC=  328 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110110; // iC=-1994 
// vC = 14'b0000001000000010; // vC=  514 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b0000000011111100; // vC=  252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011001; // iC=-2087 
// vC = 14'b0000000100111000; // vC=  312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000000111010110; // vC=  470 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101100; // iC=-2068 
// vC = 14'b0000000011110000; // vC=  240 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111011; // iC=-2245 
// vC = 14'b0000000101001111; // vC=  335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101010; // iC=-2134 
// vC = 14'b0000000111010011; // vC=  467 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011000; // iC=-2216 
// vC = 14'b0000000111011111; // vC=  479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b0000000111001110; // vC=  462 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010000; // iC=-2096 
// vC = 14'b0000000010110001; // vC=  177 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000000110010111; // vC=  407 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100111; // iC=-2201 
// vC = 14'b0000000100110011; // vC=  307 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110000; // iC=-2256 
// vC = 14'b0000000101000111; // vC=  327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010010; // iC=-2222 
// vC = 14'b0000000011001111; // vC=  207 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000000110000011; // vC=  387 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000000010100010; // vC=  162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000101; // iC=-2235 
// vC = 14'b0000000001100111; // vC=  103 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010100; // iC=-2220 
// vC = 14'b0000000110011100; // vC=  412 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b0000000001110111; // vC=  119 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001001; // iC=-2167 
// vC = 14'b0000000100001010; // vC=  266 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110000; // iC=-2128 
// vC = 14'b0000000010110100; // vC=  180 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000000001101010; // vC=  106 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110001; // iC=-1999 
// vC = 14'b0000000101010100; // vC=  340 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111111; // iC=-2177 
// vC = 14'b0000000010000101; // vC=  133 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011100; // iC=-2148 
// vC = 14'b0000000000110101; // vC=   53 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000000010110011; // vC=  179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000010; // iC=-2046 
// vC = 14'b0000000000111110; // vC=   62 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111100; // iC=-2180 
// vC = 14'b0000000010011100; // vC=  156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101110; // iC=-2130 
// vC = 14'b0000000010110110; // vC=  182 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b0000000000011100; // vC=   28 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111100; // iC=-2244 
// vC = 14'b0000000100100101; // vC=  293 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000000010001011; // vC=  139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110010; // iC=-2062 
// vC = 14'b0000000000110011; // vC=   51 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110001; // iC=-2063 
// vC = 14'b1111111111100100; // vC=  -28 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001100; // iC=-2164 
// vC = 14'b1111111111001000; // vC=  -56 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b0000000010100100; // vC=  164 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110001; // iC=-2127 
// vC = 14'b0000000010101000; // vC=  168 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101111; // iC=-2001 
// vC = 14'b0000000001101111; // vC=  111 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000000010001100; // vC=  140 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b1111111111001111; // vC=  -49 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000000000001111; // vC=   15 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b1111111110000101; // vC= -123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111100; // iC=-1924 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111001; // iC=-1991 
// vC = 14'b1111111111101100; // vC=  -20 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011101; // iC=-2083 
// vC = 14'b1111111111010110; // vC=  -42 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010111; // iC=-2217 
// vC = 14'b0000000000111101; // vC=   61 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b1111111110101001; // vC=  -87 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111111; // iC=-2177 
// vC = 14'b1111111110111101; // vC=  -67 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b1111111110111110; // vC=  -66 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011111; // iC=-2081 
// vC = 14'b0000000001101000; // vC=  104 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010111; // iC=-2217 
// vC = 14'b1111111111100101; // vC=  -27 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010111; // iC=-2153 
// vC = 14'b0000000000001100; // vC=   12 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001011; // iC=-1973 
// vC = 14'b1111111110010100; // vC= -108 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b1111111110001111; // vC= -113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100101; // iC=-2011 
// vC = 14'b1111111111000110; // vC=  -58 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b0000000000100111; // vC=   39 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011111; // iC=-2209 
// vC = 14'b1111111110001110; // vC= -114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b1111111100100111; // vC= -217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101001; // iC=-2135 
// vC = 14'b1111111101110010; // vC= -142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000000000100001; // vC=   33 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101000; // iC=-2136 
// vC = 14'b1111111110111110; // vC=  -66 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b1111111110001101; // vC= -115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b1111111110000100; // vC= -124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b1111111110100111; // vC=  -89 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100111; // iC=-1945 
// vC = 14'b1111111100001000; // vC= -248 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001110; // iC=-1906 
// vC = 14'b1111111111001011; // vC=  -53 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001001; // iC=-2167 
// vC = 14'b1111111010111111; // vC= -321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b1111111100110000; // vC= -208 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110000; // iC=-2128 
// vC = 14'b1111111010011011; // vC= -357 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101011; // iC=-2133 
// vC = 14'b1111111011110110; // vC= -266 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b1111111011101000; // vC= -280 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000101; // iC=-2107 
// vC = 14'b1111111101000000; // vC= -192 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111001; // iC=-2183 
// vC = 14'b1111111010100000; // vC= -352 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011000; // iC=-2024 
// vC = 14'b1111111100100101; // vC= -219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b1111111100111110; // vC= -194 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110011; // iC=-1997 
// vC = 14'b1111111010000110; // vC= -378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101100; // iC=-2132 
// vC = 14'b1111111010111101; // vC= -323 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001000; // iC=-2168 
// vC = 14'b1111111011001001; // vC= -311 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b1111111010110000; // vC= -336 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111100; // iC=-2116 
// vC = 14'b1111111000111111; // vC= -449 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001011; // iC=-2165 
// vC = 14'b1111111011011000; // vC= -296 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001111; // iC=-2161 
// vC = 14'b1111111010011011; // vC= -357 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101101; // iC=-2067 
// vC = 14'b1111111010000100; // vC= -380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b1111111100000111; // vC= -249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110001; // iC=-2063 
// vC = 14'b1111111100100101; // vC= -219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110010; // iC=-1934 
// vC = 14'b1111111100010110; // vC= -234 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b1111111000101110; // vC= -466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101011; // iC=-2069 
// vC = 14'b1111111001001000; // vC= -440 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b1111111001100100; // vC= -412 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011111; // iC=-2081 
// vC = 14'b1111111010111010; // vC= -326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b1111111001010100; // vC= -428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001001; // iC=-2039 
// vC = 14'b1111111011000011; // vC= -317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b1111111011101010; // vC= -278 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b1111111000000001; // vC= -511 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001001; // iC=-2039 
// vC = 14'b1111111001101011; // vC= -405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b1111111000111100; // vC= -452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011011; // iC=-2085 
// vC = 14'b1111111000011010; // vC= -486 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b1111111010001111; // vC= -369 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000110; // iC=-1850 
// vC = 14'b1111110110111001; // vC= -583 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100101; // iC=-2075 
// vC = 14'b1111111000000010; // vC= -510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b1111110110000011; // vC= -637 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000010; // iC=-2046 
// vC = 14'b1111111000110010; // vC= -462 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111010; // iC=-1798 
// vC = 14'b1111111000111110; // vC= -450 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b1111111001010101; // vC= -427 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000011; // iC=-1853 
// vC = 14'b1111111001100000; // vC= -416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100000; // iC=-2080 
// vC = 14'b1111111001011101; // vC= -419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b1111111010010000; // vC= -368 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100101; // iC=-2075 
// vC = 14'b1111111001100001; // vC= -415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b1111111001111010; // vC= -390 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010101; // iC=-1835 
// vC = 14'b1111110110000101; // vC= -635 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101010; // iC=-1814 
// vC = 14'b1111110111101000; // vC= -536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b1111110100101011; // vC= -725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101101; // iC=-1811 
// vC = 14'b1111110100100100; // vC= -732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000100; // iC=-1852 
// vC = 14'b1111110101001010; // vC= -694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b1111110111101100; // vC= -532 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b1111110111111111; // vC= -513 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b1111111000101100; // vC= -468 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b1111110011110101; // vC= -779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b1111110100001001; // vC= -759 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b1111110101111001; // vC= -647 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b1111110111000011; // vC= -573 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001000; // iC=-1784 
// vC = 14'b1111110110011101; // vC= -611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b1111110101100101; // vC= -667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010000; // iC=-1776 
// vC = 14'b1111110011010111; // vC= -809 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001110; // iC=-1842 
// vC = 14'b1111110111101010; // vC= -534 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010110; // iC=-1770 
// vC = 14'b1111110011111110; // vC= -770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b1111110111001111; // vC= -561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b1111110110111100; // vC= -580 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b1111110011011011; // vC= -805 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b1111110010011100; // vC= -868 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b1111110010011010; // vC= -870 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b1111110101100010; // vC= -670 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011001; // iC=-1895 
// vC = 14'b1111110010011101; // vC= -867 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011111; // iC=-1761 
// vC = 14'b1111110010101000; // vC= -856 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b1111110100110011; // vC= -717 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001110; // iC=-1714 
// vC = 14'b1111110110100101; // vC= -603 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010000; // iC=-1776 
// vC = 14'b1111110100011101; // vC= -739 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011111; // iC=-1761 
// vC = 14'b1111110101111101; // vC= -643 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011000; // iC=-1896 
// vC = 14'b1111110011000100; // vC= -828 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100001; // iC=-1887 
// vC = 14'b1111110101100110; // vC= -666 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b1111110001101011; // vC= -917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011010; // iC=-1766 
// vC = 14'b1111110010110110; // vC= -842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b1111110010100110; // vC= -858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b1111110001100001; // vC= -927 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b1111110010011001; // vC= -871 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101011; // iC=-1877 
// vC = 14'b1111110010111101; // vC= -835 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010100; // iC=-1772 
// vC = 14'b1111110010011010; // vC= -870 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b1111110000110111; // vC= -969 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000010; // iC=-1790 
// vC = 14'b1111110100000100; // vC= -764 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111011; // iC=-1733 
// vC = 14'b1111110000000011; // vC=-1021 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110100; // iC=-1740 
// vC = 14'b1111110100010100; // vC= -748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b1111110000100011; // vC= -989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001000; // iC=-1720 
// vC = 14'b1111110000100011; // vC= -989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111001; // iC=-1927 
// vC = 14'b1111110010111001; // vC= -839 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b1111110001111010; // vC= -902 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000001; // iC=-1663 
// vC = 14'b1111110010110011; // vC= -845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010101; // iC=-1771 
// vC = 14'b1111110001110110; // vC= -906 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001111; // iC=-1841 
// vC = 14'b1111110011110110; // vC= -778 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101101; // iC=-1811 
// vC = 14'b1111101110111111; // vC=-1089 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101000; // iC=-1688 
// vC = 14'b1111110010100110; // vC= -858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110110; // iC=-1738 
// vC = 14'b1111110000001000; // vC=-1016 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b1111110000110011; // vC= -973 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001110; // iC=-1586 
// vC = 14'b1111101111000101; // vC=-1083 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b1111101110110111; // vC=-1097 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100010; // iC=-1758 
// vC = 14'b1111101110011101; // vC=-1123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101111; // iC=-1681 
// vC = 14'b1111101111100001; // vC=-1055 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b1111110001101101; // vC= -915 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000001; // iC=-1791 
// vC = 14'b1111110001101010; // vC= -918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011000; // iC=-1768 
// vC = 14'b1111101111000001; // vC=-1087 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000011; // iC=-1661 
// vC = 14'b1111101111100111; // vC=-1049 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010010; // iC=-1582 
// vC = 14'b1111101110101100; // vC=-1108 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100011; // iC=-1821 
// vC = 14'b1111110010010101; // vC= -875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000110; // iC=-1850 
// vC = 14'b1111101101010011; // vC=-1197 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011101; // iC=-1763 
// vC = 14'b1111101110111100; // vC=-1092 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101110; // iC=-1810 
// vC = 14'b1111101111110010; // vC=-1038 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011011; // iC=-1829 
// vC = 14'b1111101111011001; // vC=-1063 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011010; // iC=-1574 
// vC = 14'b1111110001110010; // vC= -910 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100011; // iC=-1565 
// vC = 14'b1111110000001111; // vC=-1009 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100111; // iC=-1625 
// vC = 14'b1111110001010011; // vC= -941 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100000; // iC=-1568 
// vC = 14'b1111101100110011; // vC=-1229 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100001; // iC=-1567 
// vC = 14'b1111101111110110; // vC=-1034 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001111; // iC=-1521 
// vC = 14'b1111101110000111; // vC=-1145 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011100; // iC=-1508 
// vC = 14'b1111101111101010; // vC=-1046 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111110; // iC=-1666 
// vC = 14'b1111101101011000; // vC=-1192 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101101; // iC=-1811 
// vC = 14'b1111101110111010; // vC=-1094 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b1111101111100011; // vC=-1053 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001010; // iC=-1718 
// vC = 14'b1111101101111111; // vC=-1153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110000; // iC=-1488 
// vC = 14'b1111110000011110; // vC= -994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000010; // iC=-1534 
// vC = 14'b1111101111011000; // vC=-1064 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101011; // iC=-1749 
// vC = 14'b1111101101110000; // vC=-1168 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001011; // iC=-1525 
// vC = 14'b1111110000010000; // vC=-1008 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000100; // iC=-1660 
// vC = 14'b1111101100110100; // vC=-1228 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110010; // iC=-1678 
// vC = 14'b1111101110110010; // vC=-1102 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101011; // iC=-1685 
// vC = 14'b1111101111111110; // vC=-1026 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001110; // iC=-1522 
// vC = 14'b1111101111100000; // vC=-1056 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011001; // iC=-1767 
// vC = 14'b1111101110111111; // vC=-1089 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111010; // iC=-1478 
// vC = 14'b1111101110100001; // vC=-1119 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010000; // iC=-1520 
// vC = 14'b1111101100010110; // vC=-1258 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000000; // iC=-1664 
// vC = 14'b1111101011000011; // vC=-1341 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100101; // iC=-1627 
// vC = 14'b1111101010101111; // vC=-1361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110010; // iC=-1678 
// vC = 14'b1111101100101100; // vC=-1236 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000111; // iC=-1465 
// vC = 14'b1111101101000000; // vC=-1216 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010100; // iC=-1580 
// vC = 14'b1111101101110100; // vC=-1164 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110010; // iC=-1678 
// vC = 14'b1111101011011010; // vC=-1318 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101111; // iC=-1617 
// vC = 14'b1111101001111001; // vC=-1415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001100; // iC=-1460 
// vC = 14'b1111101100110111; // vC=-1225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001011; // iC=-1717 
// vC = 14'b1111101101101111; // vC=-1169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110000; // iC=-1488 
// vC = 14'b1111101001110101; // vC=-1419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100010; // iC=-1630 
// vC = 14'b1111101101101101; // vC=-1171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000111; // iC=-1657 
// vC = 14'b1111101011000100; // vC=-1340 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010110; // iC=-1450 
// vC = 14'b1111101100100000; // vC=-1248 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111011; // iC=-1669 
// vC = 14'b1111101010101100; // vC=-1364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100110; // iC=-1434 
// vC = 14'b1111101100010101; // vC=-1259 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010000; // iC=-1392 
// vC = 14'b1111101010101100; // vC=-1364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110001; // iC=-1679 
// vC = 14'b1111101001001010; // vC=-1462 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010101; // iC=-1643 
// vC = 14'b1111101001100111; // vC=-1433 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110010; // iC=-1358 
// vC = 14'b1111101011001101; // vC=-1331 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100101; // iC=-1627 
// vC = 14'b1111101001101111; // vC=-1425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110101; // iC=-1611 
// vC = 14'b1111101011100000; // vC=-1312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100010; // iC=-1566 
// vC = 14'b1111101011110110; // vC=-1290 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110110; // iC=-1418 
// vC = 14'b1111101001100101; // vC=-1435 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010101; // iC=-1643 
// vC = 14'b1111101100101010; // vC=-1238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001100; // iC=-1396 
// vC = 14'b1111101100011011; // vC=-1253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100101; // iC=-1371 
// vC = 14'b1111101100010110; // vC=-1258 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100011; // iC=-1501 
// vC = 14'b1111101011010111; // vC=-1321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110001; // iC=-1359 
// vC = 14'b1111101100101000; // vC=-1240 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010000; // iC=-1392 
// vC = 14'b1111101001001111; // vC=-1457 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001101; // iC=-1395 
// vC = 14'b1111100111101001; // vC=-1559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101101; // iC=-1363 
// vC = 14'b1111101100011101; // vC=-1251 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010110; // iC=-1450 
// vC = 14'b1111101001001001; // vC=-1463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100100; // iC=-1436 
// vC = 14'b1111101000010101; // vC=-1515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101100; // iC=-1428 
// vC = 14'b1111101010001110; // vC=-1394 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010001; // iC=-1583 
// vC = 14'b1111100111001011; // vC=-1589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000101; // iC=-1467 
// vC = 14'b1111101011010010; // vC=-1326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101000; // iC=-1560 
// vC = 14'b1111100111101100; // vC=-1556 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100110; // iC=-1306 
// vC = 14'b1111101011100000; // vC=-1312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011111; // iC=-1249 
// vC = 14'b1111100110110111; // vC=-1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001010; // iC=-1526 
// vC = 14'b1111101000000001; // vC=-1535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100110; // iC=-1498 
// vC = 14'b1111100111100000; // vC=-1568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111011; // iC=-1413 
// vC = 14'b1111101000100100; // vC=-1500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010111; // iC=-1449 
// vC = 14'b1111100111000010; // vC=-1598 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000101; // iC=-1403 
// vC = 14'b1111101011010001; // vC=-1327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010010; // iC=-1518 
// vC = 14'b1111101011000110; // vC=-1338 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101110; // iC=-1362 
// vC = 14'b1111100111100011; // vC=-1565 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001110; // iC=-1458 
// vC = 14'b1111100110101110; // vC=-1618 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001101; // iC=-1203 
// vC = 14'b1111101001001011; // vC=-1461 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111011; // iC=-1285 
// vC = 14'b1111100111110010; // vC=-1550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100010; // iC=-1502 
// vC = 14'b1111101001100011; // vC=-1437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110100; // iC=-1356 
// vC = 14'b1111101010010111; // vC=-1385 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101001; // iC=-1367 
// vC = 14'b1111101001110100; // vC=-1420 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001000; // iC=-1464 
// vC = 14'b1111101001000000; // vC=-1472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101000; // iC=-1432 
// vC = 14'b1111101000101011; // vC=-1493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100010; // iC=-1182 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001001; // iC=-1399 
// vC = 14'b1111100111110110; // vC=-1546 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001010; // iC=-1206 
// vC = 14'b1111101000100011; // vC=-1501 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010100; // iC=-1388 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010010; // iC=-1390 
// vC = 14'b1111100110011111; // vC=-1633 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000010; // iC=-1214 
// vC = 14'b1111101000111010; // vC=-1478 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000000; // iC=-1152 
// vC = 14'b1111100111111000; // vC=-1544 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111110; // iC=-1410 
// vC = 14'b1111100110001001; // vC=-1655 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000011; // iC=-1341 
// vC = 14'b1111101000110010; // vC=-1486 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000101; // iC=-1339 
// vC = 14'b1111101001000110; // vC=-1466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111100; // iC=-1284 
// vC = 14'b1111100100111010; // vC=-1734 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011100; // iC=-1124 
// vC = 14'b1111100100110111; // vC=-1737 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000001; // iC=-1407 
// vC = 14'b1111100100101111; // vC=-1745 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011001; // iC=-1255 
// vC = 14'b1111100110110010; // vC=-1614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011000; // iC=-1320 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110110; // iC=-1162 
// vC = 14'b1111100100011010; // vC=-1766 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010010; // iC=-1198 
// vC = 14'b1111101001001001; // vC=-1463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011000; // iC=-1192 
// vC = 14'b1111100100000101; // vC=-1787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011111; // iC=-1377 
// vC = 14'b1111100111000101; // vC=-1595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011110; // iC=-1122 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110100; // iC=-1228 
// vC = 14'b1111100100001001; // vC=-1783 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111100; // iC=-1220 
// vC = 14'b1111101000100110; // vC=-1498 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000000; // iC=-1216 
// vC = 14'b1111100101001110; // vC=-1714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111011; // iC=-1349 
// vC = 14'b1111100111011000; // vC=-1576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000011; // iC=-1277 
// vC = 14'b1111100100011011; // vC=-1765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000111; // iC=-1337 
// vC = 14'b1111100011100001; // vC=-1823 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101001; // iC=-1047 
// vC = 14'b1111100101011110; // vC=-1698 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011101; // iC=-1187 
// vC = 14'b1111100100000101; // vC=-1787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111111; // iC=-1089 
// vC = 14'b1111100110101000; // vC=-1624 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001000; // iC=-1080 
// vC = 14'b1111100111111111; // vC=-1537 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001101; // iC=-1011 
// vC = 14'b1111100100001100; // vC=-1780 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001100; // iC=-1076 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110010; // iC=-1038 
// vC = 14'b1111100100101011; // vC=-1749 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111101; // iC=-1091 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011001; // iC=-1191 
// vC = 14'b1111100110100100; // vC=-1628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111101; // iC=-1091 
// vC = 14'b1111100101111100; // vC=-1668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110000; // iC= -976 
// vC = 14'b1111100100110010; // vC=-1742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110111; // iC= -969 
// vC = 14'b1111100110100101; // vC=-1627 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000010; // iC= -958 
// vC = 14'b1111100011011001; // vC=-1831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100100; // iC= -988 
// vC = 14'b1111100101010001; // vC=-1711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011001; // iC=-1063 
// vC = 14'b1111100011100111; // vC=-1817 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001000; // iC= -952 
// vC = 14'b1111100111001000; // vC=-1592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000010; // iC= -958 
// vC = 14'b1111100011001010; // vC=-1846 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100111; // iC= -921 
// vC = 14'b1111100100010010; // vC=-1774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110000; // iC= -976 
// vC = 14'b1111100010111110; // vC=-1858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101011; // iC=-1045 
// vC = 14'b1111100010111100; // vC=-1860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101001; // iC=-1111 
// vC = 14'b1111100110000100; // vC=-1660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111000; // iC=-1096 
// vC = 14'b1111100100010110; // vC=-1770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110111; // iC=-1033 
// vC = 14'b1111100011001101; // vC=-1843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100110; // iC=-1050 
// vC = 14'b1111100010110010; // vC=-1870 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000001; // iC=-1023 
// vC = 14'b1111100110010011; // vC=-1645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101011; // iC= -917 
// vC = 14'b1111100101000010; // vC=-1726 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110010; // iC=-1038 
// vC = 14'b1111100001111100; // vC=-1924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001010; // iC=-1014 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000100; // iC= -892 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110110; // iC= -842 
// vC = 14'b1111100010000010; // vC=-1918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001101; // iC= -883 
// vC = 14'b1111100011110100; // vC=-1804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110101; // iC= -843 
// vC = 14'b1111100100111101; // vC=-1731 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100000; // iC=-1056 
// vC = 14'b1111100010110101; // vC=-1867 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001000; // iC=-1016 
// vC = 14'b1111100010100111; // vC=-1881 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001010; // iC= -822 
// vC = 14'b1111100001010100; // vC=-1964 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011100; // iC= -996 
// vC = 14'b1111100011100100; // vC=-1820 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111000; // iC=-1096 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010011; // iC= -941 
// vC = 14'b1111100001100011; // vC=-1949 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011100; // iC= -996 
// vC = 14'b1111100100000001; // vC=-1791 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001010; // iC= -822 
// vC = 14'b1111100011101011; // vC=-1813 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001111; // iC= -881 
// vC = 14'b1111100010011111; // vC=-1889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101001; // iC=-1047 
// vC = 14'b1111100001010010; // vC=-1966 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111111; // iC= -769 
// vC = 14'b1111100000100110; // vC=-2010 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111111; // iC=-1025 
// vC = 14'b1111100100001110; // vC=-1778 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110111; // iC= -841 
// vC = 14'b1111100100111110; // vC=-1730 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011101; // iC= -995 
// vC = 14'b1111100010111101; // vC=-1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101111; // iC= -785 
// vC = 14'b1111100001011011; // vC=-1957 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011110; // iC= -738 
// vC = 14'b1111100010011110; // vC=-1890 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b1111100011100010; // vC=-1822 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001000; // iC= -824 
// vC = 14'b1111100100101100; // vC=-1748 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110010; // iC= -718 
// vC = 14'b1111100000010010; // vC=-2030 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011101; // iC= -931 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011000; // iC= -808 
// vC = 14'b1111100011101010; // vC=-1814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110100; // iC= -908 
// vC = 14'b1111100010001111; // vC=-1905 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110111; // iC= -777 
// vC = 14'b1111100100001100; // vC=-1780 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100101; // iC= -987 
// vC = 14'b1111100001011101; // vC=-1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100010; // iC= -734 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001011; // iC= -821 
// vC = 14'b1111100000111001; // vC=-1991 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001001; // iC= -823 
// vC = 14'b1111100011001110; // vC=-1842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011001; // iC= -871 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111000; // iC= -840 
// vC = 14'b1111011111101100; // vC=-2068 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100011; // iC= -797 
// vC = 14'b1111100011011011; // vC=-1829 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100010; // iC= -798 
// vC = 14'b1111100010110100; // vC=-1868 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010001; // iC= -687 
// vC = 14'b1111100010010010; // vC=-1902 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101101; // iC= -723 
// vC = 14'b1111100001010100; // vC=-1964 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001100; // iC= -756 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101000; // iC= -920 
// vC = 14'b1111100010100001; // vC=-1887 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001110; // iC= -818 
// vC = 14'b1111100100000101; // vC=-1787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100000; // iC= -800 
// vC = 14'b1111100000001111; // vC=-2033 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010000; // iC= -688 
// vC = 14'b1111011111100100; // vC=-2076 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001111; // iC= -689 
// vC = 14'b1111100011010001; // vC=-1839 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110001; // iC= -591 
// vC = 14'b1111100010101000; // vC=-1880 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000101; // iC= -763 
// vC = 14'b1111100000111100; // vC=-1988 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000100; // iC= -636 
// vC = 14'b1111100001110000; // vC=-1936 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110101; // iC= -651 
// vC = 14'b1111100011101001; // vC=-1815 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101110; // iC= -850 
// vC = 14'b1111100000110110; // vC=-1994 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010100; // iC= -556 
// vC = 14'b1111011111011101; // vC=-2083 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101101; // iC= -531 
// vC = 14'b1111100011000011; // vC=-1853 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010010; // iC= -814 
// vC = 14'b1111100011011101; // vC=-1827 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011000; // iC= -616 
// vC = 14'b1111011111000101; // vC=-2107 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100111; // iC= -729 
// vC = 14'b1111100011010100; // vC=-1836 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110111; // iC= -713 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011101; // iC= -611 
// vC = 14'b1111011111011001; // vC=-2087 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011011; // iC= -549 
// vC = 14'b1111011111000100; // vC=-2108 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000000100; // iC= -508 
// vC = 14'b1111011110101110; // vC=-2130 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111000; // iC= -776 
// vC = 14'b1111011111101010; // vC=-2070 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000000; // iC= -576 
// vC = 14'b1111011110100010; // vC=-2142 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001001; // iC= -759 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101010; // iC= -598 
// vC = 14'b1111100000101000; // vC=-2008 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010011; // iC= -621 
// vC = 14'b1111100010000100; // vC=-1916 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011011; // iC= -485 
// vC = 14'b1111100010001011; // vC=-1909 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010100; // iC= -428 
// vC = 14'b1111100010101011; // vC=-1877 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110010; // iC= -398 
// vC = 14'b1111100000011010; // vC=-2022 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010001; // iC= -623 
// vC = 14'b1111011111011100; // vC=-2084 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011100; // iC= -420 
// vC = 14'b1111011111110001; // vC=-2063 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010100; // iC= -428 
// vC = 14'b1111100010110100; // vC=-1868 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100101; // iC= -667 
// vC = 14'b1111100011000110; // vC=-1850 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101111; // iC= -593 
// vC = 14'b1111100001010000; // vC=-1968 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110111; // iC= -329 
// vC = 14'b1111100000001000; // vC=-2040 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001101; // iC= -627 
// vC = 14'b1111100010100011; // vC=-1885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001111; // iC= -561 
// vC = 14'b1111100001010010; // vC=-1966 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011000; // iC= -424 
// vC = 14'b1111100001110101; // vC=-1931 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001001; // iC= -439 
// vC = 14'b1111100000000101; // vC=-2043 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001100; // iC= -500 
// vC = 14'b1111100001001000; // vC=-1976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011111100; // iC= -260 
// vC = 14'b1111011101111111; // vC=-2177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001011; // iC= -309 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010010; // iC= -430 
// vC = 14'b1111100000011101; // vC=-2019 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000000; // iC= -384 
// vC = 14'b1111100001011001; // vC=-1959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110100; // iC= -396 
// vC = 14'b1111011110100000; // vC=-2144 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110000; // iC= -464 
// vC = 14'b1111011111101000; // vC=-2072 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000011; // iC= -189 
// vC = 14'b1111100010110111; // vC=-1865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111010; // iC= -134 
// vC = 14'b1111100000001111; // vC=-2033 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011110; // iC= -354 
// vC = 14'b1111011101111010; // vC=-2182 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101001; // iC= -407 
// vC = 14'b1111100010011011; // vC=-1893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100100; // iC= -156 
// vC = 14'b1111011110110011; // vC=-2125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011110111; // iC= -265 
// vC = 14'b1111011110111101; // vC=-2115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100001; // iC= -351 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111010; // iC= -198 
// vC = 14'b1111011111001001; // vC=-2103 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101101; // iC= -147 
// vC = 14'b1111100001100111; // vC=-1945 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011110101; // iC= -267 
// vC = 14'b1111100010101000; // vC=-1880 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010110; // iC= -170 
// vC = 14'b1111100000111111; // vC=-1985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101010110; // iC= -170 
// vC = 14'b1111011111001011; // vC=-2101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000010; // iC= -126 
// vC = 14'b1111011101111011; // vC=-2181 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100111; // iC=  -25 
// vC = 14'b1111011111111001; // vC=-2055 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111111; // iC= -193 
// vC = 14'b1111100000011100; // vC=-2020 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111101; // iC=  -67 
// vC = 14'b1111011111100011; // vC=-2077 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010111; // iC=  151 
// vC = 14'b1111011111001111; // vC=-2097 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001000; // iC=  -56 
// vC = 14'b1111011111101001; // vC=-2071 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000100; // iC=  -60 
// vC = 14'b1111011111101101; // vC=-2067 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000101; // iC=  -59 
// vC = 14'b1111011111010100; // vC=-2092 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111110100; // iC=  -12 
// vC = 14'b1111100001011010; // vC=-1958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011001; // iC=   25 
// vC = 14'b1111011101110111; // vC=-2185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111001; // iC=  185 
// vC = 14'b1111100000110011; // vC=-1997 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001111; // iC=   79 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010001; // iC=   81 
// vC = 14'b1111100000110111; // vC=-1993 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010011; // iC=   83 
// vC = 14'b1111100000011001; // vC=-2023 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010010; // iC=  338 
// vC = 14'b1111011111111101; // vC=-2051 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100101; // iC=  165 
// vC = 14'b1111100000000011; // vC=-2045 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010000; // iC=  272 
// vC = 14'b1111100001101000; // vC=-1944 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011101; // iC=  349 
// vC = 14'b1111100001110110; // vC=-1930 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111101; // iC=  381 
// vC = 14'b1111011110011111; // vC=-2145 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010110; // iC=  342 
// vC = 14'b1111011110001110; // vC=-2162 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010001; // iC=  529 
// vC = 14'b1111100001011111; // vC=-1953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011101; // iC=  349 
// vC = 14'b1111100001011010; // vC=-1958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001001; // iC=  265 
// vC = 14'b1111011111010110; // vC=-2090 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001110; // iC=  334 
// vC = 14'b1111011110110011; // vC=-2125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000000; // iC=  448 
// vC = 14'b1111011111011111; // vC=-2081 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001111; // iC=  527 
// vC = 14'b1111100010011111; // vC=-1889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110000; // iC=  624 
// vC = 14'b1111100001001101; // vC=-1971 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011111; // iC=  479 
// vC = 14'b1111011110111101; // vC=-2115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010111; // iC=  407 
// vC = 14'b1111100011001100; // vC=-1844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000110; // iC=  582 
// vC = 14'b1111011111110111; // vC=-2057 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010101; // iC=  469 
// vC = 14'b1111011111001100; // vC=-2100 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111001; // iC=  633 
// vC = 14'b1111100000100101; // vC=-2011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111101; // iC=  573 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111011; // iC=  827 
// vC = 14'b1111011111010101; // vC=-2091 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100001; // iC=  545 
// vC = 14'b1111100011100001; // vC=-1823 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000001; // iC=  641 
// vC = 14'b1111100000000111; // vC=-2041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101111; // iC=  751 
// vC = 14'b1111100000001100; // vC=-2036 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111101; // iC=  893 
// vC = 14'b1111100001110110; // vC=-1930 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001110; // iC=  910 
// vC = 14'b1111100010101001; // vC=-1879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101000; // iC=  744 
// vC = 14'b1111100010111010; // vC=-1862 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001111; // iC=  975 
// vC = 14'b1111100000011000; // vC=-2024 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011100; // iC=  924 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111111; // iC= 1023 
// vC = 14'b1111100000010000; // vC=-2032 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100110; // iC=  870 
// vC = 14'b1111100010110011; // vC=-1869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110101; // iC= 1013 
// vC = 14'b1111100011110001; // vC=-1807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001000; // iC= 1096 
// vC = 14'b1111100010011010; // vC=-1894 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000000; // iC=  896 
// vC = 14'b1111100010001100; // vC=-1908 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010001; // iC=  913 
// vC = 14'b1111100001010101; // vC=-1963 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010110; // iC= 1046 
// vC = 14'b1111100001100110; // vC=-1946 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101010; // iC=  938 
// vC = 14'b1111100000110111; // vC=-1993 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001101; // iC= 1165 
// vC = 14'b1111100000000011; // vC=-2045 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100000; // iC= 1184 
// vC = 14'b1111100001001011; // vC=-1973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111101; // iC= 1213 
// vC = 14'b1111100100001010; // vC=-1782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111010; // iC= 1082 
// vC = 14'b1111100001000011; // vC=-1981 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000101; // iC= 1029 
// vC = 14'b1111100100100000; // vC=-1760 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111011; // iC= 1275 
// vC = 14'b1111100100000110; // vC=-1786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100101; // iC= 1189 
// vC = 14'b1111100010100000; // vC=-1888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111010; // iC= 1338 
// vC = 14'b1111100101001001; // vC=-1719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010001; // iC= 1233 
// vC = 14'b1111100001011011; // vC=-1957 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001001; // iC= 1353 
// vC = 14'b1111100000100001; // vC=-2015 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101111; // iC= 1135 
// vC = 14'b1111100000100110; // vC=-2010 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000111; // iC= 1415 
// vC = 14'b1111100001011001; // vC=-1959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100111; // iC= 1191 
// vC = 14'b1111100101011101; // vC=-1699 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000010; // iC= 1282 
// vC = 14'b1111100011001010; // vC=-1846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000101; // iC= 1413 
// vC = 14'b1111100000111100; // vC=-1988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010011; // iC= 1363 
// vC = 14'b1111100001110111; // vC=-1929 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110110; // iC= 1270 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000011; // iC= 1283 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111010; // iC= 1274 
// vC = 14'b1111100010111111; // vC=-1857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110000; // iC= 1392 
// vC = 14'b1111100110001010; // vC=-1654 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000100; // iC= 1540 
// vC = 14'b1111100001111001; // vC=-1927 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100010; // iC= 1570 
// vC = 14'b1111100110100001; // vC=-1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111001; // iC= 1465 
// vC = 14'b1111100101011111; // vC=-1697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110001; // iC= 1521 
// vC = 14'b1111100011000100; // vC=-1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001001; // iC= 1353 
// vC = 14'b1111100011111110; // vC=-1794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000111; // iC= 1607 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110010; // iC= 1394 
// vC = 14'b1111100100011010; // vC=-1766 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111011; // iC= 1467 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111001; // iC= 1401 
// vC = 14'b1111100010100000; // vC=-1888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110001; // iC= 1649 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010001; // iC= 1617 
// vC = 14'b1111100111100101; // vC=-1563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111010; // iC= 1530 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100111; // iC= 1575 
// vC = 14'b1111100101001010; // vC=-1718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110111; // iC= 1591 
// vC = 14'b1111100100001110; // vC=-1778 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000001; // iC= 1601 
// vC = 14'b1111100101101010; // vC=-1686 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010111; // iC= 1623 
// vC = 14'b1111100101010000; // vC=-1712 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111010; // iC= 1594 
// vC = 14'b1111100101010011; // vC=-1709 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100110; // iC= 1702 
// vC = 14'b1111100100110100; // vC=-1740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110111; // iC= 1591 
// vC = 14'b1111100111111100; // vC=-1540 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101111; // iC= 1711 
// vC = 14'b1111100100111100; // vC=-1732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110010; // iC= 1650 
// vC = 14'b1111100110100001; // vC=-1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011110; // iC= 1694 
// vC = 14'b1111100110010100; // vC=-1644 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000101; // iC= 1669 
// vC = 14'b1111101000010010; // vC=-1518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110101; // iC= 1909 
// vC = 14'b1111100100101000; // vC=-1752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100111; // iC= 1767 
// vC = 14'b1111101000001001; // vC=-1527 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001000; // iC= 1928 
// vC = 14'b1111100110011010; // vC=-1638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011100; // iC= 1948 
// vC = 14'b1111100110001011; // vC=-1653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100111; // iC= 1831 
// vC = 14'b1111100100101111; // vC=-1745 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111010; // iC= 1850 
// vC = 14'b1111101000100010; // vC=-1502 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001101; // iC= 1805 
// vC = 14'b1111100101010000; // vC=-1712 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001110; // iC= 1870 
// vC = 14'b1111101000010100; // vC=-1516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011100; // iC= 1884 
// vC = 14'b1111100101010011; // vC=-1709 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111111; // iC= 1791 
// vC = 14'b1111100110110001; // vC=-1615 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b1111100110100001; // vC=-1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b1111101001110001; // vC=-1423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111000; // iC= 1720 
// vC = 14'b1111101010010011; // vC=-1389 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001100; // iC= 1804 
// vC = 14'b1111100111010100; // vC=-1580 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b1111100111011101; // vC=-1571 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000010; // iC= 1858 
// vC = 14'b1111101010001101; // vC=-1395 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100111; // iC= 1895 
// vC = 14'b1111100111011010; // vC=-1574 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111011; // iC= 1915 
// vC = 14'b1111101000010000; // vC=-1520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b1111100111111101; // vC=-1539 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010101; // iC= 1877 
// vC = 14'b1111101010101011; // vC=-1365 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000111; // iC= 2055 
// vC = 14'b1111101010011011; // vC=-1381 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110111; // iC= 1911 
// vC = 14'b1111100111001110; // vC=-1586 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b1111101001111100; // vC=-1412 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111001; // iC= 1849 
// vC = 14'b1111101001111101; // vC=-1411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000011; // iC= 1859 
// vC = 14'b1111101010011001; // vC=-1383 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b1111101011111001; // vC=-1287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b1111101010110110; // vC=-1354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011010; // iC= 1818 
// vC = 14'b1111101001110001; // vC=-1423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b1111101011111000; // vC=-1288 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101100; // iC= 2092 
// vC = 14'b1111101010010101; // vC=-1387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110011; // iC= 1971 
// vC = 14'b1111101101000011; // vC=-1213 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b1111101011011000; // vC=-1320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111101; // iC= 2045 
// vC = 14'b1111101100101110; // vC=-1234 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110111; // iC= 1847 
// vC = 14'b1111101100110010; // vC=-1230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110010; // iC= 1842 
// vC = 14'b1111101001010001; // vC=-1455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000000; // iC= 2112 
// vC = 14'b1111101011000101; // vC=-1339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011111; // iC= 2079 
// vC = 14'b1111101010100100; // vC=-1372 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b1111101101111000; // vC=-1160 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011011; // iC= 1947 
// vC = 14'b1111101001111010; // vC=-1414 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011010; // iC= 2138 
// vC = 14'b1111101010110110; // vC=-1354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b1111101011110011; // vC=-1293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b1111101010111111; // vC=-1345 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111000; // iC= 2104 
// vC = 14'b1111101101001101; // vC=-1203 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111111; // iC= 1983 
// vC = 14'b1111101101110100; // vC=-1164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001110; // iC= 2126 
// vC = 14'b1111101011010111; // vC=-1321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111110; // iC= 1982 
// vC = 14'b1111101010111110; // vC=-1346 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000101; // iC= 2117 
// vC = 14'b1111101011001100; // vC=-1332 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101011; // iC= 2155 
// vC = 14'b1111101111100001; // vC=-1055 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b1111101011110000; // vC=-1296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111101110110000; // vC=-1104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011100; // iC= 2140 
// vC = 14'b1111101011011000; // vC=-1320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b1111101101100110; // vC=-1178 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110011; // iC= 1971 
// vC = 14'b1111101111010011; // vC=-1069 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100011; // iC= 1891 
// vC = 14'b1111101011010111; // vC=-1321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010011; // iC= 2195 
// vC = 14'b1111101100101001; // vC=-1239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000011; // iC= 1923 
// vC = 14'b1111101111111100; // vC=-1028 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111101110101110; // vC=-1106 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b1111101110101101; // vC=-1107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b1111101110000101; // vC=-1147 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100101; // iC= 1957 
// vC = 14'b1111101101011111; // vC=-1185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010000; // iC= 2064 
// vC = 14'b1111110000001101; // vC=-1011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b1111101111011101; // vC=-1059 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011111; // iC= 2015 
// vC = 14'b1111110000010000; // vC=-1008 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b1111101101000100; // vC=-1212 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010111; // iC= 2199 
// vC = 14'b1111110000101000; // vC= -984 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b1111101111000001; // vC=-1087 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111011; // iC= 2107 
// vC = 14'b1111110001001101; // vC= -947 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111011; // iC= 2171 
// vC = 14'b1111110000011110; // vC= -994 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b1111101110001111; // vC=-1137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100101; // iC= 2149 
// vC = 14'b1111110010011101; // vC= -867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b1111110010101100; // vC= -852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001001; // iC= 2121 
// vC = 14'b1111101110110111; // vC=-1097 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b1111110000000001; // vC=-1023 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111001; // iC= 2169 
// vC = 14'b1111110010101001; // vC= -855 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b1111110001111011; // vC= -901 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111101110111000; // vC=-1096 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b1111110010001011; // vC= -885 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001101; // iC= 1997 
// vC = 14'b1111110000101011; // vC= -981 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000100; // iC= 2244 
// vC = 14'b1111110011111110; // vC= -770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111110011000111; // vC= -825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b1111110000100001; // vC= -991 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110010; // iC= 2226 
// vC = 14'b1111110001111010; // vC= -902 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000111; // iC= 2055 
// vC = 14'b1111110001011111; // vC= -929 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110110; // iC= 2038 
// vC = 14'b1111101111101011; // vC=-1045 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110001; // iC= 2033 
// vC = 14'b1111110000101100; // vC= -980 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b1111110000011000; // vC=-1000 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b1111110100101010; // vC= -726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001011; // iC= 1995 
// vC = 14'b1111110010100000; // vC= -864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010000; // iC= 2000 
// vC = 14'b1111110011000100; // vC= -828 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111110101011001; // vC= -679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101110; // iC= 1966 
// vC = 14'b1111110011000001; // vC= -831 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111101; // iC= 2237 
// vC = 14'b1111110100000001; // vC= -767 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101000; // iC= 2152 
// vC = 14'b1111110011011011; // vC= -805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000110; // iC= 2246 
// vC = 14'b1111110010000101; // vC= -891 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b1111110101010101; // vC= -683 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110011; // iC= 2227 
// vC = 14'b1111110001110010; // vC= -910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b1111110100011001; // vC= -743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b1111110100001100; // vC= -756 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111110100100000; // vC= -736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010101; // iC= 2197 
// vC = 14'b1111110111000001; // vC= -575 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100011; // iC= 2147 
// vC = 14'b1111110010001001; // vC= -887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b1111110101110001; // vC= -655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b1111110100100101; // vC= -731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001011; // iC= 2251 
// vC = 14'b1111110111100011; // vC= -541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110101; // iC= 2229 
// vC = 14'b1111110100101011; // vC= -725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011111; // iC= 2015 
// vC = 14'b1111110011000100; // vC= -828 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011011101; // iC= 2269 
// vC = 14'b1111110111001001; // vC= -567 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011100; // iC= 2076 
// vC = 14'b1111110100111100; // vC= -708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110000; // iC= 2160 
// vC = 14'b1111110100001110; // vC= -754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001000; // iC= 2120 
// vC = 14'b1111110011111011; // vC= -773 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011111; // iC= 2079 
// vC = 14'b1111110101111000; // vC= -648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001010; // iC= 2250 
// vC = 14'b1111110110101101; // vC= -595 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111110100011001; // vC= -743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000000; // iC= 2240 
// vC = 14'b1111110110110111; // vC= -585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010001; // iC= 2257 
// vC = 14'b1111110110000101; // vC= -635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b1111110101110111; // vC= -649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b1111110111101010; // vC= -534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111110100110110; // vC= -714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000101; // iC= 2245 
// vC = 14'b1111110110001100; // vC= -628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111100; // iC= 2108 
// vC = 14'b1111110101100011; // vC= -669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110011; // iC= 2099 
// vC = 14'b1111110111010011; // vC= -557 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000110; // iC= 2182 
// vC = 14'b1111110111111000; // vC= -520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111101; // iC= 2045 
// vC = 14'b1111111010000010; // vC= -382 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011000; // iC= 2136 
// vC = 14'b1111111000100101; // vC= -475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001001; // iC= 2121 
// vC = 14'b1111111010100000; // vC= -352 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101101; // iC= 2157 
// vC = 14'b1111111001001000; // vC= -440 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010001; // iC= 2257 
// vC = 14'b1111110111001101; // vC= -563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000001; // iC= 2177 
// vC = 14'b1111110111110010; // vC= -526 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111011; // iC= 2171 
// vC = 14'b1111111010111010; // vC= -326 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100000; // iC= 2144 
// vC = 14'b1111111011010010; // vC= -302 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b1111111001101001; // vC= -407 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111011; // iC= 2107 
// vC = 14'b1111111001000000; // vC= -448 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b1111111010010000; // vC= -368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010001; // iC= 2001 
// vC = 14'b1111111000100101; // vC= -475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b1111110111110101; // vC= -523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011000; // iC= 2072 
// vC = 14'b1111110111001101; // vC= -563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111001; // iC= 2105 
// vC = 14'b1111111001001010; // vC= -438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101011; // iC= 2155 
// vC = 14'b1111110111111100; // vC= -516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110100; // iC= 2228 
// vC = 14'b1111111100100101; // vC= -219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111110; // iC= 2046 
// vC = 14'b1111111100110011; // vC= -205 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b1111111011011000; // vC= -296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000001; // iC= 2241 
// vC = 14'b1111111011000111; // vC= -313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111111001111001; // vC= -391 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b1111111100111100; // vC= -196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111001; // iC= 2169 
// vC = 14'b1111111011001101; // vC= -307 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001101; // iC= 2253 
// vC = 14'b1111111010011011; // vC= -357 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011011001; // iC= 2265 
// vC = 14'b1111111101101001; // vC= -151 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110110; // iC= 2102 
// vC = 14'b1111111001100010; // vC= -414 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b1111111011010010; // vC= -302 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b1111111010100011; // vC= -349 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b1111111001100011; // vC= -413 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101100; // iC= 2220 
// vC = 14'b1111111101101111; // vC= -145 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b1111111010100100; // vC= -348 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111110; // iC= 2110 
// vC = 14'b1111111100100011; // vC= -221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000010; // iC= 2178 
// vC = 14'b1111111101011111; // vC= -161 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100000; // iC= 2144 
// vC = 14'b1111111100100100; // vC= -220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001110; // iC= 2254 
// vC = 14'b1111111100111111; // vC= -193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111111101110110; // vC= -138 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010010; // iC= 2258 
// vC = 14'b1111111110101010; // vC=  -86 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111111011111100; // vC= -260 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110110; // iC= 2166 
// vC = 14'b1111111010110010; // vC= -334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101000; // iC= 2024 
// vC = 14'b1111111100111111; // vC= -193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000010; // iC= 1986 
// vC = 14'b1111111100101101; // vC= -211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111111100001110; // vC= -242 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100100; // iC= 2212 
// vC = 14'b1111111011110111; // vC= -265 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b1111111110110111; // vC=  -73 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b1111111100101011; // vC= -213 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111010; // iC= 2106 
// vC = 14'b1111111110111000; // vC=  -72 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b1111111100011010; // vC= -230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b1111111100000000; // vC= -256 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001100; // iC= 2252 
// vC = 14'b0000000000010100; // vC=   20 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001111; // iC= 2191 
// vC = 14'b0000000000111110; // vC=   62 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b1111111110111101; // vC=  -67 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111110; // iC= 2046 
// vC = 14'b1111111111010011; // vC=  -45 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b1111111110011010; // vC= -102 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b0000000000000111; // vC=    7 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b0000000001101000; // vC=  104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110110; // iC= 2230 
// vC = 14'b1111111110001011; // vC= -117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111111; // iC= 2175 
// vC = 14'b1111111101010111; // vC= -169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110101; // iC= 2101 
// vC = 14'b0000000001011111; // vC=   95 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b0000000001100011; // vC=   99 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001101; // iC= 2189 
// vC = 14'b0000000010011111; // vC=  159 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001000; // iC= 2120 
// vC = 14'b0000000010101011; // vC=  171 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b0000000001111110; // vC=  126 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001110; // iC= 1934 
// vC = 14'b0000000000011010; // vC=   26 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111111111000110; // vC=  -58 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011100; // iC= 2140 
// vC = 14'b1111111110110111; // vC=  -73 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110000; // iC= 2224 
// vC = 14'b0000000010000110; // vC=  134 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100100; // iC= 2148 
// vC = 14'b0000000001010111; // vC=   87 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b0000000001101110; // vC=  110 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b1111111111001101; // vC=  -51 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b0000000010101000; // vC=  168 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b0000000001000010; // vC=   66 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011011; // iC= 2203 
// vC = 14'b1111111111110010; // vC=  -14 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110110; // iC= 2038 
// vC = 14'b1111111111101000; // vC=  -24 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010011; // iC= 2131 
// vC = 14'b0000000100100001; // vC=  289 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101011; // iC= 2155 
// vC = 14'b0000000000101101; // vC=   45 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101001; // iC= 2153 
// vC = 14'b0000000000010111; // vC=   23 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b0000000000001011; // vC=   11 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010000; // iC= 2000 
// vC = 14'b0000000001010101; // vC=   85 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011110; // iC= 2078 
// vC = 14'b0000000101010100; // vC=  340 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001110; // iC= 2126 
// vC = 14'b0000000011011111; // vC=  223 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b0000000100110011; // vC=  307 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b0000000011011001; // vC=  217 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101110; // iC= 2030 
// vC = 14'b0000000001010101; // vC=   85 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010010; // iC= 2002 
// vC = 14'b0000000101010100; // vC=  340 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110101; // iC= 1909 
// vC = 14'b0000000011010100; // vC=  212 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b0000000001101011; // vC=  107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b0000000010011011; // vC=  155 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011100; // iC= 2012 
// vC = 14'b0000000001101001; // vC=  105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101110; // iC= 2158 
// vC = 14'b0000000110010101; // vC=  405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011100; // iC= 2076 
// vC = 14'b0000000101100100; // vC=  356 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001011; // iC= 1867 
// vC = 14'b0000000101011101; // vC=  349 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100100; // iC= 1892 
// vC = 14'b0000000100001111; // vC=  271 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011010; // iC= 1882 
// vC = 14'b0000000011110111; // vC=  247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011100; // iC= 2076 
// vC = 14'b0000000110100010; // vC=  418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b0000000010111000; // vC=  184 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b0000000111001000; // vC=  456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b0000000110101100; // vC=  428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110010; // iC= 2034 
// vC = 14'b0000000100010001; // vC=  273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100110; // iC= 2086 
// vC = 14'b0000000100010100; // vC=  276 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b0000001000001110; // vC=  526 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000001; // iC= 1921 
// vC = 14'b0000000111111110; // vC=  510 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100100; // iC= 2148 
// vC = 14'b0000000100000010; // vC=  258 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b0000000101011111; // vC=  351 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b0000000110100111; // vC=  423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b0000000110010101; // vC=  405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b0000001000010101; // vC=  533 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101101; // iC= 1901 
// vC = 14'b0000000111001001; // vC=  457 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101111; // iC= 2095 
// vC = 14'b0000000110001010; // vC=  394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b0000000110100001; // vC=  417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b0000000111110010; // vC=  498 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b0000001000100110; // vC=  550 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b0000000111100011; // vC=  483 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001011; // iC= 1995 
// vC = 14'b0000000111110001; // vC=  497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b0000000111101000; // vC=  488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001101; // iC= 2125 
// vC = 14'b0000000110011110; // vC=  414 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b0000001010001000; // vC=  648 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b0000001001011000; // vC=  600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001100; // iC= 1868 
// vC = 14'b0000000111011000; // vC=  472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b0000001001101010; // vC=  618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011001; // iC= 1817 
// vC = 14'b0000000111100111; // vC=  487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b0000001001000000; // vC=  576 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110101; // iC= 1909 
// vC = 14'b0000000111011011; // vC=  475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b0000001001000101; // vC=  581 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111000; // iC= 1912 
// vC = 14'b0000001001110111; // vC=  631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b0000001011010010; // vC=  722 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b0000001001000000; // vC=  576 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111100; // iC= 1916 
// vC = 14'b0000001001011000; // vC=  600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110110; // iC= 1910 
// vC = 14'b0000001011001111; // vC=  719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000101; // iC= 1861 
// vC = 14'b0000001011000001; // vC=  705 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001000; // iC= 1864 
// vC = 14'b0000000111100111; // vC=  487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010110; // iC= 2070 
// vC = 14'b0000001000011010; // vC=  538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000101; // iC= 2053 
// vC = 14'b0000000111011101; // vC=  477 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001011; // iC= 1995 
// vC = 14'b0000001010000111; // vC=  647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b0000001000000101; // vC=  517 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101111; // iC= 1967 
// vC = 14'b0000001001110001; // vC=  625 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b0000001001101111; // vC=  623 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100010; // iC= 1890 
// vC = 14'b0000001000100010; // vC=  546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b0000001011100000; // vC=  736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100010; // iC= 1762 
// vC = 14'b0000001101000111; // vC=  839 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001111; // iC= 1807 
// vC = 14'b0000001011111100; // vC=  764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010011; // iC= 1747 
// vC = 14'b0000001010000001; // vC=  641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011000; // iC= 1752 
// vC = 14'b0000001010000111; // vC=  647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000011; // iC= 1731 
// vC = 14'b0000001010101111; // vC=  687 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b0000001011001111; // vC=  719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000001; // iC= 1921 
// vC = 14'b0000001001010011; // vC=  595 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b0000001011101101; // vC=  749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b0000001011101000; // vC=  744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110101; // iC= 1717 
// vC = 14'b0000001011000111; // vC=  711 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001000; // iC= 1928 
// vC = 14'b0000001100111101; // vC=  829 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111010; // iC= 1786 
// vC = 14'b0000001100010101; // vC=  789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000110; // iC= 1862 
// vC = 14'b0000001011110010; // vC=  754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010111; // iC= 1815 
// vC = 14'b0000001110011100; // vC=  924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010000; // iC= 2000 
// vC = 14'b0000001010101001; // vC=  681 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000001; // iC= 1857 
// vC = 14'b0000001010101101; // vC=  685 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100111; // iC= 1767 
// vC = 14'b0000001100100010; // vC=  802 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110100; // iC= 1716 
// vC = 14'b0000001101010001; // vC=  849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b0000001111001011; // vC=  971 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b0000001110110111; // vC=  951 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001011; // iC= 1739 
// vC = 14'b0000001011010000; // vC=  720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011011; // iC= 1819 
// vC = 14'b0000001101110111; // vC=  887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100011; // iC= 1699 
// vC = 14'b0000001101101101; // vC=  877 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b0000001100010101; // vC=  789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000000; // iC= 1728 
// vC = 14'b0000001101000011; // vC=  835 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010000; // iC= 1744 
// vC = 14'b0000001011111010; // vC=  762 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101101; // iC= 1837 
// vC = 14'b0000001110011100; // vC=  924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111100; // iC= 1916 
// vC = 14'b0000001100000011; // vC=  771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b0000001110101110; // vC=  942 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000100; // iC= 1668 
// vC = 14'b0000010000000011; // vC= 1027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b0000001100100001; // vC=  801 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b0000001111111010; // vC= 1018 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100000; // iC= 1696 
// vC = 14'b0000001110100101; // vC=  933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111110; // iC= 1726 
// vC = 14'b0000001100101000; // vC=  808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111011; // iC= 1915 
// vC = 14'b0000001101101100; // vC=  876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000000; // iC= 1856 
// vC = 14'b0000010000010100; // vC= 1044 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011101; // iC= 1821 
// vC = 14'b0000001110010010; // vC=  914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010000; // iC= 1616 
// vC = 14'b0000010000110001; // vC= 1073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110100; // iC= 1844 
// vC = 14'b0000010000001011; // vC= 1035 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001110; // iC= 1870 
// vC = 14'b0000010000110011; // vC= 1075 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b0000001110011101; // vC=  925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011110; // iC= 1630 
// vC = 14'b0000001101111010; // vC=  890 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000000; // iC= 1728 
// vC = 14'b0000001110110011; // vC=  947 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001011; // iC= 1739 
// vC = 14'b0000010010011000; // vC= 1176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011111; // iC= 1631 
// vC = 14'b0000001111110000; // vC= 1008 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101100; // iC= 1644 
// vC = 14'b0000001111110101; // vC= 1013 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111110; // iC= 1726 
// vC = 14'b0000001111000001; // vC=  961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010100; // iC= 1876 
// vC = 14'b0000001110010101; // vC=  917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110010; // iC= 1650 
// vC = 14'b0000010001111010; // vC= 1146 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010110; // iC= 1878 
// vC = 14'b0000010010001111; // vC= 1167 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101111; // iC= 1583 
// vC = 14'b0000001110010110; // vC=  918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110100; // iC= 1780 
// vC = 14'b0000010001101111; // vC= 1135 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111011; // iC= 1595 
// vC = 14'b0000010010101011; // vC= 1195 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110000; // iC= 1648 
// vC = 14'b0000010010010000; // vC= 1168 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011100; // iC= 1628 
// vC = 14'b0000010010111111; // vC= 1215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010101; // iC= 1685 
// vC = 14'b0000001111011101; // vC=  989 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110101; // iC= 1717 
// vC = 14'b0000001111101110; // vC= 1006 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101100; // iC= 1708 
// vC = 14'b0000010011001011; // vC= 1227 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110010; // iC= 1778 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110110; // iC= 1526 
// vC = 14'b0000010000011001; // vC= 1049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011000; // iC= 1624 
// vC = 14'b0000010011001111; // vC= 1231 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010100; // iC= 1620 
// vC = 14'b0000010001110101; // vC= 1141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100000; // iC= 1504 
// vC = 14'b0000010011000110; // vC= 1222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011010; // iC= 1498 
// vC = 14'b0000010100010001; // vC= 1297 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011011; // iC= 1691 
// vC = 14'b0000010011101111; // vC= 1263 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101110; // iC= 1582 
// vC = 14'b0000010010000110; // vC= 1158 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010001; // iC= 1553 
// vC = 14'b0000010100111010; // vC= 1338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011111; // iC= 1503 
// vC = 14'b0000010010010011; // vC= 1171 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110001; // iC= 1777 
// vC = 14'b0000010000010000; // vC= 1040 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011101; // iC= 1629 
// vC = 14'b0000010000111101; // vC= 1085 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110111; // iC= 1527 
// vC = 14'b0000010100100111; // vC= 1319 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011101; // iC= 1501 
// vC = 14'b0000010011011000; // vC= 1240 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010001; // iC= 1489 
// vC = 14'b0000010001010100; // vC= 1108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011000; // iC= 1752 
// vC = 14'b0000010010101001; // vC= 1193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000011; // iC= 1667 
// vC = 14'b0000010010110010; // vC= 1202 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101000; // iC= 1704 
// vC = 14'b0000010101110101; // vC= 1397 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001010; // iC= 1482 
// vC = 14'b0000010101011011; // vC= 1371 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110011; // iC= 1651 
// vC = 14'b0000010101100111; // vC= 1383 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001001; // iC= 1737 
// vC = 14'b0000010110010011; // vC= 1427 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010110; // iC= 1494 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010111; // iC= 1495 
// vC = 14'b0000010011000001; // vC= 1217 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100110; // iC= 1638 
// vC = 14'b0000010001100000; // vC= 1120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010001; // iC= 1553 
// vC = 14'b0000010011100001; // vC= 1249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011100; // iC= 1628 
// vC = 14'b0000010100101111; // vC= 1327 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110000; // iC= 1712 
// vC = 14'b0000010011000010; // vC= 1218 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001110; // iC= 1550 
// vC = 14'b0000010110000110; // vC= 1414 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011000; // iC= 1624 
// vC = 14'b0000010101001111; // vC= 1359 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001110; // iC= 1550 
// vC = 14'b0000010110010100; // vC= 1428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101010; // iC= 1514 
// vC = 14'b0000010011011001; // vC= 1241 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101101; // iC= 1645 
// vC = 14'b0000010100001000; // vC= 1288 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110000; // iC= 1648 
// vC = 14'b0000010010110000; // vC= 1200 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b0000010100110011; // vC= 1331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100111; // iC= 1639 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010010; // iC= 1490 
// vC = 14'b0000010101111110; // vC= 1406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101111; // iC= 1519 
// vC = 14'b0000010101111011; // vC= 1403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111110; // iC= 1342 
// vC = 14'b0000010100001011; // vC= 1291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000111; // iC= 1607 
// vC = 14'b0000010011011111; // vC= 1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001101; // iC= 1485 
// vC = 14'b0000010110000100; // vC= 1412 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101101; // iC= 1453 
// vC = 14'b0000010100011111; // vC= 1311 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100111; // iC= 1447 
// vC = 14'b0000010100001011; // vC= 1291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000011; // iC= 1539 
// vC = 14'b0000010111000101; // vC= 1477 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110100; // iC= 1332 
// vC = 14'b0000010100010111; // vC= 1303 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000111; // iC= 1415 
// vC = 14'b0000010101111011; // vC= 1403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110100; // iC= 1460 
// vC = 14'b0000010100101001; // vC= 1321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111010; // iC= 1338 
// vC = 14'b0000011000001100; // vC= 1548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101110; // iC= 1518 
// vC = 14'b0000010101111010; // vC= 1402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100111; // iC= 1383 
// vC = 14'b0000011000011110; // vC= 1566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000011; // iC= 1283 
// vC = 14'b0000010110001010; // vC= 1418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100111; // iC= 1511 
// vC = 14'b0000010101100111; // vC= 1383 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001110; // iC= 1550 
// vC = 14'b0000010111000110; // vC= 1478 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101000; // iC= 1576 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111000; // iC= 1400 
// vC = 14'b0000010111011101; // vC= 1501 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010000; // iC= 1552 
// vC = 14'b0000011000010000; // vC= 1552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110100; // iC= 1396 
// vC = 14'b0000010101001010; // vC= 1354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110111; // iC= 1463 
// vC = 14'b0000010101101010; // vC= 1386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100001; // iC= 1441 
// vC = 14'b0000010111110111; // vC= 1527 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101000; // iC= 1512 
// vC = 14'b0000010110100011; // vC= 1443 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101010; // iC= 1322 
// vC = 14'b0000011001111010; // vC= 1658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101101; // iC= 1389 
// vC = 14'b0000010111000111; // vC= 1479 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000101; // iC= 1413 
// vC = 14'b0000010111010011; // vC= 1491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000111; // iC= 1351 
// vC = 14'b0000011000010001; // vC= 1553 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100101; // iC= 1381 
// vC = 14'b0000010110100110; // vC= 1446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101111; // iC= 1455 
// vC = 14'b0000010110111111; // vC= 1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010101; // iC= 1493 
// vC = 14'b0000011000100000; // vC= 1568 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111000; // iC= 1208 
// vC = 14'b0000011010000101; // vC= 1669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101001; // iC= 1385 
// vC = 14'b0000010101111110; // vC= 1406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001100; // iC= 1484 
// vC = 14'b0000011001011000; // vC= 1624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101101; // iC= 1197 
// vC = 14'b0000010111011001; // vC= 1497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110000; // iC= 1200 
// vC = 14'b0000010101111110; // vC= 1406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001010; // iC= 1418 
// vC = 14'b0000010110100111; // vC= 1447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101101; // iC= 1453 
// vC = 14'b0000011010000101; // vC= 1669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011110; // iC= 1182 
// vC = 14'b0000011000000010; // vC= 1538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000010; // iC= 1346 
// vC = 14'b0000010111111100; // vC= 1532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100101; // iC= 1317 
// vC = 14'b0000011000111001; // vC= 1593 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101100; // iC= 1196 
// vC = 14'b0000010110100100; // vC= 1444 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001011; // iC= 1419 
// vC = 14'b0000010111110000; // vC= 1520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010111; // iC= 1175 
// vC = 14'b0000011011001110; // vC= 1742 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101000; // iC= 1320 
// vC = 14'b0000010111110110; // vC= 1526 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110000; // iC= 1200 
// vC = 14'b0000011001100001; // vC= 1633 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100010; // iC= 1186 
// vC = 14'b0000011001111011; // vC= 1659 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111001; // iC= 1209 
// vC = 14'b0000011000000011; // vC= 1539 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010000; // iC= 1360 
// vC = 14'b0000011000111111; // vC= 1599 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110000; // iC= 1392 
// vC = 14'b0000010111100101; // vC= 1509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011101; // iC= 1373 
// vC = 14'b0000011001001111; // vC= 1615 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110011; // iC= 1139 
// vC = 14'b0000011011011011; // vC= 1755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100011; // iC= 1123 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101010; // iC= 1386 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010000; // iC= 1104 
// vC = 14'b0000011001000101; // vC= 1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011110; // iC= 1374 
// vC = 14'b0000011010110101; // vC= 1717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001011; // iC= 1291 
// vC = 14'b0000011100100100; // vC= 1828 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001100; // iC= 1228 
// vC = 14'b0000011001101101; // vC= 1645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000110; // iC= 1286 
// vC = 14'b0000011010011111; // vC= 1695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000010; // iC= 1282 
// vC = 14'b0000011001110110; // vC= 1654 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010100; // iC= 1044 
// vC = 14'b0000011100110111; // vC= 1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011100; // iC= 1180 
// vC = 14'b0000011100011010; // vC= 1818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001011; // iC= 1227 
// vC = 14'b0000011011001101; // vC= 1741 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101110; // iC= 1198 
// vC = 14'b0000011001110010; // vC= 1650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101110; // iC= 1134 
// vC = 14'b0000011100101001; // vC= 1833 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110111; // iC= 1207 
// vC = 14'b0000011001111000; // vC= 1656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011101; // iC= 1309 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011101; // iC=  989 
// vC = 14'b0000011101100001; // vC= 1889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001100; // iC= 1164 
// vC = 14'b0000011010011110; // vC= 1694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001011; // iC= 1035 
// vC = 14'b0000011010100001; // vC= 1697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100100; // iC= 1060 
// vC = 14'b0000011011101101; // vC= 1773 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110010; // iC= 1138 
// vC = 14'b0000011010100000; // vC= 1696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011100; // iC= 1244 
// vC = 14'b0000011010011111; // vC= 1695 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011011; // iC=  987 
// vC = 14'b0000011001011011; // vC= 1627 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100111; // iC= 1127 
// vC = 14'b0000011011001010; // vC= 1738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101011; // iC= 1195 
// vC = 14'b0000011101001101; // vC= 1869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100001; // iC= 1249 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011001; // iC=  985 
// vC = 14'b0000011010100110; // vC= 1702 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110110; // iC= 1014 
// vC = 14'b0000011100101010; // vC= 1834 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110100; // iC= 1076 
// vC = 14'b0000011010101010; // vC= 1706 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100101; // iC= 1125 
// vC = 14'b0000011010001001; // vC= 1673 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001000; // iC=  904 
// vC = 14'b0000011011110100; // vC= 1780 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011111; // iC= 1119 
// vC = 14'b0000011011011011; // vC= 1755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000000; // iC= 1088 
// vC = 14'b0000011010101110; // vC= 1710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011111; // iC=  991 
// vC = 14'b0000011010000010; // vC= 1666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001001; // iC= 1097 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000111; // iC= 1031 
// vC = 14'b0000011101011111; // vC= 1887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001111; // iC=  975 
// vC = 14'b0000011010101110; // vC= 1710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011011; // iC= 1179 
// vC = 14'b0000011101011001; // vC= 1881 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000111; // iC= 1095 
// vC = 14'b0000011100111100; // vC= 1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001000; // iC= 1032 
// vC = 14'b0000011010001010; // vC= 1674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110000; // iC= 1136 
// vC = 14'b0000011101001000; // vC= 1864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100010; // iC=  866 
// vC = 14'b0000011101000010; // vC= 1858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100001; // iC=  929 
// vC = 14'b0000011101010001; // vC= 1873 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000000; // iC=  960 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011100; // iC=  860 
// vC = 14'b0000011100100001; // vC= 1825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001001; // iC= 1097 
// vC = 14'b0000011110010111; // vC= 1943 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101010; // iC=  874 
// vC = 14'b0000011100111111; // vC= 1855 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010100; // iC= 1044 
// vC = 14'b0000011011010100; // vC= 1748 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100111; // iC=  807 
// vC = 14'b0000011100101011; // vC= 1835 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111111; // iC=  959 
// vC = 14'b0000011011110010; // vC= 1778 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110001; // iC=  945 
// vC = 14'b0000011101001001; // vC= 1865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000100; // iC=  900 
// vC = 14'b0000011101011010; // vC= 1882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111110; // iC=  830 
// vC = 14'b0000011111101110; // vC= 2030 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011101; // iC=  797 
// vC = 14'b0000011111110010; // vC= 2034 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110000; // iC=  880 
// vC = 14'b0000011110100110; // vC= 1958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010010; // iC=  914 
// vC = 14'b0000011011101101; // vC= 1773 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000010; // iC=  962 
// vC = 14'b0000011100100110; // vC= 1830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011001; // iC=  793 
// vC = 14'b0000011011110101; // vC= 1781 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000010; // iC=  834 
// vC = 14'b0000011111100111; // vC= 2023 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110110; // iC=  822 
// vC = 14'b0000011011111001; // vC= 1785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100100; // iC=  932 
// vC = 14'b0000100000000110; // vC= 2054 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101011; // iC=  939 
// vC = 14'b0000011110000100; // vC= 1924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010101; // iC=  917 
// vC = 14'b0000011111011101; // vC= 2013 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110101; // iC=  821 
// vC = 14'b0000011101110000; // vC= 1904 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001100; // iC=  716 
// vC = 14'b0000011110001001; // vC= 1929 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011100; // iC=  796 
// vC = 14'b0000011100111011; // vC= 1851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011101; // iC=  925 
// vC = 14'b0000100000100010; // vC= 2082 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010110; // iC=  854 
// vC = 14'b0000011101111110; // vC= 1918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110100; // iC=  692 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101010; // iC=  810 
// vC = 14'b0000100000011011; // vC= 2075 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001100; // iC=  716 
// vC = 14'b0000011100110001; // vC= 1841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110000; // iC=  816 
// vC = 14'b0000011111101000; // vC= 2024 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001111; // iC=  719 
// vC = 14'b0000100000010101; // vC= 2069 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000110; // iC=  646 
// vC = 14'b0000100000111011; // vC= 2107 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111001; // iC=  761 
// vC = 14'b0000011111101001; // vC= 2025 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101011; // iC=  811 
// vC = 14'b0000011101011111; // vC= 1887 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101000; // iC=  808 
// vC = 14'b0000011100110110; // vC= 1846 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000110; // iC=  774 
// vC = 14'b0000011100111010; // vC= 1850 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000101; // iC=  773 
// vC = 14'b0000100000010101; // vC= 2069 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010011; // iC=  723 
// vC = 14'b0000011111011010; // vC= 2010 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001111; // iC=  591 
// vC = 14'b0000011111111111; // vC= 2047 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100000; // iC=  736 
// vC = 14'b0000100000001000; // vC= 2056 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100101; // iC=  741 
// vC = 14'b0000011110010010; // vC= 1938 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010111; // iC=  727 
// vC = 14'b0000011110110110; // vC= 1974 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111011; // iC=  763 
// vC = 14'b0000100001000111; // vC= 2119 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101000; // iC=  872 
// vC = 14'b0000011101001111; // vC= 1871 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001101; // iC=  589 
// vC = 14'b0000100001011100; // vC= 2140 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011100; // iC=  604 
// vC = 14'b0000011110001100; // vC= 1932 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101000; // iC=  744 
// vC = 14'b0000100001010101; // vC= 2133 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101010; // iC=  618 
// vC = 14'b0000011110100110; // vC= 1958 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011111; // iC=  607 
// vC = 14'b0000011101111010; // vC= 1914 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001101; // iC=  781 
// vC = 14'b0000100000001011; // vC= 2059 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100000; // iC=  608 
// vC = 14'b0000011110011010; // vC= 1946 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110011; // iC=  755 
// vC = 14'b0000100001001111; // vC= 2127 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100110; // iC=  550 
// vC = 14'b0000011111100011; // vC= 2019 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100100; // iC=  740 
// vC = 14'b0000011100110011; // vC= 1843 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111010; // iC=  570 
// vC = 14'b0000011111111100; // vC= 2044 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101110; // iC=  750 
// vC = 14'b0000011111101011; // vC= 2027 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001011; // iC=  523 
// vC = 14'b0000011111011100; // vC= 2012 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101110; // iC=  686 
// vC = 14'b0000011111101000; // vC= 2024 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001101; // iC=  397 
// vC = 14'b0000011111111001; // vC= 2041 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110011; // iC=  499 
// vC = 14'b0000011110101010; // vC= 1962 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110110; // iC=  630 
// vC = 14'b0000100000111111; // vC= 2111 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001100; // iC=  524 
// vC = 14'b0000100001010001; // vC= 2129 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011111; // iC=  351 
// vC = 14'b0000100010001000; // vC= 2184 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111110; // iC=  446 
// vC = 14'b0000011101011011; // vC= 1883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101111; // iC=  431 
// vC = 14'b0000100000000111; // vC= 2055 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011011; // iC=  411 
// vC = 14'b0000100001000111; // vC= 2119 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111001; // iC=  505 
// vC = 14'b0000100001100001; // vC= 2145 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010001; // iC=  401 
// vC = 14'b0000011111111011; // vC= 2043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101001; // iC=  553 
// vC = 14'b0000100000101101; // vC= 2093 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101001; // iC=  553 
// vC = 14'b0000011101110010; // vC= 1906 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010110; // iC=  278 
// vC = 14'b0000100000001101; // vC= 2061 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110110; // iC=  246 
// vC = 14'b0000100001100011; // vC= 2147 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011010; // iC=  346 
// vC = 14'b0000011101101100; // vC= 1900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010011; // iC=  339 
// vC = 14'b0000011110001010; // vC= 1930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010011; // iC=  339 
// vC = 14'b0000100001110111; // vC= 2167 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111010; // iC=  378 
// vC = 14'b0000011110011100; // vC= 1948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010111; // iC=  407 
// vC = 14'b0000100000011001; // vC= 2073 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100100; // iC=  164 
// vC = 14'b0000011111010011; // vC= 2003 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000111; // iC=  391 
// vC = 14'b0000100010001011; // vC= 2187 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111100; // iC=  316 
// vC = 14'b0000100010011000; // vC= 2200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000111; // iC=  327 
// vC = 14'b0000011111011110; // vC= 2014 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001001; // iC=  137 
// vC = 14'b0000100001101010; // vC= 2154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010101; // iC=   21 
// vC = 14'b0000100001000011; // vC= 2115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101010; // iC=  106 
// vC = 14'b0000100000010000; // vC= 2064 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101100; // iC=  300 
// vC = 14'b0000011110110011; // vC= 1971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110110; // iC=  246 
// vC = 14'b0000100010010000; // vC= 2192 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001000100; // iC=   68 
// vC = 14'b0000011110101111; // vC= 1967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000101; // iC=  -59 
// vC = 14'b0000100001000001; // vC= 2113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010100; // iC=  148 
// vC = 14'b0000100000110001; // vC= 2097 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111111; // iC=  191 
// vC = 14'b0000100001010011; // vC= 2131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001101; // iC=   77 
// vC = 14'b0000100001001101; // vC= 2125 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100001; // iC=   33 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011101; // iC=   29 
// vC = 14'b0000011110011111; // vC= 1951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001001; // iC=  -55 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101111; // iC=   47 
// vC = 14'b0000100001100000; // vC= 2144 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100000; // iC=   32 
// vC = 14'b0000100001000001; // vC= 2113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000110; // iC= -186 
// vC = 14'b0000100001111100; // vC= 2172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010011; // iC=  -45 
// vC = 14'b0000100010010110; // vC= 2198 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110101110; // iC=  -82 
// vC = 14'b0000011101111011; // vC= 1915 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110111; // iC= -201 
// vC = 14'b0000011110011011; // vC= 1947 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000101; // iC= -379 
// vC = 14'b0000100001100101; // vC= 2149 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111111; // iC= -193 
// vC = 14'b0000011111101111; // vC= 2031 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100101; // iC= -155 
// vC = 14'b0000011101111101; // vC= 1917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110111; // iC= -201 
// vC = 14'b0000100001001001; // vC= 2121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101000; // iC= -472 
// vC = 14'b0000011101011111; // vC= 1887 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001011; // iC= -501 
// vC = 14'b0000011101101110; // vC= 1902 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111110010; // iC= -526 
// vC = 14'b0000100001101000; // vC= 2152 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110111; // iC= -457 
// vC = 14'b0000011110110011; // vC= 1971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001100; // iC= -436 
// vC = 14'b0000011111010100; // vC= 2004 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001101; // iC= -499 
// vC = 14'b0000100010000011; // vC= 2179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111100; // iC= -388 
// vC = 14'b0000011110101001; // vC= 1961 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110100; // iC= -652 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111001; // iC= -583 
// vC = 14'b0000011101000001; // vC= 1857 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000110; // iC= -378 
// vC = 14'b0000011111010001; // vC= 2001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011000; // iC= -424 
// vC = 14'b0000100000010001; // vC= 2065 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101100; // iC= -468 
// vC = 14'b0000100001001111; // vC= 2127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100100; // iC= -540 
// vC = 14'b0000011101101001; // vC= 1897 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000101; // iC= -763 
// vC = 14'b0000100001000011; // vC= 2115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100101; // iC= -667 
// vC = 14'b0000100001001100; // vC= 2124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001100; // iC= -692 
// vC = 14'b0000011101110111; // vC= 1911 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100100; // iC= -860 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010001; // iC= -815 
// vC = 14'b0000100000000011; // vC= 2051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101000; // iC= -600 
// vC = 14'b0000011110110000; // vC= 1968 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000111; // iC= -633 
// vC = 14'b0000100000010110; // vC= 2070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110100; // iC= -716 
// vC = 14'b0000011111010000; // vC= 2000 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110011; // iC= -781 
// vC = 14'b0000100000110000; // vC= 2096 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101010; // iC= -982 
// vC = 14'b0000011100101000; // vC= 1832 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101101; // iC= -723 
// vC = 14'b0000100000000110; // vC= 2054 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111110; // iC= -770 
// vC = 14'b0000011100000110; // vC= 1798 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010110; // iC= -746 
// vC = 14'b0000011110110010; // vC= 1970 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010111; // iC= -809 
// vC = 14'b0000011100010011; // vC= 1811 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110111; // iC= -905 
// vC = 14'b0000100000110101; // vC= 2101 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100001; // iC= -927 
// vC = 14'b0000011100100110; // vC= 1830 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011011; // iC=-1125 
// vC = 14'b0000100000110001; // vC= 2097 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111001; // iC=-1095 
// vC = 14'b0000011011110111; // vC= 1783 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101001; // iC= -983 
// vC = 14'b0000011100100100; // vC= 1828 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001000; // iC=-1144 
// vC = 14'b0000011101000101; // vC= 1861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100010; // iC= -926 
// vC = 14'b0000100000011100; // vC= 2076 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111111; // iC=-1089 
// vC = 14'b0000011111011010; // vC= 2010 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101011; // iC=-1109 
// vC = 14'b0000011101000101; // vC= 1861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101101; // iC=-1171 
// vC = 14'b0000011100011001; // vC= 1817 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001011; // iC=-1077 
// vC = 14'b0000100000001110; // vC= 2062 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011111; // iC=-1313 
// vC = 14'b0000011101111011; // vC= 1915 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000011; // iC=-1341 
// vC = 14'b0000011101000111; // vC= 1863 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100100; // iC=-1244 
// vC = 14'b0000011111010001; // vC= 2001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111100; // iC=-1156 
// vC = 14'b0000011011011000; // vC= 1752 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110101; // iC=-1099 
// vC = 14'b0000011011101100; // vC= 1772 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010011; // iC=-1389 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000100; // iC=-1404 
// vC = 14'b0000011110110101; // vC= 1973 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010111; // iC=-1385 
// vC = 14'b0000011101110111; // vC= 1911 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010111; // iC=-1193 
// vC = 14'b0000011011111001; // vC= 1785 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011110; // iC=-1442 
// vC = 14'b0000011010010010; // vC= 1682 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101000; // iC=-1304 
// vC = 14'b0000011101011100; // vC= 1884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000100; // iC=-1404 
// vC = 14'b0000011100001000; // vC= 1800 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111011; // iC=-1349 
// vC = 14'b0000011100110010; // vC= 1842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001000; // iC=-1272 
// vC = 14'b0000011100010010; // vC= 1810 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010111; // iC=-1577 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010001; // iC=-1519 
// vC = 14'b0000011101101111; // vC= 1903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010000; // iC=-1584 
// vC = 14'b0000011110010111; // vC= 1943 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010100; // iC=-1580 
// vC = 14'b0000011011011100; // vC= 1756 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001001; // iC=-1463 
// vC = 14'b0000011100100100; // vC= 1828 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111110; // iC=-1474 
// vC = 14'b0000011100011111; // vC= 1823 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010011; // iC=-1453 
// vC = 14'b0000011010110110; // vC= 1718 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101000; // iC=-1624 
// vC = 14'b0000011101100100; // vC= 1892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101110; // iC=-1682 
// vC = 14'b0000011010111101; // vC= 1725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111111; // iC=-1601 
// vC = 14'b0000011100101001; // vC= 1833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100010; // iC=-1438 
// vC = 14'b0000011011001111; // vC= 1743 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011010; // iC=-1510 
// vC = 14'b0000011011111011; // vC= 1787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110010; // iC=-1486 
// vC = 14'b0000011010001101; // vC= 1677 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100001; // iC=-1759 
// vC = 14'b0000011000111011; // vC= 1595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000010; // iC=-1534 
// vC = 14'b0000011000110111; // vC= 1591 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010001; // iC=-1647 
// vC = 14'b0000011011110000; // vC= 1776 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010000; // iC=-1648 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001001; // iC=-1591 
// vC = 14'b0000011010000110; // vC= 1670 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000010; // iC=-1790 
// vC = 14'b0000011011100101; // vC= 1765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011110; // iC=-1826 
// vC = 14'b0000011000101001; // vC= 1577 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010101; // iC=-1707 
// vC = 14'b0000011011110111; // vC= 1783 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100101; // iC=-1691 
// vC = 14'b0000011010111010; // vC= 1722 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001011; // iC=-1589 
// vC = 14'b0000011001011100; // vC= 1628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001000; // iC=-1720 
// vC = 14'b0000011000100110; // vC= 1574 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b0000011001011110; // vC= 1630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000010111100100; // vC= 1508 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000011011100111; // vC= 1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010010; // iC=-1774 
// vC = 14'b0000011000010111; // vC= 1559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000011000101010; // vC= 1578 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001010; // iC=-1910 
// vC = 14'b0000011010000111; // vC= 1671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011011; // iC=-1829 
// vC = 14'b0000011001100100; // vC= 1636 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b0000010110100000; // vC= 1440 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b0000010111001101; // vC= 1485 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111111; // iC=-1985 
// vC = 14'b0000011010011000; // vC= 1688 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000100; // iC=-1788 
// vC = 14'b0000010110100100; // vC= 1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001111; // iC=-1841 
// vC = 14'b0000011000100011; // vC= 1571 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000111; // iC=-1977 
// vC = 14'b0000010111001111; // vC= 1487 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b0000010110100010; // vC= 1442 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010010; // iC=-1838 
// vC = 14'b0000011000110101; // vC= 1589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000011000110000; // vC= 1584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b0000010110100000; // vC= 1440 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000010110010001; // vC= 1425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b0000010101001010; // vC= 1354 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b0000010101001110; // vC= 1358 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000010101110000; // vC= 1392 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101010; // iC=-1814 
// vC = 14'b0000011000000100; // vC= 1540 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b0000010101000101; // vC= 1349 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000010110111010; // vC= 1466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b0000010101000010; // vC= 1346 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b0000010011110010; // vC= 1266 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110110; // iC=-2122 
// vC = 14'b0000010101100100; // vC= 1380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110111; // iC=-1865 
// vC = 14'b0000010110000001; // vC= 1409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b0000010011011010; // vC= 1242 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110100; // iC=-1932 
// vC = 14'b0000010111010110; // vC= 1494 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b0000010110011010; // vC= 1434 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b0000010100111010; // vC= 1338 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000110; // iC=-2170 
// vC = 14'b0000010110000010; // vC= 1410 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010101; // iC=-1899 
// vC = 14'b0000010111000001; // vC= 1473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b0000010110100101; // vC= 1445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000010110011101; // vC= 1437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010010; // iC=-2094 
// vC = 14'b0000010100110111; // vC= 1335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001101; // iC=-2163 
// vC = 14'b0000010010111001; // vC= 1209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b0000010011000101; // vC= 1221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011100; // iC=-1956 
// vC = 14'b0000010101110000; // vC= 1392 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b0000010001100110; // vC= 1126 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000010011000111; // vC= 1223 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b0000010010000001; // vC= 1153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b0000010000110110; // vC= 1078 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b0000010011110010; // vC= 1266 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101111; // iC=-2001 
// vC = 14'b0000010001011111; // vC= 1119 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011111; // iC=-2209 
// vC = 14'b0000010000110001; // vC= 1073 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000100; // iC=-2108 
// vC = 14'b0000010010001111; // vC= 1167 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011100; // iC=-1956 
// vC = 14'b0000010010100001; // vC= 1185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000001111111110; // vC= 1022 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111110; // iC=-2050 
// vC = 14'b0000010011101100; // vC= 1260 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001011; // iC=-2165 
// vC = 14'b0000010010111000; // vC= 1208 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000101; // iC=-2171 
// vC = 14'b0000010010000110; // vC= 1158 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001101; // iC=-2035 
// vC = 14'b0000010011100010; // vC= 1250 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b0000010010000110; // vC= 1158 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b0000001111001100; // vC=  972 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100001; // iC=-2207 
// vC = 14'b0000001111100110; // vC=  998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100110; // iC=-2138 
// vC = 14'b0000010011110010; // vC= 1266 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100100; // iC=-1948 
// vC = 14'b0000010001101011; // vC= 1131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111111; // iC=-1921 
// vC = 14'b0000010010100110; // vC= 1190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010001; // iC=-2031 
// vC = 14'b0000001111110000; // vC= 1008 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000111; // iC=-2105 
// vC = 14'b0000010010100000; // vC= 1184 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010101; // iC=-2155 
// vC = 14'b0000010000101010; // vC= 1066 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100111; // iC=-1945 
// vC = 14'b0000010000001101; // vC= 1037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111000; // iC=-1928 
// vC = 14'b0000001111000000; // vC=  960 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011100; // iC=-1956 
// vC = 14'b0000010000111000; // vC= 1080 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b0000001110110100; // vC=  948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000010000101110; // vC= 1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000010000101110; // vC= 1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110110; // iC=-1994 
// vC = 14'b0000010000110101; // vC= 1077 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000010000000001; // vC= 1025 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b0000001111101000; // vC= 1000 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011000; // iC=-2152 
// vC = 14'b0000001101010010; // vC=  850 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000001110011001; // vC=  921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111101; // iC=-2179 
// vC = 14'b0000001110111001; // vC=  953 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000001110001001; // vC=  905 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010000; // iC=-1968 
// vC = 14'b0000001110100111; // vC=  935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111111; // iC=-1985 
// vC = 14'b0000001101110010; // vC=  882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111110; // iC=-2242 
// vC = 14'b0000001110100001; // vC=  929 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b0000010000001011; // vC= 1035 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b0000001011100100; // vC=  740 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b0000001100000000; // vC=  768 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110010; // iC=-2254 
// vC = 14'b0000001100100010; // vC=  802 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000001111111011; // vC= 1019 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100011; // iC=-1949 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101000; // iC=-2264 
// vC = 14'b0000001100001111; // vC=  783 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000001; // iC=-2239 
// vC = 14'b0000001100010111; // vC=  791 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000001111000011; // vC=  963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100001; // iC=-2079 
// vC = 14'b0000001101101010; // vC=  874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100110; // iC=-2202 
// vC = 14'b0000001110010000; // vC=  912 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001101; // iC=-2227 
// vC = 14'b0000001101000001; // vC=  833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110000; // iC=-2064 
// vC = 14'b0000001010001011; // vC=  651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010100; // iC=-2092 
// vC = 14'b0000001101011101; // vC=  861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111000; // iC=-2120 
// vC = 14'b0000001100100001; // vC=  801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b0000001010100111; // vC=  679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b0000001001110011; // vC=  627 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110100; // iC=-2252 
// vC = 14'b0000001101101010; // vC=  874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b0000001001010111; // vC=  599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000111; // iC=-2169 
// vC = 14'b0000001100001101; // vC=  781 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001010; // iC=-2230 
// vC = 14'b0000001001011101; // vC=  605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011010; // iC=-2150 
// vC = 14'b0000001001011101; // vC=  605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010010; // iC=-2094 
// vC = 14'b0000001000100001; // vC=  545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101001; // iC=-2007 
// vC = 14'b0000001010011111; // vC=  671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000010; // iC=-2238 
// vC = 14'b0000001000101111; // vC=  559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000101; // iC=-2171 
// vC = 14'b0000001000001011; // vC=  523 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000111; // iC=-1977 
// vC = 14'b0000001010010011; // vC=  659 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000011; // iC=-2237 
// vC = 14'b0000001100100000; // vC=  800 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101110; // iC=-2258 
// vC = 14'b0000001001001001; // vC=  585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000110; // iC=-2234 
// vC = 14'b0000001000110101; // vC=  565 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010101; // iC=-2091 
// vC = 14'b0000000111011111; // vC=  479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000010; // iC=-2174 
// vC = 14'b0000001000101100; // vC=  556 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001010; // iC=-2230 
// vC = 14'b0000001010000111; // vC=  647 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b0000001010100110; // vC=  678 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100101; // iC=-2011 
// vC = 14'b0000001010110011; // vC=  691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110001; // iC=-2191 
// vC = 14'b0000001001001000; // vC=  584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010010; // iC=-2158 
// vC = 14'b0000001001010000; // vC=  592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b0000001010100001; // vC=  673 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110001; // iC=-2127 
// vC = 14'b0000001011010000; // vC=  720 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110111; // iC=-2185 
// vC = 14'b0000000111000000; // vC=  448 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111101; // iC=-2243 
// vC = 14'b0000001000001100; // vC=  524 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111011; // iC=-2181 
// vC = 14'b0000001001100000; // vC=  608 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000000; // iC=-2240 
// vC = 14'b0000000110010000; // vC=  400 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100001; // iC=-2143 
// vC = 14'b0000000101111100; // vC=  380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100100; // iC=-2140 
// vC = 14'b0000000111110000; // vC=  496 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100100000; // iC=-2272 
// vC = 14'b0000001010010001; // vC=  657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b0000001001010001; // vC=  593 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011101; // iC=-2211 
// vC = 14'b0000000111010001; // vC=  465 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b0000001001000000; // vC=  576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110000; // iC=-2000 
// vC = 14'b0000001000111000; // vC=  568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100001; // iC=-2143 
// vC = 14'b0000001000000100; // vC=  516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010111; // iC=-2153 
// vC = 14'b0000001000011101; // vC=  541 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101101; // iC=-2131 
// vC = 14'b0000000101110100; // vC=  372 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000010; // iC=-2238 
// vC = 14'b0000000110010110; // vC=  406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b0000001000001000; // vC=  520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000000100110000; // vC=  304 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010111; // iC=-2089 
// vC = 14'b0000000111101110; // vC=  494 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b0000000011110110; // vC=  246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b0000000100101111; // vC=  303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110100; // iC=-2060 
// vC = 14'b0000000110010000; // vC=  400 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001000; // iC=-2168 
// vC = 14'b0000000101111110; // vC=  382 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001111; // iC=-2161 
// vC = 14'b0000000011100010; // vC=  226 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100101; // iC=-2139 
// vC = 14'b0000000101110001; // vC=  369 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010110; // iC=-2218 
// vC = 14'b0000000111001011; // vC=  459 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010000; // iC=-1968 
// vC = 14'b0000000101100101; // vC=  357 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101100; // iC=-2068 
// vC = 14'b0000000110010100; // vC=  404 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001110; // iC=-2226 
// vC = 14'b0000000011010001; // vC=  209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b0000000110100011; // vC=  419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011110; // iC=-2146 
// vC = 14'b0000000011011111; // vC=  223 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111010; // iC=-2182 
// vC = 14'b0000000101010110; // vC=  342 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000000011110010; // vC=  242 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b0000000110011101; // vC=  413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100001; // iC=-2143 
// vC = 14'b0000000010001011; // vC=  139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000000010001010; // vC=  138 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101110; // iC=-2258 
// vC = 14'b0000000110000111; // vC=  391 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010000; // iC=-2224 
// vC = 14'b0000000011000111; // vC=  199 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110000; // iC=-2256 
// vC = 14'b0000000010010010; // vC=  146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b0000000001111011; // vC=  123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b0000000010101110; // vC=  174 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b0000000101001110; // vC=  334 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b0000000100111110; // vC=  318 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000000011110000; // vC=  240 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000000100111001; // vC=  313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101011; // iC=-2069 
// vC = 14'b0000000000100000; // vC=   32 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000000011100100; // vC=  228 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000000011101000; // vC=  232 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b0000000001011110; // vC=   94 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001111; // iC=-2225 
// vC = 14'b0000000100001110; // vC=  270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011011; // iC=-2149 
// vC = 14'b0000000000010011; // vC=   19 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000000001100001; // vC=   97 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101101; // iC=-2067 
// vC = 14'b1111111111000101; // vC=  -59 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010110; // iC=-1962 
// vC = 14'b1111111111110111; // vC=   -9 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010110; // iC=-2026 
// vC = 14'b1111111111010000; // vC=  -48 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011000; // iC=-2024 
// vC = 14'b0000000010001000; // vC=  136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101001; // iC=-2071 
// vC = 14'b1111111110011111; // vC=  -97 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010111; // iC=-2153 
// vC = 14'b0000000000100001; // vC=   33 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010101; // iC=-2091 
// vC = 14'b0000000001011011; // vC=   91 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110001; // iC=-1935 
// vC = 14'b1111111110110101; // vC=  -75 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011011; // iC=-2085 
// vC = 14'b0000000001001001; // vC=   73 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111100; // iC=-2116 
// vC = 14'b1111111101100100; // vC= -156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100110; // iC=-2138 
// vC = 14'b1111111110110111; // vC=  -73 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111100; // iC=-1988 
// vC = 14'b1111111110110101; // vC=  -75 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011010; // iC=-2214 
// vC = 14'b1111111110001111; // vC= -113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111100; // iC=-2116 
// vC = 14'b1111111111000010; // vC=  -62 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111111; // iC=-2241 
// vC = 14'b1111111111111010; // vC=   -6 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b1111111111101111; // vC=  -17 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011000; // iC=-2216 
// vC = 14'b1111111100111001; // vC= -199 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010110; // iC=-1962 
// vC = 14'b1111111101011011; // vC= -165 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100001; // iC=-2143 
// vC = 14'b0000000000110010; // vC=   50 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110100; // iC=-2124 
// vC = 14'b0000000000010101; // vC=   21 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b1111111101111001; // vC= -135 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011110; // iC=-2210 
// vC = 14'b1111111110011001; // vC= -103 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101011; // iC=-2133 
// vC = 14'b1111111101100010; // vC= -158 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b1111111101000000; // vC= -192 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b1111111110011010; // vC= -102 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110001; // iC=-1935 
// vC = 14'b1111111011111000; // vC= -264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b1111111111111110; // vC=   -2 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111110; // iC=-2050 
// vC = 14'b1111111111100001; // vC=  -31 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010110; // iC=-1962 
// vC = 14'b1111111101100110; // vC= -154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010110; // iC=-2026 
// vC = 14'b1111111110001011; // vC= -117 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b1111111101000000; // vC= -192 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b1111111110111000; // vC=  -72 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b1111111101100011; // vC= -157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111100; // iC=-2180 
// vC = 14'b1111111110111111; // vC=  -65 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b1111111110001111; // vC= -113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b1111111010010000; // vC= -368 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b1111111101111101; // vC= -131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110010; // iC=-2190 
// vC = 14'b1111111001110111; // vC= -393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001001; // iC=-2039 
// vC = 14'b1111111100110110; // vC= -202 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b1111111010001100; // vC= -372 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010000; // iC=-1904 
// vC = 14'b1111111010001001; // vC= -375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b1111111010101001; // vC= -343 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011101; // iC=-2147 
// vC = 14'b1111111001101011; // vC= -405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b1111111011010010; // vC= -302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b1111111010011110; // vC= -354 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b1111111101000001; // vC= -191 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101100; // iC=-2068 
// vC = 14'b1111111010110010; // vC= -334 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101101; // iC=-2131 
// vC = 14'b1111111000010000; // vC= -496 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b1111111010000010; // vC= -382 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b1111111101000101; // vC= -187 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b1111111100111100; // vC= -196 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b1111111001101110; // vC= -402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b1111111011000100; // vC= -316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010101; // iC=-2091 
// vC = 14'b1111111011101001; // vC= -279 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101010; // iC=-2134 
// vC = 14'b1111111001001100; // vC= -436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b1111111000111100; // vC= -452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010000; // iC=-1904 
// vC = 14'b1111111010101000; // vC= -344 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011010; // iC=-2022 
// vC = 14'b1111110111011111; // vC= -545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111001; // iC=-1991 
// vC = 14'b1111111010010110; // vC= -362 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001101; // iC=-1907 
// vC = 14'b1111111010001011; // vC= -373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b1111111001110000; // vC= -400 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b1111111000000011; // vC= -509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b1111111010100111; // vC= -345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b1111111010010111; // vC= -361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111000; // iC=-2120 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000100; // iC=-2044 
// vC = 14'b1111111001001010; // vC= -438 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100100; // iC=-1884 
// vC = 14'b1111111000011100; // vC= -484 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001001; // iC=-1847 
// vC = 14'b1111110110110100; // vC= -588 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b1111111000110101; // vC= -459 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b1111111001000110; // vC= -442 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b1111111010010000; // vC= -368 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111100; // iC=-2116 
// vC = 14'b1111110111010110; // vC= -554 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b1111110110000101; // vC= -635 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b1111110111101111; // vC= -529 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b1111110110100011; // vC= -605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000101; // iC=-2043 
// vC = 14'b1111110111111100; // vC= -516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000110; // iC=-1786 
// vC = 14'b1111111001000010; // vC= -446 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101100; // iC=-2068 
// vC = 14'b1111110100101101; // vC= -723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b1111110100100000; // vC= -736 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111110; // iC=-1794 
// vC = 14'b1111110101010101; // vC= -683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001010; // iC=-1782 
// vC = 14'b1111111000000011; // vC= -509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b1111110101110101; // vC= -651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b1111111000101011; // vC= -469 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b1111111000011110; // vC= -482 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b1111110101000010; // vC= -702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b1111110110110111; // vC= -585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100001; // iC=-1887 
// vC = 14'b1111110101000001; // vC= -703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b1111110110010001; // vC= -623 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010110; // iC=-1962 
// vC = 14'b1111110110111110; // vC= -578 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011010; // iC=-1766 
// vC = 14'b1111110111010011; // vC= -557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b1111110011111010; // vC= -774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b1111110101110001; // vC= -655 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b1111110100110000; // vC= -720 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000010; // iC=-1790 
// vC = 14'b1111110100000101; // vC= -763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101010; // iC=-1814 
// vC = 14'b1111110101011111; // vC= -673 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001110; // iC=-1842 
// vC = 14'b1111110011001101; // vC= -819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b1111110110011011; // vC= -613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001001; // iC=-1719 
// vC = 14'b1111110010110110; // vC= -842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010010; // iC=-1774 
// vC = 14'b1111110011001010; // vC= -822 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110111; // iC=-1801 
// vC = 14'b1111110010100111; // vC= -857 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b1111110110010010; // vC= -622 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111110; // iC=-1794 
// vC = 14'b1111110010110101; // vC= -843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b1111110010100101; // vC= -859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100111; // iC=-1689 
// vC = 14'b1111110011010001; // vC= -815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b1111110010001011; // vC= -885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011011; // iC=-1701 
// vC = 14'b1111110001111100; // vC= -900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b1111110011110011; // vC= -781 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001001; // iC=-1719 
// vC = 14'b1111110010110011; // vC= -845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b1111110100111111; // vC= -705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b1111110011100110; // vC= -794 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b1111110001111001; // vC= -903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011101; // iC=-1827 
// vC = 14'b1111110000100011; // vC= -989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101001; // iC=-1687 
// vC = 14'b1111110100100111; // vC= -729 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111010; // iC=-1862 
// vC = 14'b1111110010010000; // vC= -880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111111; // iC=-1857 
// vC = 14'b1111110011111110; // vC= -770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001100; // iC=-1652 
// vC = 14'b1111101111100110; // vC=-1050 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001001; // iC=-1783 
// vC = 14'b1111110011111100; // vC= -772 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111100; // iC=-1796 
// vC = 14'b1111101111111000; // vC=-1032 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b1111110000000001; // vC=-1023 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001010; // iC=-1910 
// vC = 14'b1111110100001010; // vC= -758 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b1111110010110000; // vC= -848 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100110; // iC=-1690 
// vC = 14'b1111110001100011; // vC= -925 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b1111101111011110; // vC=-1058 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110011; // iC=-1741 
// vC = 14'b1111110011101001; // vC= -791 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000101; // iC=-1851 
// vC = 14'b1111101111110001; // vC=-1039 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100001; // iC=-1631 
// vC = 14'b1111110010100110; // vC= -858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001101; // iC=-1651 
// vC = 14'b1111110000101101; // vC= -979 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b1111101110001011; // vC=-1141 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111100; // iC=-1604 
// vC = 14'b1111110001010100; // vC= -940 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001000; // iC=-1592 
// vC = 14'b1111110000111011; // vC= -965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001100; // iC=-1716 
// vC = 14'b1111110010000100; // vC= -892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001001; // iC=-1655 
// vC = 14'b1111110010001101; // vC= -883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111010; // iC=-1862 
// vC = 14'b1111110010011110; // vC= -866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100011; // iC=-1757 
// vC = 14'b1111110010000100; // vC= -892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100100; // iC=-1820 
// vC = 14'b1111101110110111; // vC=-1097 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111001; // iC=-1607 
// vC = 14'b1111110000110110; // vC= -970 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111100; // iC=-1860 
// vC = 14'b1111110001011101; // vC= -931 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110011; // iC=-1805 
// vC = 14'b1111110000001100; // vC=-1012 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101011; // iC=-1685 
// vC = 14'b1111101110111010; // vC=-1094 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000101; // iC=-1787 
// vC = 14'b1111101110001101; // vC=-1139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111000; // iC=-1672 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011010; // iC=-1830 
// vC = 14'b1111101101111110; // vC=-1154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100100; // iC=-1692 
// vC = 14'b1111101111100011; // vC=-1053 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b1111110001001100; // vC= -948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111001; // iC=-1543 
// vC = 14'b1111110000100010; // vC= -990 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000011; // iC=-1533 
// vC = 14'b1111101101111111; // vC=-1153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011000; // iC=-1704 
// vC = 14'b1111110000101111; // vC= -977 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011111; // iC=-1569 
// vC = 14'b1111101101011000; // vC=-1192 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010011; // iC=-1517 
// vC = 14'b1111101110100111; // vC=-1113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b1111101100011000; // vC=-1256 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101100; // iC=-1748 
// vC = 14'b1111101101100101; // vC=-1179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011100; // iC=-1508 
// vC = 14'b1111101101011001; // vC=-1191 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000010; // iC=-1662 
// vC = 14'b1111101111010101; // vC=-1067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b1111101111010110; // vC=-1066 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101110; // iC=-1554 
// vC = 14'b1111101110010100; // vC=-1132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111111; // iC=-1601 
// vC = 14'b1111101011101100; // vC=-1300 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111000; // iC=-1608 
// vC = 14'b1111101101100000; // vC=-1184 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110110; // iC=-1482 
// vC = 14'b1111101111001010; // vC=-1078 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000000; // iC=-1536 
// vC = 14'b1111101100100101; // vC=-1243 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110011; // iC=-1613 
// vC = 14'b1111101111100111; // vC=-1049 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010001; // iC=-1519 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100011; // iC=-1501 
// vC = 14'b1111101110110100; // vC=-1100 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101110; // iC=-1554 
// vC = 14'b1111101111000011; // vC=-1085 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010000; // iC=-1456 
// vC = 14'b1111101111001011; // vC=-1077 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111101; // iC=-1667 
// vC = 14'b1111101110010001; // vC=-1135 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111010; // iC=-1478 
// vC = 14'b1111101011011000; // vC=-1320 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101100; // iC=-1684 
// vC = 14'b1111101011100110; // vC=-1306 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110010; // iC=-1486 
// vC = 14'b1111101101000001; // vC=-1215 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111100; // iC=-1476 
// vC = 14'b1111101101001100; // vC=-1204 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010101; // iC=-1579 
// vC = 14'b1111101100110101; // vC=-1227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011011; // iC=-1701 
// vC = 14'b1111101110000001; // vC=-1151 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110100; // iC=-1484 
// vC = 14'b1111101010100001; // vC=-1375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010100; // iC=-1452 
// vC = 14'b1111101010001011; // vC=-1397 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000110; // iC=-1658 
// vC = 14'b1111101100001100; // vC=-1268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010111; // iC=-1577 
// vC = 14'b1111101011111110; // vC=-1282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011100; // iC=-1444 
// vC = 14'b1111101100110101; // vC=-1227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000001; // iC=-1535 
// vC = 14'b1111101010101100; // vC=-1364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010111; // iC=-1513 
// vC = 14'b1111101010100010; // vC=-1374 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001010; // iC=-1462 
// vC = 14'b1111101101110001; // vC=-1167 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001011; // iC=-1525 
// vC = 14'b1111101011001100; // vC=-1332 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101010; // iC=-1430 
// vC = 14'b1111101101001110; // vC=-1202 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100101; // iC=-1435 
// vC = 14'b1111101001011010; // vC=-1446 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001001; // iC=-1463 
// vC = 14'b1111101100101110; // vC=-1234 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000100; // iC=-1660 
// vC = 14'b1111101000111111; // vC=-1473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110011; // iC=-1613 
// vC = 14'b1111101001101000; // vC=-1432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110011; // iC=-1421 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000001; // iC=-1407 
// vC = 14'b1111101011101110; // vC=-1298 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100001; // iC=-1631 
// vC = 14'b1111101010101011; // vC=-1365 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011011; // iC=-1637 
// vC = 14'b1111101001101001; // vC=-1431 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001011; // iC=-1333 
// vC = 14'b1111100111101010; // vC=-1558 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010011; // iC=-1517 
// vC = 14'b1111101010111101; // vC=-1347 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000101; // iC=-1467 
// vC = 14'b1111101000111110; // vC=-1474 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010010; // iC=-1454 
// vC = 14'b1111101001000100; // vC=-1468 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011100; // iC=-1508 
// vC = 14'b1111101001111010; // vC=-1414 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001110; // iC=-1586 
// vC = 14'b1111101011000010; // vC=-1342 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101000; // iC=-1304 
// vC = 14'b1111100111011011; // vC=-1573 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101001; // iC=-1495 
// vC = 14'b1111101000100011; // vC=-1501 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001110; // iC=-1394 
// vC = 14'b1111101010111111; // vC=-1345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100101; // iC=-1307 
// vC = 14'b1111100111100100; // vC=-1564 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110100; // iC=-1548 
// vC = 14'b1111100110101111; // vC=-1617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100111; // iC=-1561 
// vC = 14'b1111101001101001; // vC=-1431 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011010; // iC=-1254 
// vC = 14'b1111101010110110; // vC=-1354 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010011; // iC=-1453 
// vC = 14'b1111101010101110; // vC=-1362 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001110; // iC=-1330 
// vC = 14'b1111101000111000; // vC=-1480 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011011; // iC=-1445 
// vC = 14'b1111101010011101; // vC=-1379 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110100; // iC=-1548 
// vC = 14'b1111101010011001; // vC=-1383 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111101; // iC=-1347 
// vC = 14'b1111101010000010; // vC=-1406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001100; // iC=-1460 
// vC = 14'b1111101010110010; // vC=-1358 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100011; // iC=-1373 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101110; // iC=-1298 
// vC = 14'b1111101000101000; // vC=-1496 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110111; // iC=-1289 
// vC = 14'b1111100111110110; // vC=-1546 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101010; // iC=-1302 
// vC = 14'b1111100111111001; // vC=-1543 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000101; // iC=-1403 
// vC = 14'b1111100111110000; // vC=-1552 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100001; // iC=-1183 
// vC = 14'b1111101000101111; // vC=-1489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111010; // iC=-1478 
// vC = 14'b1111100110100010; // vC=-1630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000100; // iC=-1468 
// vC = 14'b1111100110110111; // vC=-1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100001; // iC=-1375 
// vC = 14'b1111101001010011; // vC=-1453 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001111; // iC=-1265 
// vC = 14'b1111101001011100; // vC=-1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011001; // iC=-1447 
// vC = 14'b1111100110001101; // vC=-1651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110011; // iC=-1229 
// vC = 14'b1111100111010100; // vC=-1580 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001100; // iC=-1332 
// vC = 14'b1111101000011111; // vC=-1505 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000111; // iC=-1401 
// vC = 14'b1111100101111000; // vC=-1672 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001100; // iC=-1268 
// vC = 14'b1111100101011110; // vC=-1698 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011111; // iC=-1377 
// vC = 14'b1111100111101001; // vC=-1559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111111; // iC=-1153 
// vC = 14'b1111100110011000; // vC=-1640 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100010; // iC=-1374 
// vC = 14'b1111100101000101; // vC=-1723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111110; // iC=-1154 
// vC = 14'b1111100100111111; // vC=-1729 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101100; // iC=-1172 
// vC = 14'b1111100111110101; // vC=-1547 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011101; // iC=-1187 
// vC = 14'b1111100101110000; // vC=-1680 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010100; // iC=-1388 
// vC = 14'b1111100101011100; // vC=-1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111000; // iC=-1288 
// vC = 14'b1111101000010101; // vC=-1515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101110; // iC=-1234 
// vC = 14'b1111100100000001; // vC=-1791 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011101; // iC=-1123 
// vC = 14'b1111100110010110; // vC=-1642 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000011; // iC=-1341 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001000; // iC=-1208 
// vC = 14'b1111101000011001; // vC=-1511 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001010; // iC=-1142 
// vC = 14'b1111100111010010; // vC=-1582 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111001; // iC=-1159 
// vC = 14'b1111100101010011; // vC=-1709 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010001; // iC=-1327 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011001; // iC=-1191 
// vC = 14'b1111100111000100; // vC=-1596 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000111; // iC=-1145 
// vC = 14'b1111100011011001; // vC=-1831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010110; // iC=-1066 
// vC = 14'b1111100101100100; // vC=-1692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111110; // iC=-1090 
// vC = 14'b1111100011011110; // vC=-1826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110000; // iC=-1296 
// vC = 14'b1111100101010000; // vC=-1712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001011; // iC=-1141 
// vC = 14'b1111100011001100; // vC=-1844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101111; // iC=-1041 
// vC = 14'b1111100101001010; // vC=-1718 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100000; // iC=-1056 
// vC = 14'b1111100110001101; // vC=-1651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101111; // iC=-1169 
// vC = 14'b1111100011000110; // vC=-1850 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000001; // iC=-1215 
// vC = 14'b1111100110001001; // vC=-1655 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111110; // iC=-1282 
// vC = 14'b1111100111010110; // vC=-1578 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001110; // iC=-1138 
// vC = 14'b1111100011111000; // vC=-1800 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010000; // iC=-1072 
// vC = 14'b1111100100110111; // vC=-1737 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001000; // iC=-1208 
// vC = 14'b1111100010111101; // vC=-1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100111; // iC=-1049 
// vC = 14'b1111100011010100; // vC=-1836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010000; // iC=-1200 
// vC = 14'b1111100100111100; // vC=-1732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110100; // iC=-1164 
// vC = 14'b1111100011011110; // vC=-1826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100000; // iC= -992 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111100; // iC=-1220 
// vC = 14'b1111100101000101; // vC=-1723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100111; // iC= -985 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011100; // iC=-1060 
// vC = 14'b1111100101101101; // vC=-1683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111001; // iC=-1159 
// vC = 14'b1111100101100110; // vC=-1690 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111011; // iC=-1093 
// vC = 14'b1111100011100100; // vC=-1820 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010011; // iC=-1069 
// vC = 14'b1111100101110001; // vC=-1679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010111; // iC= -937 
// vC = 14'b1111100010011011; // vC=-1893 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000100; // iC=-1020 
// vC = 14'b1111100011110010; // vC=-1806 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011110; // iC=-1186 
// vC = 14'b1111100110010111; // vC=-1641 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101101; // iC= -915 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100001; // iC=-1183 
// vC = 14'b1111100011010110; // vC=-1834 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110011; // iC=-1037 
// vC = 14'b1111100010111100; // vC=-1860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110011; // iC=-1037 
// vC = 14'b1111100001100100; // vC=-1948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110110; // iC=-1098 
// vC = 14'b1111100101100011; // vC=-1693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111000; // iC=-1096 
// vC = 14'b1111100101111011; // vC=-1669 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000100; // iC= -892 
// vC = 14'b1111100001011101; // vC=-1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111110; // iC=-1154 
// vC = 14'b1111100101111100; // vC=-1668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110000; // iC=-1040 
// vC = 14'b1111100010000110; // vC=-1914 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001110; // iC=-1138 
// vC = 14'b1111100001100100; // vC=-1948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011000; // iC=-1000 
// vC = 14'b1111100010100111; // vC=-1881 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010101; // iC=-1131 
// vC = 14'b1111100010100101; // vC=-1883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101111; // iC= -849 
// vC = 14'b1111100010011000; // vC=-1896 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000011; // iC=-1021 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100101; // iC= -987 
// vC = 14'b1111100101100010; // vC=-1694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110100; // iC= -908 
// vC = 14'b1111100101000101; // vC=-1723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000011; // iC= -957 
// vC = 14'b1111100100010110; // vC=-1770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111001; // iC= -839 
// vC = 14'b1111100011011011; // vC=-1829 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111001; // iC= -967 
// vC = 14'b1111100000111000; // vC=-1992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000100; // iC= -764 
// vC = 14'b1111100011001000; // vC=-1848 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001111; // iC= -945 
// vC = 14'b1111100001111111; // vC=-1921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000110; // iC= -954 
// vC = 14'b1111100000111011; // vC=-1989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110110; // iC= -970 
// vC = 14'b1111100000111001; // vC=-1991 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111111; // iC= -897 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011010; // iC= -934 
// vC = 14'b1111100011101100; // vC=-1812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110100; // iC= -972 
// vC = 14'b1111100011000111; // vC=-1849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100100; // iC= -988 
// vC = 14'b1111100001110001; // vC=-1935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010010; // iC= -878 
// vC = 14'b1111100000000101; // vC=-2043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010101; // iC= -747 
// vC = 14'b1111100100011100; // vC=-1764 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001110; // iC= -754 
// vC = 14'b1111100000011111; // vC=-2017 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b1111100010111111; // vC=-1857 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000111; // iC= -761 
// vC = 14'b1111100010111010; // vC=-1862 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111010; // iC= -838 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101001; // iC= -983 
// vC = 14'b1111100001010100; // vC=-1964 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111000; // iC= -840 
// vC = 14'b1111100000100110; // vC=-2010 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010011; // iC= -941 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100010; // iC= -670 
// vC = 14'b1111011111111111; // vC=-2049 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011010; // iC= -742 
// vC = 14'b1111100001010001; // vC=-1967 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010000; // iC= -816 
// vC = 14'b1111100000010010; // vC=-2030 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001001; // iC= -695 
// vC = 14'b1111011111101100; // vC=-2068 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101111; // iC= -849 
// vC = 14'b1111100000101011; // vC=-2005 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011101; // iC= -867 
// vC = 14'b1111100011000100; // vC=-1852 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010001; // iC= -623 
// vC = 14'b1111100011000001; // vC=-1855 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001001; // iC= -887 
// vC = 14'b1111100011010110; // vC=-1834 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011110; // iC= -738 
// vC = 14'b1111100000100000; // vC=-2016 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010000; // iC= -816 
// vC = 14'b1111100010111111; // vC=-1857 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110110; // iC= -586 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001100; // iC= -692 
// vC = 14'b1111100001011010; // vC=-1958 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010010; // iC= -878 
// vC = 14'b1111100001001001; // vC=-1975 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101000; // iC= -664 
// vC = 14'b1111100001001111; // vC=-1969 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000010; // iC= -830 
// vC = 14'b1111100001001110; // vC=-1970 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100111; // iC= -729 
// vC = 14'b1111011111101001; // vC=-2071 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011101; // iC= -611 
// vC = 14'b1111100010011101; // vC=-1891 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000001; // iC= -703 
// vC = 14'b1111100011010101; // vC=-1835 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110100; // iC= -780 
// vC = 14'b1111100000010111; // vC=-2025 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111101; // iC= -771 
// vC = 14'b1111100001000100; // vC=-1980 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111110110; // iC= -522 
// vC = 14'b1111100010000011; // vC=-1917 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011011; // iC= -741 
// vC = 14'b1111100010000110; // vC=-1914 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100100; // iC= -796 
// vC = 14'b1111011111010010; // vC=-2094 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101101; // iC= -659 
// vC = 14'b1111011111011110; // vC=-2082 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111010; // iC= -774 
// vC = 14'b1111100010100000; // vC=-1888 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100101; // iC= -731 
// vC = 14'b1111100000100010; // vC=-2014 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001100; // iC= -500 
// vC = 14'b1111100000010000; // vC=-2032 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111100; // iC= -516 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011001; // iC= -487 
// vC = 14'b1111100010111100; // vC=-1860 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000111; // iC= -633 
// vC = 14'b1111011110011010; // vC=-2150 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110010; // iC= -462 
// vC = 14'b1111100001110011; // vC=-1933 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001001; // iC= -631 
// vC = 14'b1111011110111001; // vC=-2119 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011100; // iC= -548 
// vC = 14'b1111100010011000; // vC=-1896 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110010; // iC= -590 
// vC = 14'b1111100010010000; // vC=-1904 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100000; // iC= -416 
// vC = 14'b1111011111101010; // vC=-2070 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010110; // iC= -426 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010111; // iC= -297 
// vC = 14'b1111100001110010; // vC=-1934 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111010; // iC= -326 
// vC = 14'b1111011111111100; // vC=-2052 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111011; // iC= -325 
// vC = 14'b1111100010011110; // vC=-1890 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001010; // iC= -246 
// vC = 14'b1111100001110111; // vC=-1929 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000110; // iC= -250 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011111; // iC= -225 
// vC = 14'b1111011111101011; // vC=-2069 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000100; // iC= -380 
// vC = 14'b1111100001101100; // vC=-1940 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011000; // iC= -488 
// vC = 14'b1111100010101101; // vC=-1875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010101; // iC= -427 
// vC = 14'b1111011111010111; // vC=-2089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100000; // iC= -160 
// vC = 14'b1111100001001011; // vC=-1973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010011; // iC= -365 
// vC = 14'b1111011110000110; // vC=-2170 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111101; // iC= -131 
// vC = 14'b1111100000010100; // vC=-2028 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111110; // iC= -322 
// vC = 14'b1111011111011101; // vC=-2083 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100111; // iC= -153 
// vC = 14'b1111100001000100; // vC=-1980 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101110000; // iC= -144 
// vC = 14'b1111011110110000; // vC=-2128 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011110; // iC= -290 
// vC = 14'b1111100000110101; // vC=-1995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000001; // iC= -319 
// vC = 14'b1111100001101101; // vC=-1939 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011111; // iC=  -97 
// vC = 14'b1111011110000001; // vC=-2175 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100110; // iC= -218 
// vC = 14'b1111011111100100; // vC=-2076 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101101; // iC= -147 
// vC = 14'b1111100000001100; // vC=-2036 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001101; // iC=  -51 
// vC = 14'b1111100010110111; // vC=-1865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110110011; // iC=  -77 
// vC = 14'b1111100010110001; // vC=-1871 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000111010; // iC=   58 
// vC = 14'b1111100010001011; // vC=-1909 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101111; // iC= -209 
// vC = 14'b1111100000010110; // vC=-2026 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001100; // iC=  -52 
// vC = 14'b1111100010100000; // vC=-1888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100001; // iC=  -95 
// vC = 14'b1111100010110101; // vC=-1867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111011001; // iC=  -39 
// vC = 14'b1111100000001011; // vC=-2037 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110110110; // iC=  -74 
// vC = 14'b1111011101111001; // vC=-2183 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101101; // iC=  -19 
// vC = 14'b1111100000100101; // vC=-2011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111011; // iC=  187 
// vC = 14'b1111100010010001; // vC=-1903 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101111; // iC=  111 
// vC = 14'b1111011110001111; // vC=-2161 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010100; // iC=  212 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011011000; // iC=  216 
// vC = 14'b1111100001101110; // vC=-1938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001001; // iC=    9 
// vC = 14'b1111100000110100; // vC=-1996 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100111; // iC=  103 
// vC = 14'b1111011111010011; // vC=-2093 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001111; // iC=  207 
// vC = 14'b1111011110001100; // vC=-2164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111001; // iC=  185 
// vC = 14'b1111011110011111; // vC=-2145 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110010; // iC=  114 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000001; // iC=  193 
// vC = 14'b1111100001110011; // vC=-1933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010100; // iC=  340 
// vC = 14'b1111011111010011; // vC=-2093 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101100; // iC=  300 
// vC = 14'b1111100000001011; // vC=-2037 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001011; // iC=  267 
// vC = 14'b1111011110100101; // vC=-2139 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001101; // iC=  397 
// vC = 14'b1111011110111100; // vC=-2116 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011110; // iC=  542 
// vC = 14'b1111011111101011; // vC=-2069 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100101; // iC=  549 
// vC = 14'b1111100000100110; // vC=-2010 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000100; // iC=  580 
// vC = 14'b1111100010000100; // vC=-1916 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100101; // iC=  357 
// vC = 14'b1111100001010001; // vC=-1967 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111001; // iC=  569 
// vC = 14'b1111011111010010; // vC=-2094 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010000; // iC=  592 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111011; // iC=  379 
// vC = 14'b1111011111011000; // vC=-2088 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000010; // iC=  514 
// vC = 14'b1111011111000111; // vC=-2105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110000; // iC=  432 
// vC = 14'b1111100001100011; // vC=-1949 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011010; // iC=  538 
// vC = 14'b1111100010000011; // vC=-1917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101011; // iC=  555 
// vC = 14'b1111100000000011; // vC=-2045 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011110; // iC=  606 
// vC = 14'b1111100011001011; // vC=-1845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011111; // iC=  735 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011111; // iC=  799 
// vC = 14'b1111011111100101; // vC=-2075 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100011; // iC=  803 
// vC = 14'b1111100011001110; // vC=-1842 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111000; // iC=  824 
// vC = 14'b1111100000101111; // vC=-2001 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000101; // iC=  901 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001011; // iC=  715 
// vC = 14'b1111011111001000; // vC=-2104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011101; // iC=  797 
// vC = 14'b1111100001001110; // vC=-1970 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010110; // iC=  726 
// vC = 14'b1111100010011001; // vC=-1895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101111; // iC=  879 
// vC = 14'b1111011111000110; // vC=-2106 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100111; // iC=  935 
// vC = 14'b1111100001010101; // vC=-1963 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101100; // iC=  748 
// vC = 14'b1111100001100001; // vC=-1951 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011101; // iC=  989 
// vC = 14'b1111100100000011; // vC=-1789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011110; // iC=  798 
// vC = 14'b1111100000110101; // vC=-1995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011111; // iC=  927 
// vC = 14'b1111011111110110; // vC=-2058 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010001; // iC= 1105 
// vC = 14'b1111100010000101; // vC=-1915 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011000; // iC=  920 
// vC = 14'b1111100010101010; // vC=-1878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011001; // iC= 1049 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100000; // iC= 1120 
// vC = 14'b1111100001010010; // vC=-1966 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110100; // iC= 1204 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101001; // iC= 1129 
// vC = 14'b1111100000100011; // vC=-2013 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011001; // iC= 1113 
// vC = 14'b1111100001011111; // vC=-1953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100100; // iC= 1124 
// vC = 14'b1111100001011001; // vC=-1959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101101; // iC= 1005 
// vC = 14'b1111100011001010; // vC=-1846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011110; // iC= 1054 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001010; // iC= 1354 
// vC = 14'b1111100101001000; // vC=-1720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010111; // iC= 1111 
// vC = 14'b1111100010000010; // vC=-1918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001011; // iC= 1163 
// vC = 14'b1111100011111011; // vC=-1797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101011; // iC= 1195 
// vC = 14'b1111100010100111; // vC=-1881 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111110; // iC= 1150 
// vC = 14'b1111100011110010; // vC=-1806 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000001; // iC= 1409 
// vC = 14'b1111100000101100; // vC=-2004 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011101; // iC= 1245 
// vC = 14'b1111100001010100; // vC=-1964 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010001; // iC= 1425 
// vC = 14'b1111100101101110; // vC=-1682 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000011; // iC= 1347 
// vC = 14'b1111100100010111; // vC=-1769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100101; // iC= 1317 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000011; // iC= 1283 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110001; // iC= 1329 
// vC = 14'b1111100110000110; // vC=-1658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010111; // iC= 1431 
// vC = 14'b1111100110000011; // vC=-1661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100000; // iC= 1568 
// vC = 14'b1111100100011100; // vC=-1764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010110; // iC= 1558 
// vC = 14'b1111100101101001; // vC=-1687 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101011; // iC= 1451 
// vC = 14'b1111100011011111; // vC=-1825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100111; // iC= 1511 
// vC = 14'b1111100101010100; // vC=-1708 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010001; // iC= 1617 
// vC = 14'b1111100010000011; // vC=-1917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110101; // iC= 1525 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000000; // iC= 1472 
// vC = 14'b1111100010110000; // vC=-1872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000010; // iC= 1666 
// vC = 14'b1111100100010110; // vC=-1770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010011; // iC= 1683 
// vC = 14'b1111100010110101; // vC=-1867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000001; // iC= 1473 
// vC = 14'b1111100111001000; // vC=-1592 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100110; // iC= 1446 
// vC = 14'b1111100110001100; // vC=-1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011100; // iC= 1756 
// vC = 14'b1111100010110100; // vC=-1868 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000110; // iC= 1670 
// vC = 14'b1111100010111101; // vC=-1859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011001; // iC= 1689 
// vC = 14'b1111100111011110; // vC=-1570 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111111; // iC= 1663 
// vC = 14'b1111100111011011; // vC=-1573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001001; // iC= 1609 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001111; // iC= 1807 
// vC = 14'b1111100011011110; // vC=-1826 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001001; // iC= 1609 
// vC = 14'b1111100110011011; // vC=-1637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000011; // iC= 1667 
// vC = 14'b1111101000000000; // vC=-1536 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000001; // iC= 1601 
// vC = 14'b1111100110011001; // vC=-1639 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011011; // iC= 1755 
// vC = 14'b1111100111101101; // vC=-1555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111001; // iC= 1593 
// vC = 14'b1111100101101100; // vC=-1684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110011; // iC= 1651 
// vC = 14'b1111100111011010; // vC=-1574 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001011; // iC= 1675 
// vC = 14'b1111100110001001; // vC=-1655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111000; // iC= 1720 
// vC = 14'b1111100111011110; // vC=-1570 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100000; // iC= 1888 
// vC = 14'b1111101000101110; // vC=-1490 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011001; // iC= 1689 
// vC = 14'b1111100101110110; // vC=-1674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010100; // iC= 1748 
// vC = 14'b1111100101000101; // vC=-1723 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000011; // iC= 1667 
// vC = 14'b1111101000111001; // vC=-1479 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001010; // iC= 1866 
// vC = 14'b1111101001110100; // vC=-1420 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111100110001011; // vC=-1653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101100; // iC= 1708 
// vC = 14'b1111100111100100; // vC=-1564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111101001111011; // vC=-1413 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111100; // iC= 1724 
// vC = 14'b1111100101011101; // vC=-1699 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b1111101000001111; // vC=-1521 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b1111100101111101; // vC=-1667 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000001; // iC= 1857 
// vC = 14'b1111100110100100; // vC=-1628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011101; // iC= 1885 
// vC = 14'b1111100111000011; // vC=-1597 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001110; // iC= 1870 
// vC = 14'b1111101010000010; // vC=-1406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b1111100111111101; // vC=-1539 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110111; // iC= 2039 
// vC = 14'b1111100111011011; // vC=-1573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101111; // iC= 1967 
// vC = 14'b1111101010100000; // vC=-1376 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001111; // iC= 2063 
// vC = 14'b1111101011000111; // vC=-1337 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b1111101001110101; // vC=-1419 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110100; // iC= 1844 
// vC = 14'b1111100111100100; // vC=-1564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010010; // iC= 1874 
// vC = 14'b1111101001001100; // vC=-1460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b1111101011101011; // vC=-1301 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001000; // iC= 1800 
// vC = 14'b1111101000111111; // vC=-1473 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001101; // iC= 1997 
// vC = 14'b1111101011110000; // vC=-1296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b1111100111111011; // vC=-1541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101111; // iC= 1967 
// vC = 14'b1111101010100101; // vC=-1371 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b1111101011011111; // vC=-1313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b1111101010010100; // vC=-1388 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100111; // iC= 1831 
// vC = 14'b1111101011000110; // vC=-1338 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110001; // iC= 1969 
// vC = 14'b1111101001010001; // vC=-1455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b1111101010110100; // vC=-1356 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b1111101010000000; // vC=-1408 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011111; // iC= 1887 
// vC = 14'b1111101101010000; // vC=-1200 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b1111101101100110; // vC=-1178 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b1111101010010000; // vC=-1392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111110; // iC= 2174 
// vC = 14'b1111101101001101; // vC=-1203 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b1111101100111101; // vC=-1219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111110; // iC= 1854 
// vC = 14'b1111101101100010; // vC=-1182 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111101011110000; // vC=-1296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000100; // iC= 2116 
// vC = 14'b1111101101101101; // vC=-1171 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b1111101011000001; // vC=-1343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000000; // iC= 2112 
// vC = 14'b1111101110010000; // vC=-1136 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b1111101101010110; // vC=-1194 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111111; // iC= 2111 
// vC = 14'b1111101100101010; // vC=-1238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001011; // iC= 1995 
// vC = 14'b1111101101001100; // vC=-1204 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111101110110101; // vC=-1099 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001101; // iC= 2125 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111101011111110; // vC=-1282 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011100; // iC= 1948 
// vC = 14'b1111101011010010; // vC=-1326 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b1111101111001001; // vC=-1079 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111001; // iC= 2105 
// vC = 14'b1111101111000111; // vC=-1081 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001000; // iC= 2184 
// vC = 14'b1111101111000110; // vC=-1082 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001111; // iC= 1999 
// vC = 14'b1111101100011101; // vC=-1251 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110110; // iC= 2166 
// vC = 14'b1111101100111100; // vC=-1220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110110; // iC= 2102 
// vC = 14'b1111101110010100; // vC=-1132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b1111101101000001; // vC=-1215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101111; // iC= 2159 
// vC = 14'b1111101110100010; // vC=-1118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101000; // iC= 2024 
// vC = 14'b1111101100100111; // vC=-1241 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100000; // iC= 2016 
// vC = 14'b1111110000101111; // vC= -977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b1111101101001101; // vC=-1203 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b1111101101011001; // vC=-1191 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110001; // iC= 1905 
// vC = 14'b1111110000100011; // vC= -989 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100010; // iC= 2210 
// vC = 14'b1111101110111111; // vC=-1089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110011; // iC= 2227 
// vC = 14'b1111101110011100; // vC=-1124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111101101101000; // vC=-1176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111101111000110; // vC=-1082 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111110001011001; // vC= -935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110000; // iC= 2160 
// vC = 14'b1111110001000010; // vC= -958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100100; // iC= 2212 
// vC = 14'b1111110000010100; // vC=-1004 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b1111110000011110; // vC= -994 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000101; // iC= 1925 
// vC = 14'b1111110010011000; // vC= -872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100111; // iC= 2215 
// vC = 14'b1111110011000110; // vC= -826 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000100; // iC= 1988 
// vC = 14'b1111110000110111; // vC= -969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000011; // iC= 2051 
// vC = 14'b1111101111001100; // vC=-1076 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111110001110110; // vC= -906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110000; // iC= 2032 
// vC = 14'b1111110011000111; // vC= -825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101010; // iC= 2154 
// vC = 14'b1111101111001100; // vC=-1076 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111001; // iC= 2169 
// vC = 14'b1111110000001101; // vC=-1011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100011; // iC= 2211 
// vC = 14'b1111101111010101; // vC=-1067 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011010; // iC= 2202 
// vC = 14'b1111110001110111; // vC= -905 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111110010011001; // vC= -871 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011101; // iC= 2205 
// vC = 14'b1111110010100101; // vC= -859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100001; // iC= 2017 
// vC = 14'b1111110000100110; // vC= -986 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b1111110000001011; // vC=-1013 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b1111110000011010; // vC= -998 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b1111110001101110; // vC= -914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101110; // iC= 1966 
// vC = 14'b1111110000111101; // vC= -963 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b1111110011101011; // vC= -789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011001; // iC= 2201 
// vC = 14'b1111110010011111; // vC= -865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101110; // iC= 2222 
// vC = 14'b1111110101001110; // vC= -690 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011100; // iC= 2076 
// vC = 14'b1111110010010010; // vC= -878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111011; // iC= 2171 
// vC = 14'b1111110010010101; // vC= -875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b1111110101000100; // vC= -700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b1111110010100001; // vC= -863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010011; // iC= 2195 
// vC = 14'b1111110100011101; // vC= -739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b1111110011101101; // vC= -787 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100111; // iC= 2023 
// vC = 14'b1111110011101010; // vC= -790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101111; // iC= 2223 
// vC = 14'b1111110010111110; // vC= -834 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000100; // iC= 2180 
// vC = 14'b1111110010110101; // vC= -843 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b1111110100000010; // vC= -766 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101000; // iC= 2152 
// vC = 14'b1111110011100011; // vC= -797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b1111110110010000; // vC= -624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111110110101001; // vC= -599 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000101; // iC= 2181 
// vC = 14'b1111110111000111; // vC= -569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000010; // iC= 1986 
// vC = 14'b1111110111101011; // vC= -533 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b1111110100101000; // vC= -728 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100111; // iC= 2215 
// vC = 14'b1111110100000010; // vC= -766 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b1111110011110101; // vC= -779 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000111; // iC= 2247 
// vC = 14'b1111110110000000; // vC= -640 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010010; // iC= 2194 
// vC = 14'b1111110100000001; // vC= -767 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111010; // iC= 1978 
// vC = 14'b1111110101100000; // vC= -672 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100101; // iC= 1957 
// vC = 14'b1111111001000010; // vC= -446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110101; // iC= 2229 
// vC = 14'b1111111001010001; // vC= -431 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000100; // iC= 2116 
// vC = 14'b1111110100011110; // vC= -738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010101; // iC= 2261 
// vC = 14'b1111111000101001; // vC= -471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001000; // iC= 1992 
// vC = 14'b1111110100111010; // vC= -710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100101; // iC= 2213 
// vC = 14'b1111111000111011; // vC= -453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111011; // iC= 2171 
// vC = 14'b1111110111111010; // vC= -518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011011; // iC= 2139 
// vC = 14'b1111111000010101; // vC= -491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b1111110110100001; // vC= -607 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011010; // iC= 2074 
// vC = 14'b1111111010000010; // vC= -382 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b1111111001100010; // vC= -414 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011011; // iC= 2139 
// vC = 14'b1111110101110011; // vC= -653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b1111110111101010; // vC= -534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001110; // iC= 2190 
// vC = 14'b1111110110101101; // vC= -595 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110100; // iC= 2100 
// vC = 14'b1111111010111000; // vC= -328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111011; // iC= 2235 
// vC = 14'b1111111000000011; // vC= -509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110101; // iC= 2165 
// vC = 14'b1111111001001111; // vC= -433 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111100; // iC= 2044 
// vC = 14'b1111111010011000; // vC= -360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b1111111000001100; // vC= -500 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111111011000000; // vC= -320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111111011110001; // vC= -271 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111111; // iC= 2175 
// vC = 14'b1111111001000000; // vC= -448 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b1111110111011000; // vC= -552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100000; // iC= 2208 
// vC = 14'b1111111011110010; // vC= -270 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100011; // iC= 2211 
// vC = 14'b1111111010011110; // vC= -354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010101; // iC= 2261 
// vC = 14'b1111111100001010; // vC= -246 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101001; // iC= 2089 
// vC = 14'b1111111011010001; // vC= -303 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111110; // iC= 2110 
// vC = 14'b1111111011110010; // vC= -270 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110111; // iC= 2167 
// vC = 14'b1111111010000010; // vC= -382 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111100; // iC= 1980 
// vC = 14'b1111111001000010; // vC= -446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000010; // iC= 1986 
// vC = 14'b1111111000011011; // vC= -485 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111111011101111; // vC= -273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110100; // iC= 2036 
// vC = 14'b1111111001101000; // vC= -408 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b1111111010101101; // vC= -339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111100; // iC= 2172 
// vC = 14'b1111111100010001; // vC= -239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000111; // iC= 2055 
// vC = 14'b1111111001111100; // vC= -388 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110101; // iC= 2101 
// vC = 14'b1111111010110111; // vC= -329 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010101; // iC= 2069 
// vC = 14'b1111111101111001; // vC= -135 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001111; // iC= 2191 
// vC = 14'b1111111100111011; // vC= -197 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b1111111010011111; // vC= -353 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011011; // iC= 1947 
// vC = 14'b1111111100010110; // vC= -234 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111100; // iC= 2172 
// vC = 14'b1111111100100101; // vC= -219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111111; // iC= 2175 
// vC = 14'b1111111101100010; // vC= -158 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101111; // iC= 2159 
// vC = 14'b1111111111000001; // vC=  -63 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000011; // iC= 2243 
// vC = 14'b1111111101111110; // vC= -130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011011; // iC= 2203 
// vC = 14'b1111111101101000; // vC= -152 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b1111111110011111; // vC=  -97 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111101; // iC= 2237 
// vC = 14'b1111111100111100; // vC= -196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100111; // iC= 2023 
// vC = 14'b1111111100000110; // vC= -250 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000011; // iC= 2115 
// vC = 14'b1111111011001011; // vC= -309 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110011; // iC= 2227 
// vC = 14'b1111111110001000; // vC= -120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000100; // iC= 1988 
// vC = 14'b1111111111111111; // vC=   -1 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011110; // iC= 2142 
// vC = 14'b0000000000011111; // vC=   31 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b1111111011111101; // vC= -259 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001100; // iC= 2252 
// vC = 14'b0000000000011101; // vC=   29 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b0000000000011000; // vC=   24 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100010; // iC= 2146 
// vC = 14'b1111111111110111; // vC=   -9 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100011; // iC= 2211 
// vC = 14'b1111111101010110; // vC= -170 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000100; // iC= 2180 
// vC = 14'b0000000000100110; // vC=   38 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001001; // iC= 2249 
// vC = 14'b1111111111100110; // vC=  -26 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b1111111101001110; // vC= -178 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000010; // iC= 2114 
// vC = 14'b1111111110010100; // vC= -108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110000; // iC= 2096 
// vC = 14'b1111111101100001; // vC= -159 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111111101011111; // vC= -161 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b0000000001000100; // vC=   68 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b1111111101110010; // vC= -142 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101110; // iC= 2094 
// vC = 14'b0000000001010000; // vC=   80 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111111110110011; // vC=  -77 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b1111111111001000; // vC=  -56 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b0000000000101101; // vC=   45 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001110; // iC= 1934 
// vC = 14'b0000000001011010; // vC=   90 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110000; // iC= 2032 
// vC = 14'b0000000000000011; // vC=    3 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111111110100111; // vC=  -89 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b0000000001101000; // vC=  104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b0000000010000101; // vC=  133 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110111; // iC= 2039 
// vC = 14'b1111111111000111; // vC=  -57 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000000; // iC= 1920 
// vC = 14'b0000000000001010; // vC=   10 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101000; // iC= 2152 
// vC = 14'b1111111111000110; // vC=  -58 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010111; // iC= 2199 
// vC = 14'b0000000010011010; // vC=  154 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010101; // iC= 2133 
// vC = 14'b1111111111100101; // vC=  -27 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000011; // iC= 1923 
// vC = 14'b0000000001101001; // vC=  105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010101; // iC= 2005 
// vC = 14'b0000000001101011; // vC=  107 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100001; // iC= 2145 
// vC = 14'b0000000010001011; // vC=  139 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100011; // iC= 2147 
// vC = 14'b0000000000011010; // vC=   26 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b0000000001011100; // vC=   92 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110111; // iC= 2167 
// vC = 14'b0000000011111010; // vC=  250 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011010; // iC= 2074 
// vC = 14'b0000000100111001; // vC=  313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111111; // iC= 2111 
// vC = 14'b0000000011101111; // vC=  239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000100; // iC= 2180 
// vC = 14'b0000000010111000; // vC=  184 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b0000000010001101; // vC=  141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111100; // iC= 1916 
// vC = 14'b0000000010100001; // vC=  161 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b0000000001000010; // vC=   66 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b0000000100101011; // vC=  299 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b0000000110010011; // vC=  403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b0000000101010111; // vC=  343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101001; // iC= 1897 
// vC = 14'b0000000110000011; // vC=  387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b0000000110010110; // vC=  406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011101; // iC= 2141 
// vC = 14'b0000000100110010; // vC=  306 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b0000000100100110; // vC=  294 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000000; // iC= 2048 
// vC = 14'b0000000110100000; // vC=  416 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111111; // iC= 1983 
// vC = 14'b0000000101100011; // vC=  355 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100000; // iC= 2016 
// vC = 14'b0000000011100001; // vC=  225 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111111; // iC= 1983 
// vC = 14'b0000000010110001; // vC=  177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b0000000100001100; // vC=  268 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001010; // iC= 1994 
// vC = 14'b0000000101010101; // vC=  341 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100010; // iC= 2146 
// vC = 14'b0000000101101011; // vC=  363 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b0000000110000100; // vC=  388 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b0000000111111111; // vC=  511 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100111; // iC= 2151 
// vC = 14'b0000000101010000; // vC=  336 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000101; // iC= 2053 
// vC = 14'b0000000100000101; // vC=  261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101011; // iC= 2155 
// vC = 14'b0000000110111100; // vC=  444 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101101; // iC= 2157 
// vC = 14'b0000000111000111; // vC=  455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b0000000101110001; // vC=  369 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000000100100011; // vC=  291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111011; // iC= 1915 
// vC = 14'b0000000110011101; // vC=  413 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000100; // iC= 1860 
// vC = 14'b0000001001001100; // vC=  588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010111; // iC= 1879 
// vC = 14'b0000001000100101; // vC=  549 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b0000001000100010; // vC=  546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110111; // iC= 1847 
// vC = 14'b0000001001011101; // vC=  605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b0000000111001010; // vC=  458 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101110; // iC= 1902 
// vC = 14'b0000000110001111; // vC=  399 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b0000000111000010; // vC=  450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000000; // iC= 1920 
// vC = 14'b0000000110000001; // vC=  385 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110101; // iC= 1845 
// vC = 14'b0000001000101110; // vC=  558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b0000001001000110; // vC=  582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b0000001000110110; // vC=  566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b0000001001110010; // vC=  626 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111111; // iC= 1983 
// vC = 14'b0000001001000001; // vC=  577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000001000101100; // vC=  556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b0000000111011010; // vC=  474 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011000; // iC= 2072 
// vC = 14'b0000000111110011; // vC=  499 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b0000001001101001; // vC=  617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100110; // iC= 2086 
// vC = 14'b0000001010000101; // vC=  645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001110; // iC= 1806 
// vC = 14'b0000000111101110; // vC=  494 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101011; // iC= 1963 
// vC = 14'b0000000110110001; // vC=  433 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010011; // iC= 2067 
// vC = 14'b0000001011100101; // vC=  741 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100010; // iC= 1890 
// vC = 14'b0000001000110000; // vC=  560 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b0000000111001101; // vC=  461 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000110; // iC= 1798 
// vC = 14'b0000000111111101; // vC=  509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b0000001000000110; // vC=  518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b0000001000001010; // vC=  522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b0000001000001010; // vC=  522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010110; // iC= 1878 
// vC = 14'b0000001010110011; // vC=  691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100001; // iC= 1761 
// vC = 14'b0000001000000111; // vC=  519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b0000001001111001; // vC=  633 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000011; // iC= 1859 
// vC = 14'b0000001011110101; // vC=  757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b0000001000011000; // vC=  536 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000000; // iC= 1920 
// vC = 14'b0000001010110110; // vC=  694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b0000001001110010; // vC=  626 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111110; // iC= 1982 
// vC = 14'b0000001101011011; // vC=  859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100100; // iC= 1764 
// vC = 14'b0000001001011001; // vC=  601 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b0000001010000000; // vC=  640 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b0000001001011101; // vC=  605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111010; // iC= 1978 
// vC = 14'b0000001100011111; // vC=  799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010001; // iC= 1809 
// vC = 14'b0000001011101110; // vC=  750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b0000001100011011; // vC=  795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111010; // iC= 1722 
// vC = 14'b0000001011011100; // vC=  732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011111; // iC= 1759 
// vC = 14'b0000001100101111; // vC=  815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b0000001100110111; // vC=  823 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b0000001011010101; // vC=  725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110000; // iC= 1840 
// vC = 14'b0000001101010010; // vC=  850 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b0000001110101001; // vC=  937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111011; // iC= 1851 
// vC = 14'b0000001010110110; // vC=  694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110010; // iC= 1906 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111000; // iC= 1848 
// vC = 14'b0000001011011100; // vC=  732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001001; // iC= 1673 
// vC = 14'b0000001011100010; // vC=  738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100010; // iC= 1954 
// vC = 14'b0000001010110101; // vC=  693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b0000001011000110; // vC=  710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b0000001100111100; // vC=  828 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011001; // iC= 1817 
// vC = 14'b0000001111101110; // vC= 1006 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010011; // iC= 1875 
// vC = 14'b0000001100111100; // vC=  828 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b0000001101011001; // vC=  857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011110; // iC= 1758 
// vC = 14'b0000001101100011; // vC=  867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111111; // iC= 1791 
// vC = 14'b0000010000010100; // vC= 1044 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111111; // iC= 1855 
// vC = 14'b0000001101001000; // vC=  840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b0000010000000010; // vC= 1026 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000110; // iC= 1862 
// vC = 14'b0000001111000010; // vC=  962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000001; // iC= 1665 
// vC = 14'b0000010000100100; // vC= 1060 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011100; // iC= 1820 
// vC = 14'b0000010000011000; // vC= 1048 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000010; // iC= 1858 
// vC = 14'b0000001110101100; // vC=  940 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010001; // iC= 1745 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b0000010000100110; // vC= 1062 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110100; // iC= 1716 
// vC = 14'b0000001110100100; // vC=  932 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110001; // iC= 1649 
// vC = 14'b0000001101100100; // vC=  868 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101001; // iC= 1769 
// vC = 14'b0000010001100111; // vC= 1127 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100110; // iC= 1638 
// vC = 14'b0000001101101010; // vC=  874 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011000; // iC= 1880 
// vC = 14'b0000001111100110; // vC=  998 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100111; // iC= 1895 
// vC = 14'b0000001110011101; // vC=  925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111010; // iC= 1594 
// vC = 14'b0000001111110111; // vC= 1015 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000011; // iC= 1795 
// vC = 14'b0000010001101011; // vC= 1131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011010; // iC= 1754 
// vC = 14'b0000001111111001; // vC= 1017 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110010; // iC= 1778 
// vC = 14'b0000001110110011; // vC=  947 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101110; // iC= 1582 
// vC = 14'b0000001110001111; // vC=  911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010110; // iC= 1878 
// vC = 14'b0000001111011100; // vC=  988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000000; // iC= 1600 
// vC = 14'b0000001111010001; // vC=  977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011010; // iC= 1562 
// vC = 14'b0000010001111000; // vC= 1144 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b0000010010001010; // vC= 1162 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000011; // iC= 1859 
// vC = 14'b0000001111001001; // vC=  969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101010; // iC= 1834 
// vC = 14'b0000001111100100; // vC=  996 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110001; // iC= 1777 
// vC = 14'b0000010000011110; // vC= 1054 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011110; // iC= 1758 
// vC = 14'b0000010011001111; // vC= 1231 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010001; // iC= 1809 
// vC = 14'b0000010000101110; // vC= 1070 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100001; // iC= 1825 
// vC = 14'b0000001111100100; // vC=  996 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000101; // iC= 1605 
// vC = 14'b0000010010001010; // vC= 1162 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000110; // iC= 1606 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101001; // iC= 1641 
// vC = 14'b0000010011000011; // vC= 1219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001000; // iC= 1544 
// vC = 14'b0000010000001100; // vC= 1036 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001001; // iC= 1737 
// vC = 14'b0000010001000110; // vC= 1094 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011011; // iC= 1819 
// vC = 14'b0000010000010101; // vC= 1045 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110110; // iC= 1782 
// vC = 14'b0000010000100011; // vC= 1059 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010001; // iC= 1553 
// vC = 14'b0000010000011100; // vC= 1052 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001000; // iC= 1736 
// vC = 14'b0000010000101010; // vC= 1066 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000111; // iC= 1479 
// vC = 14'b0000010000000000; // vC= 1024 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000110; // iC= 1670 
// vC = 14'b0000010000011111; // vC= 1055 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100001; // iC= 1569 
// vC = 14'b0000010000010111; // vC= 1047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100000; // iC= 1568 
// vC = 14'b0000010011100011; // vC= 1251 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100011; // iC= 1699 
// vC = 14'b0000010100000001; // vC= 1281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101001; // iC= 1769 
// vC = 14'b0000010001100001; // vC= 1121 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011010; // iC= 1498 
// vC = 14'b0000010010010010; // vC= 1170 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110110; // iC= 1526 
// vC = 14'b0000010010101111; // vC= 1199 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011100; // iC= 1756 
// vC = 14'b0000010001000001; // vC= 1089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001010; // iC= 1482 
// vC = 14'b0000010101011010; // vC= 1370 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011001; // iC= 1625 
// vC = 14'b0000010011110010; // vC= 1266 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101001; // iC= 1705 
// vC = 14'b0000010100011100; // vC= 1308 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100001; // iC= 1441 
// vC = 14'b0000010001111001; // vC= 1145 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011011; // iC= 1499 
// vC = 14'b0000010011111110; // vC= 1278 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111110; // iC= 1726 
// vC = 14'b0000010011011111; // vC= 1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000100; // iC= 1540 
// vC = 14'b0000010011111111; // vC= 1279 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101011; // iC= 1643 
// vC = 14'b0000010100010011; // vC= 1299 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000111; // iC= 1671 
// vC = 14'b0000010100110000; // vC= 1328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111011; // iC= 1531 
// vC = 14'b0000010110011001; // vC= 1433 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001000; // iC= 1480 
// vC = 14'b0000010010111101; // vC= 1213 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011100; // iC= 1564 
// vC = 14'b0000010110101010; // vC= 1450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b0000010010011111; // vC= 1183 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100001; // iC= 1633 
// vC = 14'b0000010011110110; // vC= 1270 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010111; // iC= 1559 
// vC = 14'b0000010100111110; // vC= 1342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000101; // iC= 1413 
// vC = 14'b0000010100011101; // vC= 1309 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111111; // iC= 1471 
// vC = 14'b0000010010111111; // vC= 1215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100101; // iC= 1509 
// vC = 14'b0000010101111010; // vC= 1402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010101; // iC= 1621 
// vC = 14'b0000010111100011; // vC= 1507 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110100; // iC= 1524 
// vC = 14'b0000010110010010; // vC= 1426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010000; // iC= 1552 
// vC = 14'b0000010011000010; // vC= 1218 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100100; // iC= 1572 
// vC = 14'b0000010110001000; // vC= 1416 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011111; // iC= 1567 
// vC = 14'b0000010110001011; // vC= 1419 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111011; // iC= 1531 
// vC = 14'b0000010111111110; // vC= 1534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111000; // iC= 1336 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111001; // iC= 1465 
// vC = 14'b0000010011100000; // vC= 1248 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010011; // iC= 1491 
// vC = 14'b0000010110111110; // vC= 1470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100010; // iC= 1314 
// vC = 14'b0000010111010100; // vC= 1492 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110000; // iC= 1520 
// vC = 14'b0000011000010101; // vC= 1557 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010101; // iC= 1365 
// vC = 14'b0000011000110001; // vC= 1585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111110; // iC= 1406 
// vC = 14'b0000010111101100; // vC= 1516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110101; // iC= 1525 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010111; // iC= 1559 
// vC = 14'b0000010111101010; // vC= 1514 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001111; // iC= 1423 
// vC = 14'b0000011000101001; // vC= 1577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010101; // iC= 1429 
// vC = 14'b0000010101000001; // vC= 1345 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010101; // iC= 1493 
// vC = 14'b0000010101001010; // vC= 1354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011100; // iC= 1436 
// vC = 14'b0000010101001000; // vC= 1352 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001010; // iC= 1546 
// vC = 14'b0000010101011110; // vC= 1374 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011010; // iC= 1434 
// vC = 14'b0000011001010110; // vC= 1622 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010110; // iC= 1430 
// vC = 14'b0000010111101011; // vC= 1515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000100; // iC= 1348 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111100; // iC= 1404 
// vC = 14'b0000011000000010; // vC= 1538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111111; // iC= 1279 
// vC = 14'b0000011010000000; // vC= 1664 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111100; // iC= 1404 
// vC = 14'b0000011000100010; // vC= 1570 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001001; // iC= 1481 
// vC = 14'b0000010101111011; // vC= 1403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100011; // iC= 1507 
// vC = 14'b0000011000010001; // vC= 1553 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010011; // iC= 1427 
// vC = 14'b0000010111101000; // vC= 1512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101110; // iC= 1390 
// vC = 14'b0000010101100010; // vC= 1378 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111010; // iC= 1274 
// vC = 14'b0000011001100011; // vC= 1635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111000; // iC= 1208 
// vC = 14'b0000010110010011; // vC= 1427 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000011; // iC= 1347 
// vC = 14'b0000011000000000; // vC= 1536 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110100; // iC= 1268 
// vC = 14'b0000010101101101; // vC= 1389 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001001; // iC= 1225 
// vC = 14'b0000010110111111; // vC= 1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110111; // iC= 1335 
// vC = 14'b0000011001101111; // vC= 1647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101101; // iC= 1261 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111011; // iC= 1211 
// vC = 14'b0000010110110110; // vC= 1462 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110111; // iC= 1463 
// vC = 14'b0000010111011000; // vC= 1496 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010011; // iC= 1171 
// vC = 14'b0000011000011011; // vC= 1563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001011; // iC= 1355 
// vC = 14'b0000011000010111; // vC= 1559 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110100; // iC= 1140 
// vC = 14'b0000011001011111; // vC= 1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101001; // iC= 1321 
// vC = 14'b0000011000100000; // vC= 1568 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010000; // iC= 1424 
// vC = 14'b0000011001011111; // vC= 1631 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001000; // iC= 1352 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110001; // iC= 1201 
// vC = 14'b0000011001101101; // vC= 1645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010100; // iC= 1428 
// vC = 14'b0000011011010011; // vC= 1747 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101010; // iC= 1322 
// vC = 14'b0000011011011101; // vC= 1757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101100; // iC= 1196 
// vC = 14'b0000011010100110; // vC= 1702 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100001; // iC= 1185 
// vC = 14'b0000011011101001; // vC= 1769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100000; // iC= 1120 
// vC = 14'b0000010111111111; // vC= 1535 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110101; // iC= 1141 
// vC = 14'b0000011001111101; // vC= 1661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011111; // iC= 1119 
// vC = 14'b0000011100000111; // vC= 1799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101000; // iC= 1064 
// vC = 14'b0000010111011110; // vC= 1502 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110110; // iC= 1334 
// vC = 14'b0000011010001010; // vC= 1674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101011; // iC= 1131 
// vC = 14'b0000011011000001; // vC= 1729 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010110; // iC= 1174 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100000; // iC= 1056 
// vC = 14'b0000010111110110; // vC= 1526 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110110; // iC= 1270 
// vC = 14'b0000011011011110; // vC= 1758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111110; // iC= 1278 
// vC = 14'b0000011001000000; // vC= 1600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001101; // iC= 1165 
// vC = 14'b0000011001111010; // vC= 1658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101011; // iC= 1067 
// vC = 14'b0000011010010101; // vC= 1685 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101100; // iC= 1324 
// vC = 14'b0000011100110000; // vC= 1840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000010; // iC= 1282 
// vC = 14'b0000011001100110; // vC= 1638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111110; // iC= 1150 
// vC = 14'b0000011001100110; // vC= 1638 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100100; // iC= 1316 
// vC = 14'b0000011011000110; // vC= 1734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100110; // iC= 1126 
// vC = 14'b0000011101011000; // vC= 1880 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010111; // iC=  983 
// vC = 14'b0000011001011110; // vC= 1630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000110; // iC= 1158 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110110; // iC= 1014 
// vC = 14'b0000011101001111; // vC= 1871 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010100; // iC= 1172 
// vC = 14'b0000011010110111; // vC= 1719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110000; // iC= 1008 
// vC = 14'b0000011001101000; // vC= 1640 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110010; // iC= 1202 
// vC = 14'b0000011100111110; // vC= 1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111010; // iC= 1018 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011100; // iC= 1052 
// vC = 14'b0000011101101101; // vC= 1901 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011100; // iC= 1244 
// vC = 14'b0000011011110100; // vC= 1780 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111001; // iC=  953 
// vC = 14'b0000011001010101; // vC= 1621 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100100; // iC=  932 
// vC = 14'b0000011010111101; // vC= 1725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011000; // iC=  920 
// vC = 14'b0000011001101111; // vC= 1647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001001; // iC=  969 
// vC = 14'b0000011011001011; // vC= 1739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010100; // iC=  980 
// vC = 14'b0000011100110000; // vC= 1840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010110; // iC=  918 
// vC = 14'b0000011101001000; // vC= 1864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010100; // iC=  916 
// vC = 14'b0000011010100100; // vC= 1700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110110; // iC= 1142 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100110; // iC=  998 
// vC = 14'b0000011011001101; // vC= 1741 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011110; // iC=  926 
// vC = 14'b0000011100001111; // vC= 1807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100110; // iC= 1062 
// vC = 14'b0000011100010111; // vC= 1815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010101; // iC=  917 
// vC = 14'b0000011010110110; // vC= 1718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110001; // iC=  945 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010110; // iC=  982 
// vC = 14'b0000011100001101; // vC= 1805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010001; // iC=  849 
// vC = 14'b0000011010000111; // vC= 1671 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010110; // iC=  982 
// vC = 14'b0000011110110001; // vC= 1969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111001; // iC= 1081 
// vC = 14'b0000011111001001; // vC= 1993 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010111; // iC=  983 
// vC = 14'b0000011011010100; // vC= 1748 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010111; // iC= 1111 
// vC = 14'b0000011010100110; // vC= 1702 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001100; // iC= 1036 
// vC = 14'b0000011010100110; // vC= 1702 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111000; // iC=  888 
// vC = 14'b0000011111001001; // vC= 1993 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001110; // iC=  974 
// vC = 14'b0000011011001111; // vC= 1743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000011; // iC= 1027 
// vC = 14'b0000011010111101; // vC= 1725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111111; // iC=  959 
// vC = 14'b0000011010101001; // vC= 1705 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010101; // iC=  917 
// vC = 14'b0000011011011001; // vC= 1753 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001001; // iC=  905 
// vC = 14'b0000011101100000; // vC= 1888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001001; // iC=  841 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011111; // iC=  991 
// vC = 14'b0000011101110111; // vC= 1911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110101; // iC=  821 
// vC = 14'b0000011100010011; // vC= 1811 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110001; // iC=  817 
// vC = 14'b0000011011110111; // vC= 1783 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110010; // iC=  818 
// vC = 14'b0000011101001101; // vC= 1869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011001; // iC=  921 
// vC = 14'b0000011111010000; // vC= 2000 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110010; // iC= 1010 
// vC = 14'b0000011101100000; // vC= 1888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010101; // iC=  917 
// vC = 14'b0000011100111001; // vC= 1849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111000; // iC=  824 
// vC = 14'b0000011100001010; // vC= 1802 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100010; // iC=  866 
// vC = 14'b0000100000001101; // vC= 2061 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001000; // iC=  776 
// vC = 14'b0000011100100010; // vC= 1826 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001100; // iC=  972 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000010; // iC=  834 
// vC = 14'b0000011100110101; // vC= 1845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001100; // iC=  972 
// vC = 14'b0000011101101110; // vC= 1902 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001101; // iC=  717 
// vC = 14'b0000100000001101; // vC= 2061 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001110; // iC=  718 
// vC = 14'b0000011110011100; // vC= 1948 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001111; // iC=  975 
// vC = 14'b0000011111110110; // vC= 2038 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001101; // iC=  845 
// vC = 14'b0000011111010000; // vC= 2000 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001100; // iC=  844 
// vC = 14'b0000011111101100; // vC= 2028 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000001; // iC=  961 
// vC = 14'b0000011110010101; // vC= 1941 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110001; // iC=  689 
// vC = 14'b0000100000001010; // vC= 2058 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111101; // iC=  701 
// vC = 14'b0000011110010001; // vC= 1937 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100101; // iC=  805 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101011; // iC=  747 
// vC = 14'b0000011111101001; // vC= 2025 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111111; // iC=  831 
// vC = 14'b0000011111111101; // vC= 2045 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101101010; // iC=  874 
// vC = 14'b0000100000011010; // vC= 2074 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010101; // iC=  661 
// vC = 14'b0000011111111001; // vC= 2041 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111001; // iC=  825 
// vC = 14'b0000011100000110; // vC= 1798 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100010; // iC=  674 
// vC = 14'b0000011101110110; // vC= 1910 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110011; // iC=  627 
// vC = 14'b0000100001000010; // vC= 2114 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011101; // iC=  797 
// vC = 14'b0000011111010000; // vC= 2000 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100110; // iC=  742 
// vC = 14'b0000100000000111; // vC= 2055 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010110; // iC=  854 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110111; // iC=  567 
// vC = 14'b0000011100110011; // vC= 1843 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110011; // iC=  691 
// vC = 14'b0000011111100011; // vC= 2019 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100100; // iC=  804 
// vC = 14'b0000011111111100; // vC= 2044 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010111; // iC=  727 
// vC = 14'b0000011110100011; // vC= 1955 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110010; // iC=  754 
// vC = 14'b0000100000101111; // vC= 2095 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011001; // iC=  537 
// vC = 14'b0000011101011000; // vC= 1880 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111101; // iC=  701 
// vC = 14'b0000011101001100; // vC= 1868 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101110; // iC=  686 
// vC = 14'b0000100000011011; // vC= 2075 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000000; // iC=  576 
// vC = 14'b0000100000110111; // vC= 2103 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000011; // iC=  451 
// vC = 14'b0000011111011111; // vC= 2015 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111111; // iC=  511 
// vC = 14'b0000100000101101; // vC= 2093 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011101; // iC=  605 
// vC = 14'b0000100000111010; // vC= 2106 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011111; // iC=  671 
// vC = 14'b0000011111101111; // vC= 2031 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000010; // iC=  578 
// vC = 14'b0000100001011110; // vC= 2142 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101101; // iC=  557 
// vC = 14'b0000011101010011; // vC= 1875 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100000; // iC=  608 
// vC = 14'b0000011110100100; // vC= 1956 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001001; // iC=  457 
// vC = 14'b0000011110010101; // vC= 1941 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001011; // iC=  523 
// vC = 14'b0000100001110101; // vC= 2165 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110011; // iC=  371 
// vC = 14'b0000011111011001; // vC= 2009 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000111; // iC=  327 
// vC = 14'b0000100001010011; // vC= 2131 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100010; // iC=  418 
// vC = 14'b0000100000010110; // vC= 2070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100000010; // iC=  258 
// vC = 14'b0000011110001001; // vC= 1929 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000101; // iC=  389 
// vC = 14'b0000100000100000; // vC= 2080 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010111; // iC=  215 
// vC = 14'b0000011110011100; // vC= 1948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101101; // iC=  301 
// vC = 14'b0000011101010101; // vC= 1877 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000000; // iC=  320 
// vC = 14'b0000011101101111; // vC= 1903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001010; // iC=  266 
// vC = 14'b0000011111101001; // vC= 2025 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100110; // iC=  358 
// vC = 14'b0000100001111000; // vC= 2168 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101000; // iC=  232 
// vC = 14'b0000100001010000; // vC= 2128 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101001; // iC=  361 
// vC = 14'b0000011101101010; // vC= 1898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000001; // iC=  129 
// vC = 14'b0000011110001010; // vC= 1930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001110; // iC=  142 
// vC = 14'b0000011110000001; // vC= 1921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100010; // iC=  162 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011011000; // iC=  216 
// vC = 14'b0000011101011000; // vC= 1880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111000; // iC=  248 
// vC = 14'b0000011110110101; // vC= 1973 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010101; // iC=  149 
// vC = 14'b0000100000011010; // vC= 2074 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000000; // iC=  128 
// vC = 14'b0000011101101010; // vC= 1898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101110; // iC=   46 
// vC = 14'b0000100010001110; // vC= 2190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110011; // iC=  243 
// vC = 14'b0000011110001011; // vC= 1931 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010001; // iC=   17 
// vC = 14'b0000011101101000; // vC= 1896 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101110; // iC=   46 
// vC = 14'b0000100000001100; // vC= 2060 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000011; // iC=  195 
// vC = 14'b0000011111010101; // vC= 2005 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111100; // iC=  124 
// vC = 14'b0000100001111000; // vC= 2168 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001100; // iC=  140 
// vC = 14'b0000011111000011; // vC= 1987 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101110; // iC= -146 
// vC = 14'b0000100001110010; // vC= 2162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001111; // iC=  143 
// vC = 14'b0000011101011010; // vC= 1882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100001; // iC=  -31 
// vC = 14'b0000011111001011; // vC= 1995 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101011101; // iC= -163 
// vC = 14'b0000100001010010; // vC= 2130 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111111110; // iC=   -2 
// vC = 14'b0000100001001100; // vC= 2124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001101; // iC= -179 
// vC = 14'b0000011101110011; // vC= 1907 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111011; // iC= -133 
// vC = 14'b0000011110001010; // vC= 1930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111110; // iC=  -66 
// vC = 14'b0000011101010101; // vC= 1877 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000001; // iC= -127 
// vC = 14'b0000011110111010; // vC= 1978 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101110110; // iC= -138 
// vC = 14'b0000011101011101; // vC= 1885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110101; // iC= -331 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000111; // iC= -313 
// vC = 14'b0000100000111110; // vC= 2110 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100111; // iC= -409 
// vC = 14'b0000011111010100; // vC= 2004 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001110; // iC= -242 
// vC = 14'b0000011111100101; // vC= 2021 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000000; // iC= -448 
// vC = 14'b0000100000111101; // vC= 2109 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000110; // iC= -186 
// vC = 14'b0000011101110101; // vC= 1909 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001101; // iC= -435 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010111; // iC= -489 
// vC = 14'b0000011110101001; // vC= 1961 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000011; // iC= -317 
// vC = 14'b0000011111000101; // vC= 1989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011100; // iC= -420 
// vC = 14'b0000011111100110; // vC= 2022 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111100; // iC= -580 
// vC = 14'b0000011111100001; // vC= 2017 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011100; // iC= -612 
// vC = 14'b0000100001110101; // vC= 2165 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101010; // iC= -470 
// vC = 14'b0000100001001000; // vC= 2120 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101111; // iC= -593 
// vC = 14'b0000011111001001; // vC= 1993 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001111; // iC= -625 
// vC = 14'b0000100001100011; // vC= 2147 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011110; // iC= -482 
// vC = 14'b0000011110100100; // vC= 1956 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110010111; // iC= -617 
// vC = 14'b0000011111100101; // vC= 2021 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000111; // iC= -761 
// vC = 14'b0000011111010101; // vC= 2005 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001011; // iC= -757 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011000; // iC= -616 
// vC = 14'b0000011110010011; // vC= 1939 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011001; // iC= -679 
// vC = 14'b0000011101110111; // vC= 1911 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100111; // iC= -601 
// vC = 14'b0000011111100001; // vC= 2017 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101100; // iC= -724 
// vC = 14'b0000011100111011; // vC= 1851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110101; // iC= -651 
// vC = 14'b0000011110010000; // vC= 1936 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111100; // iC= -836 
// vC = 14'b0000011110111100; // vC= 1980 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010110; // iC= -810 
// vC = 14'b0000100000000101; // vC= 2053 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000011; // iC= -701 
// vC = 14'b0000011111111000; // vC= 2040 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111010; // iC= -774 
// vC = 14'b0000100000111000; // vC= 2104 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111000; // iC= -712 
// vC = 14'b0000011111101000; // vC= 2024 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110001; // iC= -847 
// vC = 14'b0000011111101111; // vC= 2031 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110000; // iC= -912 
// vC = 14'b0000011100010101; // vC= 1813 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001000; // iC=-1016 
// vC = 14'b0000011111111100; // vC= 2044 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001011; // iC=-1077 
// vC = 14'b0000011101111101; // vC= 1917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001011; // iC= -821 
// vC = 14'b0000011111100101; // vC= 2021 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111000; // iC=-1096 
// vC = 14'b0000011111101101; // vC= 2029 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001001; // iC=-1079 
// vC = 14'b0000011100010000; // vC= 1808 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010001; // iC=-1071 
// vC = 14'b0000011111110101; // vC= 2037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001000; // iC=-1016 
// vC = 14'b0000011111101010; // vC= 2026 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110111; // iC= -969 
// vC = 14'b0000011111011010; // vC= 2010 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000110; // iC= -954 
// vC = 14'b0000011110011100; // vC= 1948 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010000; // iC=-1008 
// vC = 14'b0000011111110010; // vC= 2034 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001011; // iC=-1013 
// vC = 14'b0000011111011001; // vC= 2009 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111000; // iC=-1096 
// vC = 14'b0000011101101100; // vC= 1900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011011; // iC=-1189 
// vC = 14'b0000011101111110; // vC= 1918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110111; // iC=-1097 
// vC = 14'b0000011011110011; // vC= 1779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111100; // iC=-1220 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111111; // iC=-1345 
// vC = 14'b0000011110011000; // vC= 1944 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110010; // iC=-1230 
// vC = 14'b0000011101011000; // vC= 1880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100000; // iC=-1312 
// vC = 14'b0000011101110000; // vC= 1904 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100110; // iC=-1434 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110011; // iC=-1293 
// vC = 14'b0000011011000011; // vC= 1731 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110100; // iC=-1484 
// vC = 14'b0000011110101010; // vC= 1962 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011000; // iC=-1512 
// vC = 14'b0000011110101111; // vC= 1967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011101; // iC=-1315 
// vC = 14'b0000011011111001; // vC= 1785 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101001; // iC=-1367 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111101; // iC=-1475 
// vC = 14'b0000011011001101; // vC= 1741 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001111; // iC=-1521 
// vC = 14'b0000011010110001; // vC= 1713 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100101; // iC=-1435 
// vC = 14'b0000011001100100; // vC= 1636 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110101; // iC=-1419 
// vC = 14'b0000011001100000; // vC= 1632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010010; // iC=-1518 
// vC = 14'b0000011101011110; // vC= 1886 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111010; // iC=-1414 
// vC = 14'b0000011010000011; // vC= 1667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110100; // iC=-1420 
// vC = 14'b0000011001010100; // vC= 1620 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100011; // iC=-1629 
// vC = 14'b0000011010000001; // vC= 1665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100010; // iC=-1438 
// vC = 14'b0000011010101001; // vC= 1705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001011; // iC=-1461 
// vC = 14'b0000011100010111; // vC= 1815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000101; // iC=-1467 
// vC = 14'b0000011101011100; // vC= 1884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001110; // iC=-1522 
// vC = 14'b0000011011100011; // vC= 1763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111101; // iC=-1603 
// vC = 14'b0000011010000001; // vC= 1665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100010; // iC=-1694 
// vC = 14'b0000011100001100; // vC= 1804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011110; // iC=-1506 
// vC = 14'b0000011100101101; // vC= 1837 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111110; // iC=-1538 
// vC = 14'b0000011000001111; // vC= 1551 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100000; // iC=-1632 
// vC = 14'b0000011001011010; // vC= 1626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010011; // iC=-1709 
// vC = 14'b0000011001011101; // vC= 1629 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101101; // iC=-1619 
// vC = 14'b0000011000001010; // vC= 1546 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011111; // iC=-1633 
// vC = 14'b0000011001101100; // vC= 1644 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111110; // iC=-1666 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101111; // iC=-1809 
// vC = 14'b0000011010110100; // vC= 1716 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011010; // iC=-1702 
// vC = 14'b0000011010010101; // vC= 1685 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001001; // iC=-1719 
// vC = 14'b0000011000111010; // vC= 1594 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b0000011001111010; // vC= 1658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001110; // iC=-1714 
// vC = 14'b0000011000100001; // vC= 1569 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010101; // iC=-1707 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000011; // iC=-1725 
// vC = 14'b0000010111010111; // vC= 1495 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b0000011000101000; // vC= 1576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001101; // iC=-1907 
// vC = 14'b0000011000011111; // vC= 1567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b0000011010100000; // vC= 1696 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111000; // iC=-1736 
// vC = 14'b0000011000011001; // vC= 1561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b0000011010001101; // vC= 1677 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010010; // iC=-1774 
// vC = 14'b0000011001100000; // vC= 1632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001111; // iC=-1777 
// vC = 14'b0000010111101011; // vC= 1515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101110; // iC=-1874 
// vC = 14'b0000010110100100; // vC= 1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b0000011000010101; // vC= 1557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101001; // iC=-1879 
// vC = 14'b0000010101000101; // vC= 1349 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b0000010111000101; // vC= 1477 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001100; // iC=-1908 
// vC = 14'b0000011000011011; // vC= 1563 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110101; // iC=-1803 
// vC = 14'b0000011000001110; // vC= 1550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100011; // iC=-2077 
// vC = 14'b0000010111010001; // vC= 1489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010110; // iC=-2026 
// vC = 14'b0000010101101100; // vC= 1388 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111001; // iC=-1991 
// vC = 14'b0000010110101100; // vC= 1452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000010101100111; // vC= 1383 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b0000010100100010; // vC= 1314 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b0000010110110110; // vC= 1462 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b0000010101001111; // vC= 1359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b0000010101000011; // vC= 1347 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000010100100100; // vC= 1316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110001; // iC=-1935 
// vC = 14'b0000010101011011; // vC= 1371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100100; // iC=-1884 
// vC = 14'b0000010101000110; // vC= 1350 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b0000010111101011; // vC= 1515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011001; // iC=-2151 
// vC = 14'b0000010011100110; // vC= 1254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110010; // iC=-1870 
// vC = 14'b0000010101011010; // vC= 1370 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b0000010110010011; // vC= 1427 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000010011000111; // vC= 1223 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000101; // iC=-2107 
// vC = 14'b0000010101100000; // vC= 1376 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000010010111000; // vC= 1208 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100000; // iC=-2080 
// vC = 14'b0000010101000110; // vC= 1350 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000010100100111; // vC= 1319 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b0000010001110110; // vC= 1142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000010110100100; // vC= 1444 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101101; // iC=-2067 
// vC = 14'b0000010010101100; // vC= 1196 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111001; // iC=-1927 
// vC = 14'b0000010011011010; // vC= 1242 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000100; // iC=-1916 
// vC = 14'b0000010001011001; // vC= 1113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010110; // iC=-2154 
// vC = 14'b0000010010111110; // vC= 1214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001100; // iC=-1908 
// vC = 14'b0000010010010011; // vC= 1171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b0000010010000010; // vC= 1154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b0000010010111111; // vC= 1215 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000010001011111; // vC= 1119 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101010; // iC=-2070 
// vC = 14'b0000010001011110; // vC= 1118 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000000; // iC=-2176 
// vC = 14'b0000010011100100; // vC= 1252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011100; // iC=-1956 
// vC = 14'b0000010100010010; // vC= 1298 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b0000010000110111; // vC= 1079 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111111; // iC=-1985 
// vC = 14'b0000010000110110; // vC= 1078 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b0000010001110110; // vC= 1142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100001; // iC=-2143 
// vC = 14'b0000010001100111; // vC= 1127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b0000001111100100; // vC=  996 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011111; // iC=-2145 
// vC = 14'b0000010001110001; // vC= 1137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100000; // iC=-1952 
// vC = 14'b0000010001001001; // vC= 1097 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111001; // iC=-2119 
// vC = 14'b0000001110111111; // vC=  959 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b0000001110111100; // vC=  956 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011101; // iC=-2147 
// vC = 14'b0000010010111110; // vC= 1214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011000; // iC=-2216 
// vC = 14'b0000010011100010; // vC= 1250 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100101; // iC=-2203 
// vC = 14'b0000001111011011; // vC=  987 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110100; // iC=-1932 
// vC = 14'b0000001110100000; // vC=  928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b0000010011001011; // vC= 1227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b0000010001100011; // vC= 1123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100101; // iC=-2075 
// vC = 14'b0000010001111011; // vC= 1147 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100101; // iC=-2011 
// vC = 14'b0000010001010101; // vC= 1109 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000011; // iC=-2173 
// vC = 14'b0000001110101110; // vC=  942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b0000001111100110; // vC=  998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000001111011001; // vC=  985 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100010; // iC=-2014 
// vC = 14'b0000010000101100; // vC= 1068 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010000; // iC=-2160 
// vC = 14'b0000001111011101; // vC=  989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b0000001101101111; // vC=  879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001001; // iC=-2039 
// vC = 14'b0000001110001011; // vC=  907 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011011; // iC=-2085 
// vC = 14'b0000001110011000; // vC=  920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000010000000100; // vC= 1028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000111; // iC=-2233 
// vC = 14'b0000001110000001; // vC=  897 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011111; // iC=-2145 
// vC = 14'b0000001110011100; // vC=  924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b0000001111011000; // vC=  984 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110100; // iC=-2188 
// vC = 14'b0000010000000100; // vC= 1028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b0000001111110001; // vC= 1009 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b0000001100101011; // vC=  811 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b0000001101010110; // vC=  854 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110000; // iC=-2064 
// vC = 14'b0000001111000111; // vC=  967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b0000001111100010; // vC=  994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b0000001111010010; // vC=  978 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b0000001101011001; // vC=  857 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110000; // iC=-2000 
// vC = 14'b0000001101110010; // vC=  882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101011; // iC=-2197 
// vC = 14'b0000001110010101; // vC=  917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000001110111010; // vC=  954 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b0000001110111110; // vC=  958 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100011; // iC=-2077 
// vC = 14'b0000001101110101; // vC=  885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111110; // iC=-2178 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010001; // iC=-2095 
// vC = 14'b0000001110011010; // vC=  922 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b0000001010100010; // vC=  674 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101101; // iC=-2131 
// vC = 14'b0000001110011110; // vC=  926 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b0000001101101110; // vC=  878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001001; // iC=-2103 
// vC = 14'b0000001101011111; // vC=  863 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101110; // iC=-2258 
// vC = 14'b0000001011111110; // vC=  766 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b0000001101100001; // vC=  865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001011; // iC=-2165 
// vC = 14'b0000001011001000; // vC=  712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000001010100000; // vC=  672 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000001011111011; // vC=  763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b0000001010110001; // vC=  689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011010; // iC=-2214 
// vC = 14'b0000001011001100; // vC=  716 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111111; // iC=-2113 
// vC = 14'b0000001011110001; // vC=  753 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011110; // iC=-2210 
// vC = 14'b0000001011010111; // vC=  727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b0000001000111010; // vC=  570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b0000001011010010; // vC=  722 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101101; // iC=-2131 
// vC = 14'b0000001011000000; // vC=  704 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b0000000111101001; // vC=  489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b0000001000001011; // vC=  523 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000000111101101; // vC=  493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110001; // iC=-2063 
// vC = 14'b0000000111001010; // vC=  458 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000001001011110; // vC=  606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000001011011011; // vC=  731 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000000110011111; // vC=  415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111110; // iC=-2050 
// vC = 14'b0000001000101011; // vC=  555 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101110; // iC=-2194 
// vC = 14'b0000000110001111; // vC=  399 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001000; // iC=-2040 
// vC = 14'b0000000111001111; // vC=  463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001111; // iC=-2161 
// vC = 14'b0000000111100100; // vC=  484 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b0000000111110011; // vC=  499 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b0000000111010000; // vC=  464 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010111; // iC=-2153 
// vC = 14'b0000001000000000; // vC=  512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b0000001001100110; // vC=  614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000000111011101; // vC=  477 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101001; // iC=-2199 
// vC = 14'b0000001001001110; // vC=  590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000000; // iC=-2240 
// vC = 14'b0000000110110010; // vC=  434 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b0000001001100110; // vC=  614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100001; // iC=-2207 
// vC = 14'b0000001001011101; // vC=  605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000000111010111; // vC=  471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000000110111101; // vC=  445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b0000000110011011; // vC=  411 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100100; // iC=-2204 
// vC = 14'b0000000111100010; // vC=  482 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b0000001000011000; // vC=  536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011100; // iC=-2212 
// vC = 14'b0000000110000101; // vC=  389 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010011; // iC=-2093 
// vC = 14'b0000001000000110; // vC=  518 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100100111; // iC=-2265 
// vC = 14'b0000000100101011; // vC=  299 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111111; // iC=-2113 
// vC = 14'b0000000101001001; // vC=  329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b0000000011101101; // vC=  237 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010110; // iC=-2026 
// vC = 14'b0000000110010010; // vC=  402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110100; // iC=-2124 
// vC = 14'b0000000110000000; // vC=  384 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000000011010000; // vC=  208 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011000; // iC=-2216 
// vC = 14'b0000000111000001; // vC=  449 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111010; // iC=-2246 
// vC = 14'b0000000100010101; // vC=  277 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b0000000011101111; // vC=  239 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b0000000100001000; // vC=  264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000110; // iC=-2106 
// vC = 14'b0000000100100111; // vC=  295 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101110; // iC=-2258 
// vC = 14'b0000000011110001; // vC=  241 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010010; // iC=-2222 
// vC = 14'b0000000011001101; // vC=  205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b0000000010101111; // vC=  175 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101010; // iC=-2198 
// vC = 14'b0000000001011111; // vC=   95 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110000; // iC=-2064 
// vC = 14'b0000000001011101; // vC=   93 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110111; // iC=-2249 
// vC = 14'b0000000101101011; // vC=  363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011010; // iC=-2214 
// vC = 14'b0000000010010101; // vC=  149 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000000010100010; // vC=  162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b0000000101010110; // vC=  342 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110101; // iC=-2123 
// vC = 14'b0000000101000111; // vC=  327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010010; // iC=-1966 
// vC = 14'b0000000100000001; // vC=  257 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110001; // iC=-2191 
// vC = 14'b0000000010101111; // vC=  175 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001011; // iC=-2229 
// vC = 14'b0000000010110000; // vC=  176 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001011; // iC=-1973 
// vC = 14'b0000000000010001; // vC=   17 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011101; // iC=-2147 
// vC = 14'b0000000100100000; // vC=  288 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b0000000010010011; // vC=  147 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111101; // iC=-2115 
// vC = 14'b0000000100101000; // vC=  296 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101110; // iC=-2130 
// vC = 14'b0000000011000010; // vC=  194 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000110; // iC=-2106 
// vC = 14'b1111111111001111; // vC=  -49 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100100; // iC=-1948 
// vC = 14'b0000000010010111; // vC=  151 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111000; // iC=-1928 
// vC = 14'b0000000000001110; // vC=   14 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b0000000001001111; // vC=   79 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111110; // iC=-2178 
// vC = 14'b0000000000101101; // vC=   45 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b0000000010100000; // vC=  160 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b0000000010000011; // vC=  131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b1111111111101110; // vC=  -18 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b0000000010111001; // vC=  185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111000; // iC=-2056 
// vC = 14'b0000000000001000; // vC=    8 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100000; // iC=-1952 
// vC = 14'b1111111110010101; // vC= -107 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000000000010100; // vC=   20 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011001; // iC=-2215 
// vC = 14'b0000000000001000; // vC=    8 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000111; // iC=-2105 
// vC = 14'b1111111111101011; // vC=  -21 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000000000000011; // vC=    3 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011000; // iC=-2216 
// vC = 14'b1111111111100001; // vC=  -31 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b1111111111110110; // vC=  -10 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100000; // iC=-1952 
// vC = 14'b1111111110000000; // vC= -128 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b1111111111001011; // vC=  -53 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000000001001011; // vC=   75 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110000; // iC=-2192 
// vC = 14'b1111111101000010; // vC= -190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010010; // iC=-2222 
// vC = 14'b0000000000001000; // vC=    8 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111011; // iC=-2181 
// vC = 14'b1111111110101001; // vC=  -87 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b1111111101100010; // vC= -158 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b1111111111110101; // vC=  -11 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b1111111110011011; // vC= -101 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110111; // iC=-2185 
// vC = 14'b1111111111000001; // vC=  -63 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000001; // iC=-1983 
// vC = 14'b1111111101110111; // vC= -137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001111; // iC=-2161 
// vC = 14'b0000000000010100; // vC=   20 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111100; // iC=-2116 
// vC = 14'b1111111100000100; // vC= -252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b1111111111100101; // vC=  -27 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111111; // iC=-2177 
// vC = 14'b1111111101110101; // vC= -139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b1111111011000010; // vC= -318 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b1111111011001100; // vC= -308 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111111; // iC=-1921 
// vC = 14'b1111111100001110; // vC= -242 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110101; // iC=-2187 
// vC = 14'b1111111010111111; // vC= -321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100010; // iC=-1886 
// vC = 14'b1111111101110100; // vC= -140 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010010; // iC=-2094 
// vC = 14'b1111111010110101; // vC= -331 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010101; // iC=-2091 
// vC = 14'b1111111100100001; // vC= -223 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100000; // iC=-2080 
// vC = 14'b1111111010111110; // vC= -322 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b1111111101000111; // vC= -185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b1111111001110011; // vC= -397 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101010; // iC=-2134 
// vC = 14'b1111111001110010; // vC= -398 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b1111111101001101; // vC= -179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b1111111100100011; // vC= -221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b1111111010001000; // vC= -376 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b1111111101101011; // vC= -149 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011010; // iC=-1894 
// vC = 14'b1111111101000000; // vC= -192 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101111; // iC=-1873 
// vC = 14'b1111111100011110; // vC= -226 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b1111111100000110; // vC= -250 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b1111111100001111; // vC= -241 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b1111111001111100; // vC= -388 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010110; // iC=-1898 
// vC = 14'b1111111010100000; // vC= -352 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b1111111001101000; // vC= -408 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000100; // iC=-1916 
// vC = 14'b1111111100001111; // vC= -241 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b1111111100000010; // vC= -254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b1111111010100010; // vC= -350 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b1111111000000101; // vC= -507 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b1111110111101000; // vC= -536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100010; // iC=-1886 
// vC = 14'b1111111010111010; // vC= -326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010010; // iC=-2094 
// vC = 14'b1111111001101010; // vC= -406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100111; // iC=-2073 
// vC = 14'b1111111010101000; // vC= -344 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100101; // iC=-1819 
// vC = 14'b1111111011110100; // vC= -268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111001; // iC=-1991 
// vC = 14'b1111111000010001; // vC= -495 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111101; // iC=-1923 
// vC = 14'b1111111010000110; // vC= -378 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b1111111001100011; // vC= -413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b1111110110001111; // vC= -625 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110001; // iC=-2127 
// vC = 14'b1111111000110111; // vC= -457 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000100; // iC=-1980 
// vC = 14'b1111110111111001; // vC= -519 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b1111110101111010; // vC= -646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001110; // iC=-1906 
// vC = 14'b1111110111001001; // vC= -567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b1111110111000100; // vC= -572 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011001; // iC=-2087 
// vC = 14'b1111111001110100; // vC= -396 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000011; // iC=-1789 
// vC = 14'b1111111000011011; // vC= -485 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b1111110111100111; // vC= -537 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011001; // iC=-1831 
// vC = 14'b1111110111100110; // vC= -538 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010100; // iC=-2092 
// vC = 14'b1111110110011110; // vC= -610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b1111110110001110; // vC= -626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001001; // iC=-1783 
// vC = 14'b1111110110101100; // vC= -596 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001011; // iC=-1845 
// vC = 14'b1111110101001011; // vC= -693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b1111110101001011; // vC= -693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011000; // iC=-2024 
// vC = 14'b1111111000101111; // vC= -465 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b1111110100111010; // vC= -710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b1111111001000011; // vC= -445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100101; // iC=-2011 
// vC = 14'b1111110111001000; // vC= -568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011111; // iC=-1825 
// vC = 14'b1111111000000110; // vC= -506 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011100; // iC=-1956 
// vC = 14'b1111110111011111; // vC= -545 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b1111110100010001; // vC= -751 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b1111110011111010; // vC= -774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b1111110111110100; // vC= -524 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000011; // iC=-1789 
// vC = 14'b1111110110010111; // vC= -617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101111; // iC=-1937 
// vC = 14'b1111110100000000; // vC= -768 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b1111110100111011; // vC= -709 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011010; // iC=-1894 
// vC = 14'b1111110011000001; // vC= -831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b1111110011001100; // vC= -820 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101111; // iC=-2001 
// vC = 14'b1111110111000100; // vC= -572 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011111; // iC=-1953 
// vC = 14'b1111110110011010; // vC= -614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101000; // iC=-1816 
// vC = 14'b1111110010101111; // vC= -849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101001; // iC=-1751 
// vC = 14'b1111110100001110; // vC= -754 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111100; // iC=-1796 
// vC = 14'b1111110101100101; // vC= -667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b1111110010101000; // vC= -856 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000000; // iC=-1792 
// vC = 14'b1111110011100000; // vC= -800 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b1111110100111100; // vC= -708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001100; // iC=-1972 
// vC = 14'b1111110001101110; // vC= -914 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100001; // iC=-1695 
// vC = 14'b1111110001111000; // vC= -904 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110011; // iC=-1741 
// vC = 14'b1111110010111100; // vC= -836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110100; // iC=-1932 
// vC = 14'b1111110010110011; // vC= -845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001010; // iC=-1782 
// vC = 14'b1111110100111100; // vC= -708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b1111110010000111; // vC= -889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000101; // iC=-1851 
// vC = 14'b1111110101010111; // vC= -681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101100; // iC=-1748 
// vC = 14'b1111110010100101; // vC= -859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110100; // iC=-1932 
// vC = 14'b1111110001101010; // vC= -918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101110; // iC=-1746 
// vC = 14'b1111110100010011; // vC= -749 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110000; // iC=-1936 
// vC = 14'b1111110010000100; // vC= -892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b1111110001101100; // vC= -916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111010; // iC=-1862 
// vC = 14'b1111110101000111; // vC= -697 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b1111110001010011; // vC= -941 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111000; // iC=-1672 
// vC = 14'b1111110010000001; // vC= -895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110001; // iC=-1935 
// vC = 14'b1111110000100001; // vC= -991 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010111; // iC=-1897 
// vC = 14'b1111110001100100; // vC= -924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001011; // iC=-1781 
// vC = 14'b1111110100000010; // vC= -766 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000011; // iC=-1661 
// vC = 14'b1111110010110011; // vC= -845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100111; // iC=-1881 
// vC = 14'b1111110010000110; // vC= -890 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000101; // iC=-1787 
// vC = 14'b1111110010010101; // vC= -875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101001; // iC=-1687 
// vC = 14'b1111110010001010; // vC= -886 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010111; // iC=-1833 
// vC = 14'b1111101111001001; // vC=-1079 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100100; // iC=-1884 
// vC = 14'b1111110000100010; // vC= -990 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001110; // iC=-1778 
// vC = 14'b1111110001100100; // vC= -924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100100; // iC=-1628 
// vC = 14'b1111110000101100; // vC= -980 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110000; // iC=-1616 
// vC = 14'b1111110010011100; // vC= -868 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011000; // iC=-1640 
// vC = 14'b1111110000010000; // vC=-1008 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111001; // iC=-1671 
// vC = 14'b1111110010111110; // vC= -834 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010101; // iC=-1707 
// vC = 14'b1111101110100100; // vC=-1116 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011110; // iC=-1634 
// vC = 14'b1111110010100110; // vC= -858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010110; // iC=-1898 
// vC = 14'b1111101110010100; // vC=-1132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100011; // iC=-1629 
// vC = 14'b1111101110001101; // vC=-1139 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001001; // iC=-1591 
// vC = 14'b1111110001001001; // vC= -951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110001; // iC=-1615 
// vC = 14'b1111110001100111; // vC= -921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000010; // iC=-1790 
// vC = 14'b1111101101011101; // vC=-1187 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011011; // iC=-1701 
// vC = 14'b1111110001001110; // vC= -946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b1111110000011101; // vC= -995 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001001; // iC=-1847 
// vC = 14'b1111101101111111; // vC=-1153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111101; // iC=-1667 
// vC = 14'b1111101111010101; // vC=-1067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001100; // iC=-1588 
// vC = 14'b1111101111111000; // vC=-1032 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100100; // iC=-1564 
// vC = 14'b1111110001010001; // vC= -943 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000001; // iC=-1535 
// vC = 14'b1111101111010001; // vC=-1071 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100101; // iC=-1691 
// vC = 14'b1111101101010010; // vC=-1198 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101011; // iC=-1685 
// vC = 14'b1111110000111010; // vC= -966 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000000; // iC=-1664 
// vC = 14'b1111110000110100; // vC= -972 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010111; // iC=-1577 
// vC = 14'b1111101110110110; // vC=-1098 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011011; // iC=-1509 
// vC = 14'b1111101110110101; // vC=-1099 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110011; // iC=-1549 
// vC = 14'b1111101101111011; // vC=-1157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110111; // iC=-1673 
// vC = 14'b1111101111010010; // vC=-1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111100; // iC=-1796 
// vC = 14'b1111101101001100; // vC=-1204 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011100; // iC=-1636 
// vC = 14'b1111101101111000; // vC=-1160 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110001; // iC=-1615 
// vC = 14'b1111110000000111; // vC=-1017 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011100; // iC=-1636 
// vC = 14'b1111101110001111; // vC=-1137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b1111101110010010; // vC=-1134 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001101; // iC=-1651 
// vC = 14'b1111101100100000; // vC=-1248 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101001; // iC=-1751 
// vC = 14'b1111101100011111; // vC=-1249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010101; // iC=-1771 
// vC = 14'b1111101011111101; // vC=-1283 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100001; // iC=-1503 
// vC = 14'b1111101100011001; // vC=-1255 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100101; // iC=-1563 
// vC = 14'b1111101100101111; // vC=-1233 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101011; // iC=-1621 
// vC = 14'b1111101111101010; // vC=-1046 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010111; // iC=-1641 
// vC = 14'b1111101011011101; // vC=-1315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100000; // iC=-1440 
// vC = 14'b1111101111000001; // vC=-1087 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101111; // iC=-1489 
// vC = 14'b1111101111010110; // vC=-1066 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000001; // iC=-1471 
// vC = 14'b1111101011011000; // vC=-1320 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001110; // iC=-1458 
// vC = 14'b1111101100100101; // vC=-1243 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100100; // iC=-1628 
// vC = 14'b1111101010001101; // vC=-1395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110110; // iC=-1546 
// vC = 14'b1111101110011001; // vC=-1127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010100; // iC=-1452 
// vC = 14'b1111101101111111; // vC=-1153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110000; // iC=-1424 
// vC = 14'b1111101011011110; // vC=-1314 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000000; // iC=-1664 
// vC = 14'b1111101010100101; // vC=-1371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110110; // iC=-1482 
// vC = 14'b1111101011010111; // vC=-1321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011110; // iC=-1506 
// vC = 14'b1111101100011111; // vC=-1249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000011; // iC=-1533 
// vC = 14'b1111101011000000; // vC=-1344 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111100; // iC=-1540 
// vC = 14'b1111101100111100; // vC=-1220 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011110; // iC=-1570 
// vC = 14'b1111101101110100; // vC=-1164 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110110; // iC=-1610 
// vC = 14'b1111101100000101; // vC=-1275 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101011; // iC=-1557 
// vC = 14'b1111101011000001; // vC=-1343 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011000; // iC=-1448 
// vC = 14'b1111101001000001; // vC=-1471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101001; // iC=-1623 
// vC = 14'b1111101100001111; // vC=-1265 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100111; // iC=-1625 
// vC = 14'b1111101001001101; // vC=-1459 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011111; // iC=-1441 
// vC = 14'b1111101001110011; // vC=-1421 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010110; // iC=-1578 
// vC = 14'b1111101001001001; // vC=-1463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111001; // iC=-1543 
// vC = 14'b1111101001101001; // vC=-1431 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111100; // iC=-1476 
// vC = 14'b1111101001100100; // vC=-1436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111100; // iC=-1348 
// vC = 14'b1111101010011010; // vC=-1382 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001010; // iC=-1590 
// vC = 14'b1111101000100110; // vC=-1498 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010111; // iC=-1513 
// vC = 14'b1111101011101000; // vC=-1304 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101100; // iC=-1492 
// vC = 14'b1111101100000111; // vC=-1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101011; // iC=-1365 
// vC = 14'b1111101100110110; // vC=-1226 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101111; // iC=-1553 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100110; // iC=-1370 
// vC = 14'b1111101100011101; // vC=-1251 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110100; // iC=-1292 
// vC = 14'b1111101000010101; // vC=-1515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110110; // iC=-1354 
// vC = 14'b1111101001110101; // vC=-1419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001101; // iC=-1459 
// vC = 14'b1111101010011111; // vC=-1377 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101100; // iC=-1364 
// vC = 14'b1111100111010110; // vC=-1578 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101010; // iC=-1494 
// vC = 14'b1111101011010100; // vC=-1324 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110101; // iC=-1355 
// vC = 14'b1111101001101011; // vC=-1429 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000000; // iC=-1472 
// vC = 14'b1111100111011001; // vC=-1575 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110011; // iC=-1549 
// vC = 14'b1111101000010101; // vC=-1515 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000110; // iC=-1530 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111010; // iC=-1478 
// vC = 14'b1111101010011111; // vC=-1377 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010000; // iC=-1392 
// vC = 14'b1111101001011011; // vC=-1445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010011; // iC=-1261 
// vC = 14'b1111101001110001; // vC=-1423 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001100; // iC=-1524 
// vC = 14'b1111101000110101; // vC=-1483 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000100; // iC=-1404 
// vC = 14'b1111101000010010; // vC=-1518 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110101; // iC=-1483 
// vC = 14'b1111100111001101; // vC=-1587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111100; // iC=-1476 
// vC = 14'b1111101000110111; // vC=-1481 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111011; // iC=-1221 
// vC = 14'b1111100110101010; // vC=-1622 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011110; // iC=-1250 
// vC = 14'b1111101000111001; // vC=-1479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000011; // iC=-1469 
// vC = 14'b1111101010101110; // vC=-1362 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001110; // iC=-1202 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111000; // iC=-1480 
// vC = 14'b1111100110011011; // vC=-1637 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111101; // iC=-1411 
// vC = 14'b1111101000011111; // vC=-1505 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101000; // iC=-1368 
// vC = 14'b1111100110110111; // vC=-1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110010; // iC=-1230 
// vC = 14'b1111101000011101; // vC=-1507 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111011; // iC=-1221 
// vC = 14'b1111101000001111; // vC=-1521 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000111; // iC=-1273 
// vC = 14'b1111101001111000; // vC=-1416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101110; // iC=-1362 
// vC = 14'b1111101000110010; // vC=-1486 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101100; // iC=-1300 
// vC = 14'b1111100111101111; // vC=-1553 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100101; // iC=-1179 
// vC = 14'b1111101000001001; // vC=-1527 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110001; // iC=-1231 
// vC = 14'b1111101001011001; // vC=-1447 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111001; // iC=-1159 
// vC = 14'b1111101001110100; // vC=-1420 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001111; // iC=-1265 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000110; // iC=-1210 
// vC = 14'b1111100111000100; // vC=-1596 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100010; // iC=-1310 
// vC = 14'b1111100101111001; // vC=-1671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010110; // iC=-1258 
// vC = 14'b1111101000010011; // vC=-1517 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100111; // iC=-1369 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011110; // iC=-1314 
// vC = 14'b1111101000111101; // vC=-1475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000000; // iC=-1216 
// vC = 14'b1111100111101000; // vC=-1560 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100110; // iC=-1114 
// vC = 14'b1111101001001001; // vC=-1463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111000; // iC=-1288 
// vC = 14'b1111100101100111; // vC=-1689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000110; // iC=-1146 
// vC = 14'b1111100100101010; // vC=-1750 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011011; // iC=-1253 
// vC = 14'b1111100110010000; // vC=-1648 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111011; // iC=-1349 
// vC = 14'b1111100110110100; // vC=-1612 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010011; // iC=-1197 
// vC = 14'b1111100111110001; // vC=-1551 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111000; // iC=-1352 
// vC = 14'b1111100101011101; // vC=-1699 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111110; // iC=-1282 
// vC = 14'b1111100101010001; // vC=-1711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111001; // iC=-1351 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010010; // iC=-1070 
// vC = 14'b1111101000000110; // vC=-1530 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101111; // iC=-1233 
// vC = 14'b1111100100001100; // vC=-1780 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000110; // iC=-1146 
// vC = 14'b1111100011101010; // vC=-1814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111011; // iC=-1221 
// vC = 14'b1111100111101110; // vC=-1554 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001001; // iC=-1015 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100100; // iC=-1244 
// vC = 14'b1111100111110110; // vC=-1546 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001101; // iC=-1203 
// vC = 14'b1111100111111111; // vC=-1537 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101110; // iC=-1170 
// vC = 14'b1111100111010100; // vC=-1580 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011110; // iC=-1186 
// vC = 14'b1111100110010011; // vC=-1645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111010; // iC=-1158 
// vC = 14'b1111100111001000; // vC=-1592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010111; // iC=-1001 
// vC = 14'b1111100111100000; // vC=-1568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111000; // iC=-1160 
// vC = 14'b1111100101110100; // vC=-1676 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010100; // iC=-1068 
// vC = 14'b1111100110100001; // vC=-1631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000010; // iC=-1214 
// vC = 14'b1111100100111011; // vC=-1733 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010101; // iC=-1259 
// vC = 14'b1111100101000011; // vC=-1725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110011; // iC=-1229 
// vC = 14'b1111100110011001; // vC=-1639 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001110; // iC= -946 
// vC = 14'b1111100100101010; // vC=-1750 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001110; // iC= -946 
// vC = 14'b1111100100100110; // vC=-1754 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001111; // iC= -945 
// vC = 14'b1111100011101101; // vC=-1811 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110111; // iC=-1161 
// vC = 14'b1111100011110111; // vC=-1801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000010; // iC=-1150 
// vC = 14'b1111100011100011; // vC=-1821 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100011; // iC= -925 
// vC = 14'b1111100010011010; // vC=-1894 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000000; // iC=-1024 
// vC = 14'b1111100100000101; // vC=-1787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110001; // iC= -975 
// vC = 14'b1111100100011011; // vC=-1765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011010; // iC=-1190 
// vC = 14'b1111100101111100; // vC=-1668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010010; // iC=-1198 
// vC = 14'b1111100110010011; // vC=-1645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011100; // iC= -932 
// vC = 14'b1111100010001001; // vC=-1911 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000010; // iC= -894 
// vC = 14'b1111100010001110; // vC=-1906 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100010; // iC=-1182 
// vC = 14'b1111100011010101; // vC=-1835 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001000; // iC=-1080 
// vC = 14'b1111100110000110; // vC=-1658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010100; // iC=-1068 
// vC = 14'b1111100010011010; // vC=-1894 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001000; // iC=-1080 
// vC = 14'b1111100010100000; // vC=-1888 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001101; // iC= -947 
// vC = 14'b1111100001011101; // vC=-1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000000; // iC=-1152 
// vC = 14'b1111100100101110; // vC=-1746 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010001; // iC= -943 
// vC = 14'b1111100011001011; // vC=-1845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010110; // iC=-1066 
// vC = 14'b1111100011111001; // vC=-1799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000000; // iC= -896 
// vC = 14'b1111100001011100; // vC=-1956 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101101; // iC= -851 
// vC = 14'b1111100001000111; // vC=-1977 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100100; // iC= -988 
// vC = 14'b1111100010111101; // vC=-1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111110; // iC=-1090 
// vC = 14'b1111100101100110; // vC=-1690 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001001; // iC= -887 
// vC = 14'b1111100010101010; // vC=-1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111100; // iC= -964 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111000; // iC= -904 
// vC = 14'b1111100001011001; // vC=-1959 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011000; // iC= -936 
// vC = 14'b1111100010100000; // vC=-1888 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110100; // iC= -972 
// vC = 14'b1111100101110000; // vC=-1680 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011010; // iC= -870 
// vC = 14'b1111100001111111; // vC=-1921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111101; // iC= -963 
// vC = 14'b1111100001001111; // vC=-1969 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101100; // iC= -980 
// vC = 14'b1111100010101101; // vC=-1875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000010; // iC=-1022 
// vC = 14'b1111100010010010; // vC=-1902 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111011; // iC= -773 
// vC = 14'b1111100010010100; // vC=-1900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101101; // iC= -723 
// vC = 14'b1111100000101001; // vC=-2007 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100001; // iC= -735 
// vC = 14'b1111100000100000; // vC=-2016 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011001; // iC= -807 
// vC = 14'b1111100011000111; // vC=-1849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101101; // iC= -851 
// vC = 14'b1111100100101110; // vC=-1746 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011101; // iC= -867 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001010; // iC= -950 
// vC = 14'b1111100010010011; // vC=-1901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010111; // iC= -745 
// vC = 14'b1111100000011001; // vC=-2023 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001011; // iC= -821 
// vC = 14'b1111100001000000; // vC=-1984 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111101; // iC= -899 
// vC = 14'b1111100001001000; // vC=-1976 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111011; // iC= -901 
// vC = 14'b1111100010001011; // vC=-1909 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001110; // iC= -754 
// vC = 14'b1111011111111110; // vC=-2050 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010110; // iC= -746 
// vC = 14'b1111011111111000; // vC=-2056 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110011; // iC= -717 
// vC = 14'b1111100011101111; // vC=-1809 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100010; // iC= -734 
// vC = 14'b1111100011101100; // vC=-1812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001100; // iC= -692 
// vC = 14'b1111011111110010; // vC=-2062 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100001; // iC= -863 
// vC = 14'b1111100001100011; // vC=-1949 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110001; // iC= -719 
// vC = 14'b1111100000100111; // vC=-2009 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101101; // iC= -659 
// vC = 14'b1111100001000111; // vC=-1977 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001010; // iC= -630 
// vC = 14'b1111100010000001; // vC=-1919 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000111; // iC= -761 
// vC = 14'b1111100001011101; // vC=-1955 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101010; // iC= -790 
// vC = 14'b1111100010100111; // vC=-1881 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001001; // iC= -631 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111110; // iC= -898 
// vC = 14'b1111100001000000; // vC=-1984 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100111; // iC= -793 
// vC = 14'b1111100011101100; // vC=-1812 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001000; // iC= -824 
// vC = 14'b1111100000100111; // vC=-2009 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000000; // iC= -768 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100111; // iC= -665 
// vC = 14'b1111011111101011; // vC=-2069 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001110; // iC= -626 
// vC = 14'b1111100010000100; // vC=-1916 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000111; // iC= -633 
// vC = 14'b1111011111000010; // vC=-2110 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110100; // iC= -588 
// vC = 14'b1111100001011011; // vC=-1957 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010011; // iC= -685 
// vC = 14'b1111011111100110; // vC=-2074 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111001; // iC= -839 
// vC = 14'b1111011111001111; // vC=-2097 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101000; // iC= -728 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011011; // iC= -549 
// vC = 14'b1111011111111000; // vC=-2056 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011000; // iC= -552 
// vC = 14'b1111100011101110; // vC=-1810 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001001; // iC= -567 
// vC = 14'b1111100011110000; // vC=-1808 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001001; // iC= -631 
// vC = 14'b1111100011110000; // vC=-1808 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000100; // iC= -700 
// vC = 14'b1111011111001101; // vC=-2099 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101011; // iC= -597 
// vC = 14'b1111011110111000; // vC=-2120 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011011; // iC= -549 
// vC = 14'b1111100011101001; // vC=-1815 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011100; // iC= -740 
// vC = 14'b1111011111000110; // vC=-2106 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100101; // iC= -603 
// vC = 14'b1111011110101000; // vC=-2136 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111010; // iC= -582 
// vC = 14'b1111100000110010; // vC=-1998 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111100; // iC= -452 
// vC = 14'b1111100000110000; // vC=-2000 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110000; // iC= -464 
// vC = 14'b1111100001110110; // vC=-1930 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011110; // iC= -674 
// vC = 14'b1111100000010011; // vC=-2029 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100100; // iC= -412 
// vC = 14'b1111100000100011; // vC=-2013 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011001; // iC= -359 
// vC = 14'b1111011111110110; // vC=-2058 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000011; // iC= -573 
// vC = 14'b1111011111111011; // vC=-2053 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110101; // iC= -331 
// vC = 14'b1111100011010101; // vC=-1835 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110001; // iC= -591 
// vC = 14'b1111100000000001; // vC=-2047 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101101; // iC= -531 
// vC = 14'b1111011110111101; // vC=-2115 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111111; // iC= -321 
// vC = 14'b1111100000100010; // vC=-2014 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011111010; // iC= -262 
// vC = 14'b1111100000110000; // vC=-2000 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001100; // iC= -372 
// vC = 14'b1111011110001010; // vC=-2166 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001111; // iC= -241 
// vC = 14'b1111100000111000; // vC=-1992 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001001; // iC= -311 
// vC = 14'b1111011111010111; // vC=-2089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011100111; // iC= -281 
// vC = 14'b1111100001110001; // vC=-1935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111110; // iC= -194 
// vC = 14'b1111100000000000; // vC=-2048 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111011; // iC= -389 
// vC = 14'b1111100010100001; // vC=-1887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101011110; // iC= -162 
// vC = 14'b1111100001001110; // vC=-1970 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000111; // iC= -121 
// vC = 14'b1111011111011011; // vC=-2085 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011111; // iC= -353 
// vC = 14'b1111100000010101; // vC=-2027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011011; // iC= -293 
// vC = 14'b1111011111010100; // vC=-2092 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100000; // iC= -224 
// vC = 14'b1111100001001111; // vC=-1969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010011111; // iC= -353 
// vC = 14'b1111011110000011; // vC=-2173 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101011001; // iC= -167 
// vC = 14'b1111011111111101; // vC=-2051 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001111; // iC= -305 
// vC = 14'b1111011110101000; // vC=-2136 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110001110; // iC= -114 
// vC = 14'b1111100001101011; // vC=-1941 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000000; // iC=  -64 
// vC = 14'b1111011111010101; // vC=-2091 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000110; // iC= -186 
// vC = 14'b1111100000100111; // vC=-2009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001110; // iC=  -50 
// vC = 14'b1111011110010011; // vC=-2157 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101110010; // iC= -142 
// vC = 14'b1111100001101111; // vC=-1937 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110001; // iC= -207 
// vC = 14'b1111100000110101; // vC=-1995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011110; // iC=  -98 
// vC = 14'b1111011110001110; // vC=-2162 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000001; // iC=  -63 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100010; // iC=  -94 
// vC = 14'b1111100001001000; // vC=-1976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100111; // iC=  103 
// vC = 14'b1111011110010100; // vC=-2156 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000100; // iC=  132 
// vC = 14'b1111011110011100; // vC=-2148 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101000; // iC=   40 
// vC = 14'b1111011110011100; // vC=-2148 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000111; // iC=  135 
// vC = 14'b1111011111110110; // vC=-2058 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001100; // iC=  140 
// vC = 14'b1111011110101100; // vC=-2132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100001; // iC=  289 
// vC = 14'b1111100010101000; // vC=-1880 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010100; // iC=  148 
// vC = 14'b1111100010111110; // vC=-1858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110111; // iC=  247 
// vC = 14'b1111100000000100; // vC=-2044 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001110; // iC=  206 
// vC = 14'b1111011110000111; // vC=-2169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101111; // iC=  367 
// vC = 14'b1111011110011011; // vC=-2149 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100000; // iC=  288 
// vC = 14'b1111100000000111; // vC=-2041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110000; // iC=  304 
// vC = 14'b1111100010000111; // vC=-1913 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110000; // iC=  176 
// vC = 14'b1111100010101010; // vC=-1878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110101; // iC=  181 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100101; // iC=  229 
// vC = 14'b1111100001011001; // vC=-1959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110111; // iC=  439 
// vC = 14'b1111100000010010; // vC=-2030 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010101; // iC=  341 
// vC = 14'b1111011110101010; // vC=-2134 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111010; // iC=  314 
// vC = 14'b1111100010101000; // vC=-1880 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001111; // iC=  399 
// vC = 14'b1111100000111001; // vC=-1991 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010011; // iC=  531 
// vC = 14'b1111100000101101; // vC=-2003 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001111; // iC=  591 
// vC = 14'b1111100011100001; // vC=-1823 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010100; // iC=  532 
// vC = 14'b1111100001001100; // vC=-1972 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001011; // iC=  523 
// vC = 14'b1111100011010011; // vC=-1837 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100111; // iC=  551 
// vC = 14'b1111100000010100; // vC=-2028 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101000; // iC=  616 
// vC = 14'b1111100010011001; // vC=-1895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101011; // iC=  619 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111010; // iC=  506 
// vC = 14'b1111011111001100; // vC=-2100 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011101; // iC=  605 
// vC = 14'b1111100001011110; // vC=-1954 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000001; // iC=  513 
// vC = 14'b1111100010011011; // vC=-1893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100110; // iC=  614 
// vC = 14'b1111100010001001; // vC=-1911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110011; // iC=  563 
// vC = 14'b1111011111001111; // vC=-2097 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010111; // iC=  791 
// vC = 14'b1111100011101101; // vC=-1811 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011101; // iC=  797 
// vC = 14'b1111100011000001; // vC=-1855 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000110; // iC=  710 
// vC = 14'b1111100000011011; // vC=-2021 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000000; // iC=  704 
// vC = 14'b1111100010111101; // vC=-1859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101001; // iC=  745 
// vC = 14'b1111011111100110; // vC=-2074 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000001; // iC=  833 
// vC = 14'b1111100010111101; // vC=-1859 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001100; // iC=  716 
// vC = 14'b1111100010000101; // vC=-1915 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110010; // iC= 1010 
// vC = 14'b1111100011111110; // vC=-1794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000111; // iC=  903 
// vC = 14'b1111100001011100; // vC=-1956 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011100; // iC=  796 
// vC = 14'b1111100000001001; // vC=-2039 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101000; // iC= 1000 
// vC = 14'b1111100001010111; // vC=-1961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100110; // iC=  998 
// vC = 14'b1111100011110111; // vC=-1801 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101001; // iC= 1001 
// vC = 14'b1111100100100100; // vC=-1756 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010011; // iC= 1171 
// vC = 14'b1111100011100101; // vC=-1819 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110100; // iC= 1140 
// vC = 14'b1111100000001100; // vC=-2036 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001001; // iC=  969 
// vC = 14'b1111100010101000; // vC=-1880 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011100; // iC=  988 
// vC = 14'b1111100011001100; // vC=-1844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101000; // iC= 1000 
// vC = 14'b1111100000001101; // vC=-2035 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100111; // iC=  999 
// vC = 14'b1111100010111000; // vC=-1864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111110; // iC= 1086 
// vC = 14'b1111100001110000; // vC=-1936 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000100; // iC= 1284 
// vC = 14'b1111100011100101; // vC=-1819 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010000; // iC= 1104 
// vC = 14'b1111100010001001; // vC=-1911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110101; // iC= 1205 
// vC = 14'b1111100000100010; // vC=-2014 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101010; // iC= 1066 
// vC = 14'b1111100001100100; // vC=-1948 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100111; // iC= 1319 
// vC = 14'b1111100011011110; // vC=-1826 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010110; // iC= 1174 
// vC = 14'b1111100000101111; // vC=-2001 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010110; // iC= 1238 
// vC = 14'b1111100100001011; // vC=-1781 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011000; // iC= 1368 
// vC = 14'b1111100100011011; // vC=-1765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000101; // iC= 1477 
// vC = 14'b1111100101011011; // vC=-1701 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101001; // iC= 1193 
// vC = 14'b1111100011110011; // vC=-1805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010100; // iC= 1236 
// vC = 14'b1111100011100110; // vC=-1818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000011; // iC= 1411 
// vC = 14'b1111100001101110; // vC=-1938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101110; // iC= 1454 
// vC = 14'b1111100101110110; // vC=-1674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011001; // iC= 1369 
// vC = 14'b1111100001111111; // vC=-1921 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000001; // iC= 1281 
// vC = 14'b1111100101111111; // vC=-1665 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111111; // iC= 1599 
// vC = 14'b1111100010110100; // vC=-1868 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000000; // iC= 1536 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010111; // iC= 1367 
// vC = 14'b1111100101011101; // vC=-1699 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000000; // iC= 1344 
// vC = 14'b1111100101001000; // vC=-1720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010110; // iC= 1558 
// vC = 14'b1111100110111100; // vC=-1604 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100001; // iC= 1569 
// vC = 14'b1111100010011100; // vC=-1892 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110011; // iC= 1651 
// vC = 14'b1111100110100011; // vC=-1629 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001011; // iC= 1675 
// vC = 14'b1111100110110010; // vC=-1614 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101100; // iC= 1644 
// vC = 14'b1111100100010010; // vC=-1774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000001; // iC= 1601 
// vC = 14'b1111100100010001; // vC=-1775 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110010; // iC= 1714 
// vC = 14'b1111100110110010; // vC=-1614 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111110; // iC= 1726 
// vC = 14'b1111100011110000; // vC=-1808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101001; // iC= 1769 
// vC = 14'b1111100011101001; // vC=-1815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000001; // iC= 1537 
// vC = 14'b1111100110110111; // vC=-1609 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111000; // iC= 1784 
// vC = 14'b1111100110011111; // vC=-1633 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101111; // iC= 1711 
// vC = 14'b1111100111100110; // vC=-1562 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001100; // iC= 1740 
// vC = 14'b1111100011011110; // vC=-1826 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100101; // iC= 1573 
// vC = 14'b1111100110001100; // vC=-1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010001; // iC= 1553 
// vC = 14'b1111100111111111; // vC=-1537 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001111; // iC= 1871 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b1111100101011011; // vC=-1701 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b1111100110111001; // vC=-1607 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010110; // iC= 1686 
// vC = 14'b1111100101000101; // vC=-1723 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010111; // iC= 1751 
// vC = 14'b1111100101101100; // vC=-1684 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000110; // iC= 1670 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100001; // iC= 1825 
// vC = 14'b1111100110011000; // vC=-1640 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010111; // iC= 1687 
// vC = 14'b1111101001001100; // vC=-1460 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110000; // iC= 1648 
// vC = 14'b1111100111101101; // vC=-1555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b1111100110101001; // vC=-1623 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b1111100110011101; // vC=-1635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b1111100111100011; // vC=-1565 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011011; // iC= 1947 
// vC = 14'b1111100111000011; // vC=-1597 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111110; // iC= 1726 
// vC = 14'b1111100110101101; // vC=-1619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001000; // iC= 1800 
// vC = 14'b1111100110010011; // vC=-1645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101101; // iC= 1709 
// vC = 14'b1111101000000101; // vC=-1531 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101111; // iC= 1839 
// vC = 14'b1111101001110011; // vC=-1421 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b1111101001010100; // vC=-1452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010101; // iC= 2005 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b1111101000000000; // vC=-1536 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110100; // iC= 1844 
// vC = 14'b1111100111000100; // vC=-1596 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110101; // iC= 2037 
// vC = 14'b1111101000000111; // vC=-1529 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100100; // iC= 1828 
// vC = 14'b1111101010001111; // vC=-1393 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b1111101011000010; // vC=-1342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110110; // iC= 1782 
// vC = 14'b1111101011110011; // vC=-1293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b1111101011011010; // vC=-1318 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010000; // iC= 2000 
// vC = 14'b1111101011000100; // vC=-1340 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111101000101000; // vC=-1496 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b1111101001100100; // vC=-1436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b1111101011101010; // vC=-1302 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110111; // iC= 1847 
// vC = 14'b1111101011101101; // vC=-1299 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111101011010000; // vC=-1328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001000; // iC= 2120 
// vC = 14'b1111101000011111; // vC=-1505 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000001; // iC= 1921 
// vC = 14'b1111101001010011; // vC=-1453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000010; // iC= 2114 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010101; // iC= 1877 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b1111101011001001; // vC=-1335 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000001; // iC= 2049 
// vC = 14'b1111101011100101; // vC=-1307 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101000; // iC= 2024 
// vC = 14'b1111101101000110; // vC=-1210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010110; // iC= 2134 
// vC = 14'b1111101001001111; // vC=-1457 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000100; // iC= 2116 
// vC = 14'b1111101101111000; // vC=-1160 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011110; // iC= 2078 
// vC = 14'b1111101010000110; // vC=-1402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100000; // iC= 1888 
// vC = 14'b1111101011010110; // vC=-1322 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000000; // iC= 2048 
// vC = 14'b1111101011101111; // vC=-1297 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111101; // iC= 2109 
// vC = 14'b1111101100101111; // vC=-1233 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111101100011111; // vC=-1249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110000; // iC= 2096 
// vC = 14'b1111101110011110; // vC=-1122 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b1111101010111110; // vC=-1346 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011011; // iC= 2075 
// vC = 14'b1111101110011100; // vC=-1124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b1111101100110010; // vC=-1230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100011; // iC= 2083 
// vC = 14'b1111101111001000; // vC=-1080 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011111; // iC= 2079 
// vC = 14'b1111101100011100; // vC=-1252 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001001; // iC= 2185 
// vC = 14'b1111101111101101; // vC=-1043 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111110; // iC= 1982 
// vC = 14'b1111101100001001; // vC=-1271 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b1111101111101001; // vC=-1047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111101110010001; // vC=-1135 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111111; // iC= 2111 
// vC = 14'b1111101100000111; // vC=-1273 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b1111101011100010; // vC=-1310 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110010; // iC= 1970 
// vC = 14'b1111101110110010; // vC=-1102 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b1111101100101100; // vC=-1236 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110001; // iC= 2097 
// vC = 14'b1111101110111100; // vC=-1092 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111110000001000; // vC=-1016 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b1111101101110010; // vC=-1166 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000011; // iC= 2179 
// vC = 14'b1111101101000101; // vC=-1211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111100; // iC= 1980 
// vC = 14'b1111101100101000; // vC=-1240 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b1111101110101100; // vC=-1108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b1111101101110110; // vC=-1162 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011110; // iC= 2078 
// vC = 14'b1111110000101001; // vC= -983 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111101; // iC= 2173 
// vC = 14'b1111101101000001; // vC=-1215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110001; // iC= 1969 
// vC = 14'b1111101101110111; // vC=-1161 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b1111101111110101; // vC=-1035 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b1111110001000011; // vC= -957 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111100; // iC= 2044 
// vC = 14'b1111110010000010; // vC= -894 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b1111110000110111; // vC= -969 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101011; // iC= 2155 
// vC = 14'b1111101110010000; // vC=-1136 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b1111110010111010; // vC= -838 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000001; // iC= 2049 
// vC = 14'b1111101110111001; // vC=-1095 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b1111101110101001; // vC=-1111 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101011; // iC= 2219 
// vC = 14'b1111110011010010; // vC= -814 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101101; // iC= 2157 
// vC = 14'b1111110001101000; // vC= -920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b1111110010010001; // vC= -879 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110100; // iC= 1972 
// vC = 14'b1111110010110010; // vC= -846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b1111110001001001; // vC= -951 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b1111110000000101; // vC=-1019 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011111; // iC= 2143 
// vC = 14'b1111110000001000; // vC=-1016 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b1111110011010100; // vC= -812 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100111; // iC= 2023 
// vC = 14'b1111110011011000; // vC= -808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b1111110100100000; // vC= -736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100010; // iC= 2210 
// vC = 14'b1111110011011111; // vC= -801 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101000; // iC= 2152 
// vC = 14'b1111110011110110; // vC= -778 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000010; // iC= 2242 
// vC = 14'b1111110001111101; // vC= -899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101001; // iC= 2153 
// vC = 14'b1111110011000010; // vC= -830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001010; // iC= 1994 
// vC = 14'b1111110011100001; // vC= -799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b1111110101100011; // vC= -669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b1111110001000001; // vC= -959 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110000; // iC= 2096 
// vC = 14'b1111110100011110; // vC= -738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101001; // iC= 2217 
// vC = 14'b1111110011110010; // vC= -782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100011; // iC= 2211 
// vC = 14'b1111110100010000; // vC= -752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110000; // iC= 2032 
// vC = 14'b1111110010100110; // vC= -858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001111; // iC= 2191 
// vC = 14'b1111110110010100; // vC= -620 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111011; // iC= 2235 
// vC = 14'b1111110101110111; // vC= -649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011111; // iC= 2079 
// vC = 14'b1111110101011000; // vC= -680 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110000; // iC= 2224 
// vC = 14'b1111110110100000; // vC= -608 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b1111110011101110; // vC= -786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000011; // iC= 2243 
// vC = 14'b1111110011111110; // vC= -770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110100; // iC= 2100 
// vC = 14'b1111110011011111; // vC= -801 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011111; // iC= 2079 
// vC = 14'b1111110010101000; // vC= -856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101110; // iC= 2158 
// vC = 14'b1111110111000111; // vC= -569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111100; // iC= 2108 
// vC = 14'b1111110101110111; // vC= -649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111110010111100; // vC= -836 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110100; // iC= 2164 
// vC = 14'b1111110100000110; // vC= -762 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100100; // iC= 2212 
// vC = 14'b1111110011100100; // vC= -796 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111110; // iC= 2174 
// vC = 14'b1111110110110100; // vC= -588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111110111000111; // vC= -569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111111; // iC= 1983 
// vC = 14'b1111110110101110; // vC= -594 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b1111110111010111; // vC= -553 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111111; // iC= 2111 
// vC = 14'b1111110110010001; // vC= -623 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100000; // iC= 2144 
// vC = 14'b1111110100100010; // vC= -734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111110101010111; // vC= -681 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010010; // iC= 2130 
// vC = 14'b1111110101110011; // vC= -653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111110111010101; // vC= -555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110011; // iC= 2163 
// vC = 14'b1111111001001010; // vC= -438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100011; // iC= 2147 
// vC = 14'b1111110110101110; // vC= -594 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100011; // iC= 2211 
// vC = 14'b1111110101001100; // vC= -692 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b1111111001111101; // vC= -387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b1111110111010100; // vC= -556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010010; // iC= 2066 
// vC = 14'b1111110101110111; // vC= -649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010000; // iC= 2256 
// vC = 14'b1111111000110011; // vC= -461 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010101; // iC= 2069 
// vC = 14'b1111111001110100; // vC= -396 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011011110; // iC= 2270 
// vC = 14'b1111110111111111; // vC= -513 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b1111111010011111; // vC= -353 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111111011000101; // vC= -315 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000010; // iC= 2114 
// vC = 14'b1111111010101001; // vC= -343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100100; // iC= 2148 
// vC = 14'b1111110110100001; // vC= -607 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010000; // iC= 2256 
// vC = 14'b1111111011010110; // vC= -298 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010111; // iC= 2199 
// vC = 14'b1111111000011110; // vC= -482 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010000; // iC= 2000 
// vC = 14'b1111111001000011; // vC= -445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100011; // iC= 2211 
// vC = 14'b1111111000010100; // vC= -492 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000111; // iC= 2247 
// vC = 14'b1111111011100101; // vC= -283 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110111; // iC= 2231 
// vC = 14'b1111111010010011; // vC= -365 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000010; // iC= 2178 
// vC = 14'b1111111011000100; // vC= -316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011010; // iC= 2202 
// vC = 14'b1111111010111000; // vC= -328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010001; // iC= 2065 
// vC = 14'b1111111100100101; // vC= -219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111010; // iC= 2170 
// vC = 14'b1111111100000100; // vC= -252 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101111; // iC= 2159 
// vC = 14'b1111111100110011; // vC= -205 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100000; // iC= 2080 
// vC = 14'b1111111001111101; // vC= -387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b1111111001001101; // vC= -435 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101110; // iC= 2158 
// vC = 14'b1111111100000100; // vC= -252 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b1111111100000011; // vC= -253 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b1111111101001111; // vC= -177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b1111111101110011; // vC= -141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001110; // iC= 2190 
// vC = 14'b1111111101111100; // vC= -132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110001; // iC= 2161 
// vC = 14'b1111111110000000; // vC= -128 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011010; // iC= 2202 
// vC = 14'b1111111101010110; // vC= -170 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111111001010110; // vC= -426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010000; // iC= 2000 
// vC = 14'b1111111011100110; // vC= -282 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010010; // iC= 2194 
// vC = 14'b1111111010010010; // vC= -366 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100101; // iC= 2149 
// vC = 14'b1111111011011110; // vC= -290 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010101; // iC= 2261 
// vC = 14'b1111111110101101; // vC=  -83 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110101; // iC= 2037 
// vC = 14'b1111111100000110; // vC= -250 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000111; // iC= 2247 
// vC = 14'b1111111010001001; // vC= -375 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000101; // iC= 2053 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b1111111010110001; // vC= -335 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010111; // iC= 2199 
// vC = 14'b1111111101010011; // vC= -173 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100010; // iC= 2018 
// vC = 14'b1111111100111101; // vC= -195 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000010; // iC= 1986 
// vC = 14'b1111111110001000; // vC= -120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111110; // iC= 2046 
// vC = 14'b0000000000000110; // vC=    6 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b1111111100101101; // vC= -211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111011; // iC= 2107 
// vC = 14'b1111111100000001; // vC= -255 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100011; // iC= 2083 
// vC = 14'b1111111110101011; // vC=  -85 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101000; // iC= 2152 
// vC = 14'b0000000000000110; // vC=    6 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111011; // iC= 2171 
// vC = 14'b1111111011101101; // vC= -275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b1111111100101000; // vC= -216 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010001; // iC= 2129 
// vC = 14'b1111111100111101; // vC= -195 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110011; // iC= 2099 
// vC = 14'b1111111110000001; // vC= -127 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011011; // iC= 2203 
// vC = 14'b1111111100011011; // vC= -229 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101000; // iC= 2216 
// vC = 14'b1111111111011111; // vC=  -33 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101101; // iC= 2157 
// vC = 14'b1111111111000001; // vC=  -63 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111111100101011; // vC= -213 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111100; // iC= 2236 
// vC = 14'b0000000001011110; // vC=   94 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001010; // iC= 2186 
// vC = 14'b0000000000001000; // vC=    8 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b0000000000011110; // vC=   30 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110000; // iC= 2160 
// vC = 14'b0000000001001111; // vC=   79 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101100; // iC= 2156 
// vC = 14'b1111111110101100; // vC=  -84 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001100; // iC= 2060 
// vC = 14'b0000000000100000; // vC=   32 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111100; // iC= 2044 
// vC = 14'b1111111110010011; // vC= -109 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110001; // iC= 2097 
// vC = 14'b0000000010010011; // vC=  147 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b0000000010001000; // vC=  136 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010110; // iC= 2198 
// vC = 14'b0000000000010001; // vC=   17 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111011; // iC= 2171 
// vC = 14'b1111111110100110; // vC=  -90 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100010; // iC= 2210 
// vC = 14'b0000000000001011; // vC=   11 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001111; // iC= 1999 
// vC = 14'b0000000001001010; // vC=   74 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110110; // iC= 1974 
// vC = 14'b0000000010101111; // vC=  175 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b0000000011110001; // vC=  241 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b0000000011111001; // vC=  249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000010; // iC= 2114 
// vC = 14'b0000000010110000; // vC=  176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101101; // iC= 2157 
// vC = 14'b1111111111111111; // vC=   -1 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b0000000100001011; // vC=  267 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100010; // iC= 2146 
// vC = 14'b0000000001101101; // vC=  109 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b1111111111110010; // vC=  -14 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100010; // iC= 2018 
// vC = 14'b0000000011011110; // vC=  222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110010; // iC= 2034 
// vC = 14'b0000000001000110; // vC=   70 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000000; // iC= 2048 
// vC = 14'b0000000001101110; // vC=  110 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001001; // iC= 2121 
// vC = 14'b0000000001001111; // vC=   79 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b0000000010001011; // vC=  139 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000100; // iC= 1988 
// vC = 14'b0000000010001010; // vC=  138 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010100; // iC= 2068 
// vC = 14'b0000000100000100; // vC=  260 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b0000000011110111; // vC=  247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001110; // iC= 1934 
// vC = 14'b0000000000110100; // vC=   52 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111010; // iC= 2170 
// vC = 14'b0000000101010101; // vC=  341 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010100; // iC= 2132 
// vC = 14'b0000000101111011; // vC=  379 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001001; // iC= 1865 
// vC = 14'b0000000001010111; // vC=   87 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111001; // iC= 2105 
// vC = 14'b0000000101011101; // vC=  349 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b0000000110100001; // vC=  417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101101; // iC= 2157 
// vC = 14'b0000000011111100; // vC=  252 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101100; // iC= 2156 
// vC = 14'b0000000110100110; // vC=  422 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100001; // iC= 2081 
// vC = 14'b0000000101001100; // vC=  332 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b0000000011000001; // vC=  193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011110; // iC= 2014 
// vC = 14'b0000000110010110; // vC=  406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010011; // iC= 2067 
// vC = 14'b0000000101110111; // vC=  375 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001000; // iC= 1928 
// vC = 14'b0000000011111100; // vC=  252 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b0000000011001100; // vC=  204 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b0000000100100011; // vC=  291 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011011; // iC= 1947 
// vC = 14'b0000000011101111; // vC=  239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b0000000011100110; // vC=  230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001001; // iC= 2057 
// vC = 14'b0000000011100000; // vC=  224 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b0000000110000000; // vC=  384 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b0000000100101100; // vC=  300 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100110; // iC= 1830 
// vC = 14'b0000000110100001; // vC=  417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110101; // iC= 1845 
// vC = 14'b0000000111101100; // vC=  492 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001101; // iC= 1997 
// vC = 14'b0000000101011111; // vC=  351 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000100; // iC= 1988 
// vC = 14'b0000000101110100; // vC=  372 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b0000000101000010; // vC=  322 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010010; // iC= 1874 
// vC = 14'b0000001001001010; // vC=  586 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100111; // iC= 1831 
// vC = 14'b0000000100011001; // vC=  281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101111; // iC= 2095 
// vC = 14'b0000000100111111; // vC=  319 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b0000000101111010; // vC=  378 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011110; // iC= 1822 
// vC = 14'b0000000100111010; // vC=  314 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011010; // iC= 2074 
// vC = 14'b0000001001000011; // vC=  579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b0000001001111101; // vC=  637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111111; // iC= 2111 
// vC = 14'b0000000111011110; // vC=  478 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101010; // iC= 1834 
// vC = 14'b0000001001111011; // vC=  635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b0000000111010010; // vC=  466 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011100; // iC= 1948 
// vC = 14'b0000001000000100; // vC=  516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b0000001001001001; // vC=  585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100100; // iC= 1892 
// vC = 14'b0000001010010100; // vC=  660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b0000001001110011; // vC=  627 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110100; // iC= 2036 
// vC = 14'b0000000111000100; // vC=  452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110010; // iC= 2098 
// vC = 14'b0000001001000000; // vC=  576 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111001; // iC= 1849 
// vC = 14'b0000000110101010; // vC=  426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b0000001011001100; // vC=  716 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b0000000111110011; // vC=  499 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b0000000111111111; // vC=  511 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100101; // iC= 1893 
// vC = 14'b0000000111000010; // vC=  450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110111; // iC= 1783 
// vC = 14'b0000001001100010; // vC=  610 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111011; // iC= 1787 
// vC = 14'b0000001011110000; // vC=  752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b0000000111111100; // vC=  508 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100101; // iC= 1765 
// vC = 14'b0000001000000011; // vC=  515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b0000001011010001; // vC=  721 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010010; // iC= 2066 
// vC = 14'b0000001000111010; // vC=  570 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100110; // iC= 1830 
// vC = 14'b0000001000010010; // vC=  530 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101111; // iC= 1839 
// vC = 14'b0000001010111000; // vC=  696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000100; // iC= 1924 
// vC = 14'b0000001011001010; // vC=  714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b0000001010001111; // vC=  655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b0000001011001101; // vC=  717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110111; // iC= 1847 
// vC = 14'b0000001001111011; // vC=  635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b0000001001101100; // vC=  620 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101001; // iC= 1833 
// vC = 14'b0000001000111110; // vC=  574 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b0000001010010101; // vC=  661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b0000001001000101; // vC=  581 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000000; // iC= 1920 
// vC = 14'b0000001010011111; // vC=  671 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101110; // iC= 2030 
// vC = 14'b0000001001011110; // vC=  606 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b0000001101111001; // vC=  889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100101; // iC= 1701 
// vC = 14'b0000001101010110; // vC=  854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b0000001011110111; // vC=  759 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001100; // iC= 1804 
// vC = 14'b0000001010010010; // vC=  658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101101; // iC= 1709 
// vC = 14'b0000001010100101; // vC=  677 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011011; // iC= 1755 
// vC = 14'b0000001011000110; // vC=  710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101111; // iC= 1903 
// vC = 14'b0000001100110110; // vC=  822 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010001; // iC= 2001 
// vC = 14'b0000001100001110; // vC=  782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100111; // iC= 1703 
// vC = 14'b0000001100000000; // vC=  768 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011000; // iC= 1816 
// vC = 14'b0000001100101001; // vC=  809 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111110; // iC= 1918 
// vC = 14'b0000001110101011; // vC=  939 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101110; // iC= 1774 
// vC = 14'b0000001111001101; // vC=  973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101111; // iC= 1711 
// vC = 14'b0000001100010100; // vC=  788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100111; // iC= 1831 
// vC = 14'b0000001110111110; // vC=  958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110010; // iC= 1842 
// vC = 14'b0000001100011001; // vC=  793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001011; // iC= 1803 
// vC = 14'b0000001111110101; // vC= 1013 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b0000001111001010; // vC=  970 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111010; // iC= 1658 
// vC = 14'b0000001101011101; // vC=  861 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b0000001110000010; // vC=  898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111001; // iC= 1721 
// vC = 14'b0000001101110001; // vC=  881 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111000; // iC= 1784 
// vC = 14'b0000001110011000; // vC=  920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010010; // iC= 1874 
// vC = 14'b0000001110000000; // vC=  896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111001; // iC= 1849 
// vC = 14'b0000001100100101; // vC=  805 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111111; // iC= 1855 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001000; // iC= 1928 
// vC = 14'b0000001110000000; // vC=  896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b0000001110000111; // vC=  903 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001111; // iC= 1743 
// vC = 14'b0000001101101011; // vC=  875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010000; // iC= 1680 
// vC = 14'b0000001100011001; // vC=  793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100010; // iC= 1890 
// vC = 14'b0000001101100101; // vC=  869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111110; // iC= 1662 
// vC = 14'b0000001110001110; // vC=  910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111001; // iC= 1785 
// vC = 14'b0000001100111011; // vC=  827 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101010; // iC= 1770 
// vC = 14'b0000001101010011; // vC=  851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110100; // iC= 1844 
// vC = 14'b0000010001101100; // vC= 1132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100101; // iC= 1893 
// vC = 14'b0000001101110111; // vC=  887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101100; // iC= 1708 
// vC = 14'b0000010000001111; // vC= 1039 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000110; // iC= 1606 
// vC = 14'b0000010001100100; // vC= 1124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001011; // iC= 1611 
// vC = 14'b0000010001000111; // vC= 1095 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101111; // iC= 1839 
// vC = 14'b0000010000011010; // vC= 1050 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100001; // iC= 1697 
// vC = 14'b0000010010001100; // vC= 1164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100100; // iC= 1572 
// vC = 14'b0000001111011000; // vC=  984 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011010; // iC= 1754 
// vC = 14'b0000010001011010; // vC= 1114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111011; // iC= 1595 
// vC = 14'b0000010001010101; // vC= 1109 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111111; // iC= 1855 
// vC = 14'b0000010001011001; // vC= 1113 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001011; // iC= 1803 
// vC = 14'b0000010001101100; // vC= 1132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110011; // iC= 1715 
// vC = 14'b0000001111101101; // vC= 1005 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111110; // iC= 1534 
// vC = 14'b0000010010100000; // vC= 1184 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000100; // iC= 1540 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100111; // iC= 1575 
// vC = 14'b0000010010110001; // vC= 1201 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101001; // iC= 1769 
// vC = 14'b0000010010101101; // vC= 1197 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111010; // iC= 1594 
// vC = 14'b0000010000100101; // vC= 1061 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001011; // iC= 1611 
// vC = 14'b0000010011010110; // vC= 1238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101111; // iC= 1519 
// vC = 14'b0000010001001101; // vC= 1101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010111; // iC= 1751 
// vC = 14'b0000001111011000; // vC=  984 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101111; // iC= 1711 
// vC = 14'b0000001111010011; // vC=  979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100111; // iC= 1767 
// vC = 14'b0000010010001011; // vC= 1163 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111110; // iC= 1534 
// vC = 14'b0000010011001100; // vC= 1228 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111100; // iC= 1724 
// vC = 14'b0000010100011001; // vC= 1305 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000111; // iC= 1671 
// vC = 14'b0000010011000101; // vC= 1221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100000; // iC= 1696 
// vC = 14'b0000010011100001; // vC= 1249 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100111; // iC= 1703 
// vC = 14'b0000010000000100; // vC= 1028 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000000; // iC= 1536 
// vC = 14'b0000010011010111; // vC= 1239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011101; // iC= 1629 
// vC = 14'b0000010011000110; // vC= 1222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001100; // iC= 1548 
// vC = 14'b0000010011000001; // vC= 1217 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101100; // iC= 1708 
// vC = 14'b0000010101010011; // vC= 1363 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110101; // iC= 1461 
// vC = 14'b0000010010011111; // vC= 1183 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011000; // iC= 1752 
// vC = 14'b0000010010010100; // vC= 1172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110101; // iC= 1461 
// vC = 14'b0000010101010011; // vC= 1363 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000100; // iC= 1732 
// vC = 14'b0000010001011011; // vC= 1115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110111; // iC= 1463 
// vC = 14'b0000010100010010; // vC= 1298 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111000; // iC= 1464 
// vC = 14'b0000010010000000; // vC= 1152 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010100; // iC= 1620 
// vC = 14'b0000010001011111; // vC= 1119 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010011; // iC= 1683 
// vC = 14'b0000010110000000; // vC= 1408 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111011; // iC= 1595 
// vC = 14'b0000010100001101; // vC= 1293 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000100; // iC= 1668 
// vC = 14'b0000010101011011; // vC= 1371 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b0000010110010100; // vC= 1428 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111110; // iC= 1534 
// vC = 14'b0000010011110011; // vC= 1267 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101100; // iC= 1580 
// vC = 14'b0000010011010000; // vC= 1232 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100101; // iC= 1637 
// vC = 14'b0000010100000110; // vC= 1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110110; // iC= 1398 
// vC = 14'b0000010100010011; // vC= 1299 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100111; // iC= 1639 
// vC = 14'b0000010110101001; // vC= 1449 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011011; // iC= 1499 
// vC = 14'b0000010100011000; // vC= 1304 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100101; // iC= 1381 
// vC = 14'b0000010110100010; // vC= 1442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000001; // iC= 1409 
// vC = 14'b0000010010110110; // vC= 1206 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110001; // iC= 1649 
// vC = 14'b0000010011001001; // vC= 1225 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110110; // iC= 1590 
// vC = 14'b0000010100011000; // vC= 1304 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011100; // iC= 1564 
// vC = 14'b0000010110111010; // vC= 1466 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110110; // iC= 1526 
// vC = 14'b0000010100101000; // vC= 1320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111111; // iC= 1599 
// vC = 14'b0000010011010110; // vC= 1238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100101; // iC= 1381 
// vC = 14'b0000010111100011; // vC= 1507 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101101; // iC= 1325 
// vC = 14'b0000010100001100; // vC= 1292 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001101; // iC= 1613 
// vC = 14'b0000010100100000; // vC= 1312 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110111; // iC= 1591 
// vC = 14'b0000010100011001; // vC= 1305 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001010; // iC= 1418 
// vC = 14'b0000010100101011; // vC= 1323 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100100; // iC= 1316 
// vC = 14'b0000011000011101; // vC= 1565 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011011; // iC= 1563 
// vC = 14'b0000010101111001; // vC= 1401 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001111; // iC= 1359 
// vC = 14'b0000010011111110; // vC= 1278 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110010; // iC= 1330 
// vC = 14'b0000010110111100; // vC= 1468 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001111; // iC= 1551 
// vC = 14'b0000010110100101; // vC= 1445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101101; // iC= 1581 
// vC = 14'b0000010110011010; // vC= 1434 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011011; // iC= 1371 
// vC = 14'b0000010110001101; // vC= 1421 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101100; // iC= 1516 
// vC = 14'b0000011001000100; // vC= 1604 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001101; // iC= 1485 
// vC = 14'b0000010110001111; // vC= 1423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100001; // iC= 1505 
// vC = 14'b0000010111010100; // vC= 1492 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101110; // iC= 1454 
// vC = 14'b0000011000001100; // vC= 1548 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111001; // iC= 1273 
// vC = 14'b0000011000110100; // vC= 1588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010110; // iC= 1558 
// vC = 14'b0000010111111111; // vC= 1535 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b0000010111101110; // vC= 1518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101100; // iC= 1452 
// vC = 14'b0000011001010010; // vC= 1618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011010; // iC= 1306 
// vC = 14'b0000011001101010; // vC= 1642 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001010; // iC= 1418 
// vC = 14'b0000010111111000; // vC= 1528 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110101; // iC= 1333 
// vC = 14'b0000011000010001; // vC= 1553 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100000; // iC= 1248 
// vC = 14'b0000010110110001; // vC= 1457 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001110; // iC= 1486 
// vC = 14'b0000010110101100; // vC= 1452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001100; // iC= 1356 
// vC = 14'b0000011001110001; // vC= 1649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001110; // iC= 1422 
// vC = 14'b0000011000010000; // vC= 1552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010110; // iC= 1366 
// vC = 14'b0000011001000010; // vC= 1602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110111; // iC= 1207 
// vC = 14'b0000011010010001; // vC= 1681 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100101; // iC= 1445 
// vC = 14'b0000011000110111; // vC= 1591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110000; // iC= 1200 
// vC = 14'b0000011001111111; // vC= 1663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011101; // iC= 1309 
// vC = 14'b0000010111010010; // vC= 1490 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010110; // iC= 1238 
// vC = 14'b0000010110100111; // vC= 1447 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100000; // iC= 1376 
// vC = 14'b0000011001000000; // vC= 1600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001101; // iC= 1421 
// vC = 14'b0000011010001000; // vC= 1672 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001001; // iC= 1161 
// vC = 14'b0000011001000010; // vC= 1602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010010; // iC= 1426 
// vC = 14'b0000011001001010; // vC= 1610 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101010; // iC= 1450 
// vC = 14'b0000010110110001; // vC= 1457 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101100; // iC= 1132 
// vC = 14'b0000011001011001; // vC= 1625 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101110; // iC= 1198 
// vC = 14'b0000011000100010; // vC= 1570 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011001; // iC= 1369 
// vC = 14'b0000011010101101; // vC= 1709 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001000; // iC= 1288 
// vC = 14'b0000011010111000; // vC= 1720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001010; // iC= 1418 
// vC = 14'b0000011010110011; // vC= 1715 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111111; // iC= 1407 
// vC = 14'b0000010110111110; // vC= 1470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010100; // iC= 1236 
// vC = 14'b0000011001011000; // vC= 1624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111000; // iC= 1400 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100001; // iC= 1313 
// vC = 14'b0000011001000001; // vC= 1601 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111100; // iC= 1340 
// vC = 14'b0000011011011101; // vC= 1757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110101; // iC= 1269 
// vC = 14'b0000011000111111; // vC= 1599 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000101; // iC= 1093 
// vC = 14'b0000011000100101; // vC= 1573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001001; // iC= 1289 
// vC = 14'b0000011100001001; // vC= 1801 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001111; // iC= 1359 
// vC = 14'b0000010111010111; // vC= 1495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100011; // iC= 1251 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100000; // iC= 1184 
// vC = 14'b0000011100011010; // vC= 1818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000101; // iC= 1285 
// vC = 14'b0000011000000000; // vC= 1536 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111101; // iC= 1341 
// vC = 14'b0000011011100001; // vC= 1761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100010; // iC= 1058 
// vC = 14'b0000011011011010; // vC= 1754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100011; // iC= 1251 
// vC = 14'b0000011100101100; // vC= 1836 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000010; // iC= 1218 
// vC = 14'b0000011100011011; // vC= 1819 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000101; // iC= 1285 
// vC = 14'b0000011100011111; // vC= 1823 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010001; // iC= 1041 
// vC = 14'b0000011010110011; // vC= 1715 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100110; // iC= 1318 
// vC = 14'b0000011010100010; // vC= 1698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111110; // iC= 1214 
// vC = 14'b0000011000001101; // vC= 1549 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011110; // iC= 1182 
// vC = 14'b0000011000110111; // vC= 1591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000100; // iC= 1284 
// vC = 14'b0000011100111000; // vC= 1848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000100; // iC= 1284 
// vC = 14'b0000011011110000; // vC= 1776 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001000; // iC= 1096 
// vC = 14'b0000011011010110; // vC= 1750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110010; // iC= 1010 
// vC = 14'b0000011010011100; // vC= 1692 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011110; // iC= 1246 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110110; // iC= 1014 
// vC = 14'b0000011100111011; // vC= 1851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110000; // iC= 1264 
// vC = 14'b0000011100111111; // vC= 1855 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100010; // iC=  994 
// vC = 14'b0000011010101000; // vC= 1704 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110110; // iC= 1142 
// vC = 14'b0000011010001111; // vC= 1679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010101; // iC= 1237 
// vC = 14'b0000011100101000; // vC= 1832 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010010; // iC= 1106 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011101; // iC= 1181 
// vC = 14'b0000011010111101; // vC= 1725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010110; // iC= 1046 
// vC = 14'b0000011100111110; // vC= 1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001010; // iC=  906 
// vC = 14'b0000011011011011; // vC= 1755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010010; // iC=  978 
// vC = 14'b0000011010000110; // vC= 1670 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000011; // iC= 1091 
// vC = 14'b0000011101000000; // vC= 1856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010000; // iC=  976 
// vC = 14'b0000011101001000; // vC= 1864 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001000; // iC= 1032 
// vC = 14'b0000011001110111; // vC= 1655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001111; // iC= 1103 
// vC = 14'b0000011011100010; // vC= 1762 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111100; // iC= 1084 
// vC = 14'b0000011010110110; // vC= 1718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001101; // iC= 1165 
// vC = 14'b0000011011100010; // vC= 1762 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100011; // iC=  867 
// vC = 14'b0000011101000111; // vC= 1863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000111; // iC= 1095 
// vC = 14'b0000011011011110; // vC= 1758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001000; // iC= 1096 
// vC = 14'b0000011101011111; // vC= 1887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110100; // iC= 1076 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110101; // iC= 1077 
// vC = 14'b0000011010111110; // vC= 1726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010100; // iC=  916 
// vC = 14'b0000011110000101; // vC= 1925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101101; // iC=  813 
// vC = 14'b0000011100101011; // vC= 1835 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110110; // iC=  822 
// vC = 14'b0000011010101110; // vC= 1710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100011; // iC=  867 
// vC = 14'b0000011100111110; // vC= 1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011010; // iC=  986 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001000; // iC= 1032 
// vC = 14'b0000011111000000; // vC= 1984 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011110; // iC=  798 
// vC = 14'b0000011111001101; // vC= 1997 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101110; // iC=  814 
// vC = 14'b0000011100001000; // vC= 1800 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011111; // iC=  991 
// vC = 14'b0000011100100001; // vC= 1825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111001; // iC=  953 
// vC = 14'b0000011100001110; // vC= 1806 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000000; // iC=  768 
// vC = 14'b0000011100111001; // vC= 1849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011011; // iC=  987 
// vC = 14'b0000011111100000; // vC= 2016 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001101; // iC=  781 
// vC = 14'b0000011011110100; // vC= 1780 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001001; // iC=  969 
// vC = 14'b0000011110000100; // vC= 1924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110100; // iC=  820 
// vC = 14'b0000011011011101; // vC= 1757 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100000; // iC=  992 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100110; // iC=  806 
// vC = 14'b0000011101101100; // vC= 1900 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011001; // iC=  921 
// vC = 14'b0000011111111010; // vC= 2042 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100100; // iC=  996 
// vC = 14'b0000011110111101; // vC= 1981 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011111; // iC=  735 
// vC = 14'b0000011111101000; // vC= 2024 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101100; // iC=  940 
// vC = 14'b0000011111001111; // vC= 1999 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110100; // iC= 1012 
// vC = 14'b0000011100000010; // vC= 1794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010011; // iC=  723 
// vC = 14'b0000011100010001; // vC= 1809 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110111; // iC=  951 
// vC = 14'b0000011111010010; // vC= 2002 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010000; // iC=  720 
// vC = 14'b0000100000010110; // vC= 2070 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101011; // iC=  683 
// vC = 14'b0000100000011100; // vC= 2076 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100000; // iC=  672 
// vC = 14'b0000011100000001; // vC= 1793 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111000; // iC=  952 
// vC = 14'b0000011110111001; // vC= 1977 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111100; // iC=  956 
// vC = 14'b0000011111111110; // vC= 2046 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011111; // iC=  799 
// vC = 14'b0000011100011000; // vC= 1816 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100010; // iC=  866 
// vC = 14'b0000011111100001; // vC= 2017 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000010; // iC=  642 
// vC = 14'b0000011110110111; // vC= 1975 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010111; // iC=  663 
// vC = 14'b0000011100110001; // vC= 1841 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000011; // iC=  643 
// vC = 14'b0000011111110110; // vC= 2038 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010010; // iC=  914 
// vC = 14'b0000100000011010; // vC= 2074 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001000; // iC=  712 
// vC = 14'b0000011100011111; // vC= 1823 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110101; // iC=  693 
// vC = 14'b0000011110100100; // vC= 1956 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000010; // iC=  898 
// vC = 14'b0000011110011100; // vC= 1948 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000000; // iC=  576 
// vC = 14'b0000011111111001; // vC= 2041 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001011; // iC=  587 
// vC = 14'b0000011101011010; // vC= 1882 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111101; // iC=  829 
// vC = 14'b0000100000000001; // vC= 2049 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010111; // iC=  855 
// vC = 14'b0000100001001100; // vC= 2124 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000010; // iC=  834 
// vC = 14'b0000011110000000; // vC= 1920 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111000; // iC=  824 
// vC = 14'b0000011111001111; // vC= 1999 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000101; // iC=  581 
// vC = 14'b0000011100110110; // vC= 1846 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100100; // iC=  548 
// vC = 14'b0000100000110010; // vC= 2098 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001110; // iC=  526 
// vC = 14'b0000011111111100; // vC= 2044 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100010; // iC=  802 
// vC = 14'b0000100000011110; // vC= 2078 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011011; // iC=  795 
// vC = 14'b0000011101101001; // vC= 1897 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111011; // iC=  763 
// vC = 14'b0000100000000100; // vC= 2052 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000110; // iC=  710 
// vC = 14'b0000011110000000; // vC= 1920 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010111; // iC=  535 
// vC = 14'b0000011101010001; // vC= 1873 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111110; // iC=  574 
// vC = 14'b0000011100101001; // vC= 1833 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001001; // iC=  713 
// vC = 14'b0000011101010010; // vC= 1874 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001100; // iC=  716 
// vC = 14'b0000011101100100; // vC= 1892 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110000; // iC=  624 
// vC = 14'b0000100000000100; // vC= 2052 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100100; // iC=  420 
// vC = 14'b0000011111110001; // vC= 2033 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110000; // iC=  624 
// vC = 14'b0000011111010011; // vC= 2003 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010011; // iC=  659 
// vC = 14'b0000011100110001; // vC= 1841 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101111; // iC=  431 
// vC = 14'b0000011111011111; // vC= 2015 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101100; // iC=  492 
// vC = 14'b0000011100110111; // vC= 1847 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100100; // iC=  484 
// vC = 14'b0000100000000100; // vC= 2052 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000111; // iC=  327 
// vC = 14'b0000011110000011; // vC= 1923 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111110; // iC=  318 
// vC = 14'b0000011110110110; // vC= 1974 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111110; // iC=  254 
// vC = 14'b0000011110100111; // vC= 1959 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001111; // iC=  527 
// vC = 14'b0000011111111010; // vC= 2042 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100010; // iC=  226 
// vC = 14'b0000100001001010; // vC= 2122 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011101; // iC=  285 
// vC = 14'b0000100000010101; // vC= 2069 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101010; // iC=  298 
// vC = 14'b0000011110101011; // vC= 1963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010001; // iC=  401 
// vC = 14'b0000100000101011; // vC= 2091 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000111; // iC=  199 
// vC = 14'b0000011101111001; // vC= 1913 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101000; // iC=  232 
// vC = 14'b0000011111001010; // vC= 1994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101001; // iC=  169 
// vC = 14'b0000011111110011; // vC= 2035 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001000; // iC=  136 
// vC = 14'b0000100001010000; // vC= 2128 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011010; // iC=  282 
// vC = 14'b0000011111100001; // vC= 2017 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100001; // iC=  225 
// vC = 14'b0000011110101001; // vC= 1961 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111010; // iC=  250 
// vC = 14'b0000100001010011; // vC= 2131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001110; // iC=  142 
// vC = 14'b0000100000000010; // vC= 2050 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101010; // iC=   42 
// vC = 14'b0000100001111000; // vC= 2168 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000000; // iC=  128 
// vC = 14'b0000100001001000; // vC= 2120 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101101; // iC=   45 
// vC = 14'b0000100000101010; // vC= 2090 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100111; // iC=  231 
// vC = 14'b0000011110000001; // vC= 1921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111011111; // iC=  -33 
// vC = 14'b0000100001111011; // vC= 2171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001000; // iC=  -56 
// vC = 14'b0000100000010000; // vC= 2064 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100010; // iC=  162 
// vC = 14'b0000100010000010; // vC= 2178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010110; // iC=  150 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110100001; // iC=  -95 
// vC = 14'b0000100001111101; // vC= 2173 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100010; // iC=  -30 
// vC = 14'b0000011111010100; // vC= 2004 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101000; // iC=   40 
// vC = 14'b0000011101100010; // vC= 1890 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101011000; // iC= -168 
// vC = 14'b0000011101111011; // vC= 1915 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010011; // iC=  -45 
// vC = 14'b0000011110011111; // vC= 1951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111110011; // iC=  -13 
// vC = 14'b0000100010001101; // vC= 2189 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010000; // iC=  -48 
// vC = 14'b0000011110011001; // vC= 1945 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000000; // iC= -256 
// vC = 14'b0000100001001001; // vC= 2121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101011111; // iC= -161 
// vC = 14'b0000100010000010; // vC= 2178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010101; // iC= -107 
// vC = 14'b0000100000110010; // vC= 2098 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000101; // iC= -251 
// vC = 14'b0000100001100010; // vC= 2146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100100; // iC= -156 
// vC = 14'b0000100001011110; // vC= 2142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100110; // iC= -218 
// vC = 14'b0000100001101100; // vC= 2156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001010; // iC= -182 
// vC = 14'b0000100001111110; // vC= 2174 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010100; // iC= -300 
// vC = 14'b0000100001001011; // vC= 2123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111110; // iC= -386 
// vC = 14'b0000100001011110; // vC= 2142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100001; // iC= -223 
// vC = 14'b0000100000000110; // vC= 2054 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011010; // iC= -230 
// vC = 14'b0000011110111111; // vC= 1983 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001100; // iC= -372 
// vC = 14'b0000100001101100; // vC= 2156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010100; // iC= -364 
// vC = 14'b0000011111111110; // vC= 2046 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000111; // iC= -377 
// vC = 14'b0000100000010100; // vC= 2068 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001101; // iC= -371 
// vC = 14'b0000011101111111; // vC= 1919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000101; // iC= -443 
// vC = 14'b0000011101111100; // vC= 1916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000000; // iC= -640 
// vC = 14'b0000011111100100; // vC= 2020 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000101; // iC= -571 
// vC = 14'b0000011110011101; // vC= 1949 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001111; // iC= -433 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011110; // iC= -482 
// vC = 14'b0000011101101110; // vC= 1902 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001011; // iC= -501 
// vC = 14'b0000011101101111; // vC= 1903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111101; // iC= -579 
// vC = 14'b0000011111110100; // vC= 2036 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001000; // iC= -504 
// vC = 14'b0000100000010011; // vC= 2067 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000100; // iC= -700 
// vC = 14'b0000100000110000; // vC= 2096 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100000; // iC= -736 
// vC = 14'b0000100001001011; // vC= 2123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011000; // iC= -680 
// vC = 14'b0000011111100100; // vC= 2020 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101100; // iC= -724 
// vC = 14'b0000011110000000; // vC= 1920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010100; // iC= -748 
// vC = 14'b0000011100100011; // vC= 1827 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111101; // iC= -835 
// vC = 14'b0000011101010010; // vC= 1874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000100; // iC= -828 
// vC = 14'b0000011111011110; // vC= 2014 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110111; // iC= -969 
// vC = 14'b0000011100110111; // vC= 1847 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011010; // iC= -934 
// vC = 14'b0000011111011101; // vC= 2013 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011100; // iC= -932 
// vC = 14'b0000011111100110; // vC= 2022 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010111; // iC= -809 
// vC = 14'b0000011111011000; // vC= 2008 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010010; // iC=-1006 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110111; // iC=-1033 
// vC = 14'b0000011011111011; // vC= 1787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101110; // iC= -978 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111011; // iC= -965 
// vC = 14'b0000011101010001; // vC= 1873 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101001; // iC=-1047 
// vC = 14'b0000011111010010; // vC= 2002 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011011; // iC=-1061 
// vC = 14'b0000011101100011; // vC= 1891 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110010; // iC=-1166 
// vC = 14'b0000011111110110; // vC= 2038 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101001; // iC= -919 
// vC = 14'b0000011101101111; // vC= 1903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011011; // iC=-1189 
// vC = 14'b0000100000001110; // vC= 2062 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110101; // iC=-1163 
// vC = 14'b0000011111011100; // vC= 2012 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000000; // iC= -960 
// vC = 14'b0000011110001001; // vC= 1929 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101011; // iC=-1045 
// vC = 14'b0000011110101000; // vC= 1960 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000101; // iC=-1147 
// vC = 14'b0000011111101000; // vC= 2024 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001100; // iC=-1204 
// vC = 14'b0000011110001001; // vC= 1929 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010011; // iC=-1325 
// vC = 14'b0000011101110010; // vC= 1906 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011110; // iC=-1058 
// vC = 14'b0000011111001110; // vC= 1998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001101; // iC=-1267 
// vC = 14'b0000011111010100; // vC= 2004 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011001; // iC=-1255 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110001; // iC=-1423 
// vC = 14'b0000011100110010; // vC= 1842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001011; // iC=-1397 
// vC = 14'b0000011010100001; // vC= 1697 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011010; // iC=-1190 
// vC = 14'b0000011111001110; // vC= 1998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101101; // iC=-1427 
// vC = 14'b0000011010100101; // vC= 1701 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010010; // iC=-1262 
// vC = 14'b0000011100110111; // vC= 1847 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000110; // iC=-1466 
// vC = 14'b0000011001111100; // vC= 1660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000010; // iC=-1406 
// vC = 14'b0000011011100011; // vC= 1763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111010; // iC=-1478 
// vC = 14'b0000011110001001; // vC= 1929 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000101; // iC=-1275 
// vC = 14'b0000011001111111; // vC= 1663 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000011; // iC=-1341 
// vC = 14'b0000011011101101; // vC= 1773 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010000; // iC=-1328 
// vC = 14'b0000011010101000; // vC= 1704 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111101; // iC=-1603 
// vC = 14'b0000011011110010; // vC= 1778 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110000; // iC=-1552 
// vC = 14'b0000011100010110; // vC= 1814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011111; // iC=-1505 
// vC = 14'b0000011001000110; // vC= 1606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110010; // iC=-1486 
// vC = 14'b0000011001100011; // vC= 1635 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010010; // iC=-1518 
// vC = 14'b0000011000110110; // vC= 1590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010111; // iC=-1385 
// vC = 14'b0000011100001110; // vC= 1806 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000110; // iC=-1722 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111100; // iC=-1412 
// vC = 14'b0000011100100110; // vC= 1830 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001100; // iC=-1716 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000010; // iC=-1662 
// vC = 14'b0000011100000111; // vC= 1799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000111; // iC=-1593 
// vC = 14'b0000011011101010; // vC= 1770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000011; // iC=-1725 
// vC = 14'b0000011000000111; // vC= 1543 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100001; // iC=-1759 
// vC = 14'b0000011011101010; // vC= 1770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100110; // iC=-1754 
// vC = 14'b0000011010111001; // vC= 1721 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b0000011100110011; // vC= 1843 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111010; // iC=-1542 
// vC = 14'b0000011010010111; // vC= 1687 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b0000011000100101; // vC= 1573 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100011; // iC=-1565 
// vC = 14'b0000011011101001; // vC= 1769 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010001; // iC=-1839 
// vC = 14'b0000010111110111; // vC= 1527 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100110; // iC=-1690 
// vC = 14'b0000010111110011; // vC= 1523 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101100; // iC=-1812 
// vC = 14'b0000011001101100; // vC= 1644 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010000; // iC=-1712 
// vC = 14'b0000011001100111; // vC= 1639 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100100; // iC=-1692 
// vC = 14'b0000010111010010; // vC= 1490 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001101; // iC=-1779 
// vC = 14'b0000011010101100; // vC= 1708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b0000011011001111; // vC= 1743 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b0000011000000111; // vC= 1543 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100111; // iC=-1881 
// vC = 14'b0000010111011100; // vC= 1500 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001100; // iC=-1780 
// vC = 14'b0000011000101010; // vC= 1578 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111110; // iC=-1922 
// vC = 14'b0000011010101000; // vC= 1704 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b0000011010111100; // vC= 1724 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b0000011010001101; // vC= 1677 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b0000011000100010; // vC= 1570 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b0000010111111000; // vC= 1528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001011; // iC=-1973 
// vC = 14'b0000010110000111; // vC= 1415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b0000010110110001; // vC= 1457 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011101; // iC=-1827 
// vC = 14'b0000010110010001; // vC= 1425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b0000011000111101; // vC= 1597 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b0000010111000111; // vC= 1479 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110111; // iC=-1865 
// vC = 14'b0000010111011101; // vC= 1501 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000011000011010; // vC= 1562 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000010110001010; // vC= 1418 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000001; // iC=-1983 
// vC = 14'b0000011000001110; // vC= 1550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b0000010110001110; // vC= 1422 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010101; // iC=-1835 
// vC = 14'b0000010111001111; // vC= 1487 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b0000010110010101; // vC= 1429 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111110; // iC=-2050 
// vC = 14'b0000010101111110; // vC= 1406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100010; // iC=-1822 
// vC = 14'b0000010110100000; // vC= 1440 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b0000010100010110; // vC= 1302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000010101100111; // vC= 1383 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b0000010111110111; // vC= 1527 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000010100100000; // vC= 1312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b0000010011000000; // vC= 1216 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b0000010011101111; // vC= 1263 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b0000010100100100; // vC= 1316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101011; // iC=-2069 
// vC = 14'b0000010110011101; // vC= 1437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b0000010111000011; // vC= 1475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b0000010100111111; // vC= 1343 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b0000010011100101; // vC= 1253 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b0000010110100011; // vC= 1443 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101000; // iC=-1880 
// vC = 14'b0000010011111110; // vC= 1278 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000010011001011; // vC= 1227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101011; // iC=-1877 
// vC = 14'b0000010011100111; // vC= 1255 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100100; // iC=-2140 
// vC = 14'b0000010100100001; // vC= 1313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101001; // iC=-2007 
// vC = 14'b0000010001010111; // vC= 1111 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b0000010001010001; // vC= 1105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110000; // iC=-2192 
// vC = 14'b0000010011101000; // vC= 1256 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101100; // iC=-2004 
// vC = 14'b0000010100010000; // vC= 1296 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100100; // iC=-1884 
// vC = 14'b0000010001100010; // vC= 1122 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111010; // iC=-2182 
// vC = 14'b0000010010000111; // vC= 1159 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111111; // iC=-1921 
// vC = 14'b0000010011010110; // vC= 1238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b0000010000101101; // vC= 1069 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110111; // iC=-2185 
// vC = 14'b0000010010110000; // vC= 1200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000001111111010; // vC= 1018 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000001111111110; // vC= 1022 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010101; // iC=-2027 
// vC = 14'b0000010100000111; // vC= 1287 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111000; // iC=-2184 
// vC = 14'b0000010010110001; // vC= 1201 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001100; // iC=-1908 
// vC = 14'b0000010000010000; // vC= 1040 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011001; // iC=-2215 
// vC = 14'b0000010001111010; // vC= 1146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b0000010000001111; // vC= 1039 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111000; // iC=-2056 
// vC = 14'b0000010010101001; // vC= 1193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100110; // iC=-2202 
// vC = 14'b0000010010000001; // vC= 1153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010000; // iC=-2160 
// vC = 14'b0000010001111101; // vC= 1149 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b0000010011000011; // vC= 1219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100011; // iC=-2141 
// vC = 14'b0000010000101000; // vC= 1064 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110000; // iC=-2064 
// vC = 14'b0000001110111100; // vC=  956 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b0000010010101101; // vC= 1197 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100010; // iC=-2142 
// vC = 14'b0000010000010011; // vC= 1043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100100; // iC=-2204 
// vC = 14'b0000010010011010; // vC= 1178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b0000010001010000; // vC= 1104 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111110; // iC=-2050 
// vC = 14'b0000001110001011; // vC=  907 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100110; // iC=-2202 
// vC = 14'b0000010000111011; // vC= 1083 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010111; // iC=-2025 
// vC = 14'b0000001110000001; // vC=  897 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b0000010000001110; // vC= 1038 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010100; // iC=-2220 
// vC = 14'b0000001110000010; // vC=  898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110010; // iC=-1934 
// vC = 14'b0000010000110111; // vC= 1079 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101111; // iC=-2001 
// vC = 14'b0000001110001001; // vC=  905 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101010; // iC=-2134 
// vC = 14'b0000001100101111; // vC=  815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b0000001111001110; // vC=  974 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010111; // iC=-2153 
// vC = 14'b0000001110111010; // vC=  954 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101110; // iC=-2130 
// vC = 14'b0000001100010011; // vC=  787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001101; // iC=-2163 
// vC = 14'b0000010000101001; // vC= 1065 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b0000010000000011; // vC= 1027 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110011; // iC=-2253 
// vC = 14'b0000001110101011; // vC=  939 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010001; // iC=-2159 
// vC = 14'b0000001101000001; // vC=  833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101111; // iC=-2193 
// vC = 14'b0000001100100101; // vC=  805 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110011; // iC=-2253 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100101; // iC=-2203 
// vC = 14'b0000001101110010; // vC=  882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000001101101111; // vC=  879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101111; // iC=-2257 
// vC = 14'b0000001110010011; // vC=  915 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100011; // iC=-2077 
// vC = 14'b0000001010100100; // vC=  676 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000101; // iC=-2171 
// vC = 14'b0000001010111100; // vC=  700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000011; // iC=-2237 
// vC = 14'b0000001011110111; // vC=  759 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111101; // iC=-2179 
// vC = 14'b0000001100010100; // vC=  788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b0000001011001010; // vC=  714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b0000001110100100; // vC=  932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000001010011010; // vC=  666 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111100; // iC=-2244 
// vC = 14'b0000001010101011; // vC=  683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001101; // iC=-2035 
// vC = 14'b0000001001010010; // vC=  594 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110000; // iC=-2256 
// vC = 14'b0000001011100010; // vC=  738 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110000; // iC=-2128 
// vC = 14'b0000001011000100; // vC=  708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010111; // iC=-2153 
// vC = 14'b0000001100100111; // vC=  807 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100100; // iC=-2140 
// vC = 14'b0000001011011000; // vC=  728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b0000001101000100; // vC=  836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110000; // iC=-2064 
// vC = 14'b0000001010101000; // vC=  680 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000101; // iC=-2171 
// vC = 14'b0000001100001011; // vC=  779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b0000001100110101; // vC=  821 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101111; // iC=-2257 
// vC = 14'b0000001011000111; // vC=  711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110001; // iC=-2191 
// vC = 14'b0000001001001110; // vC=  590 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b0000001011001110; // vC=  718 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b0000001011110001; // vC=  753 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b0000001011010011; // vC=  723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111110; // iC=-2242 
// vC = 14'b0000000111100111; // vC=  487 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011111; // iC=-1953 
// vC = 14'b0000001000111000; // vC=  568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001100; // iC=-2228 
// vC = 14'b0000001011100110; // vC=  742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b0000001011010100; // vC=  724 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011100; // iC=-1956 
// vC = 14'b0000001011000011; // vC=  707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011111; // iC=-2209 
// vC = 14'b0000000111010111; // vC=  471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101000; // iC=-2264 
// vC = 14'b0000000111010110; // vC=  470 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100011101; // iC=-2275 
// vC = 14'b0000000110110100; // vC=  436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b0000000111011011; // vC=  475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b0000000110101010; // vC=  426 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111000; // iC=-2184 
// vC = 14'b0000000111100000; // vC=  480 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b0000000111000100; // vC=  452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b0000001010010000; // vC=  656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101010; // iC=-2134 
// vC = 14'b0000001001110001; // vC=  625 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000001001011010; // vC=  602 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011110; // iC=-2018 
// vC = 14'b0000001001011111; // vC=  607 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010101; // iC=-2155 
// vC = 14'b0000001000010100; // vC=  532 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b0000000101011111; // vC=  351 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100100; // iC=-2140 
// vC = 14'b0000000101001000; // vC=  328 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111110; // iC=-2050 
// vC = 14'b0000000100110110; // vC=  310 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b0000000111010000; // vC=  464 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010101; // iC=-2155 
// vC = 14'b0000000110110011; // vC=  435 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100011; // iC=-1949 
// vC = 14'b0000001000101011; // vC=  555 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000101; // iC=-2043 
// vC = 14'b0000000110011011; // vC=  411 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100100110; // iC=-2266 
// vC = 14'b0000001000001101; // vC=  525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b0000000101001001; // vC=  329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100110; // iC=-2202 
// vC = 14'b0000000100100101; // vC=  293 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b0000000011011001; // vC=  217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b0000000100001110; // vC=  270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100100101; // iC=-2267 
// vC = 14'b0000000011100010; // vC=  226 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b0000000100000110; // vC=  262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000000011001010; // vC=  202 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b0000000111001100; // vC=  460 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010111; // iC=-2217 
// vC = 14'b0000000101101010; // vC=  362 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b0000000101101011; // vC=  363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b0000000101101111; // vC=  367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011110; // iC=-2018 
// vC = 14'b0000000111000110; // vC=  454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001100; // iC=-2164 
// vC = 14'b0000000010010001; // vC=  145 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000000011110010; // vC=  242 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000000110010010; // vC=  402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000100; // iC=-2108 
// vC = 14'b0000000110000111; // vC=  391 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110100; // iC=-2124 
// vC = 14'b0000000001100010; // vC=   98 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b0000000011100100; // vC=  228 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000101; // iC=-2235 
// vC = 14'b0000000100100111; // vC=  295 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111011; // iC=-2117 
// vC = 14'b0000000010111010; // vC=  186 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110101; // iC=-2187 
// vC = 14'b0000000011101111; // vC=  239 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100111; // iC=-2201 
// vC = 14'b0000000001011100; // vC=   92 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000000001001110; // vC=   78 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011100; // iC=-2148 
// vC = 14'b0000000100111101; // vC=  317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000000010010010; // vC=  146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001000; // iC=-2232 
// vC = 14'b0000000001111110; // vC=  126 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000000011000111; // vC=  199 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010101; // iC=-2219 
// vC = 14'b1111111111111111; // vC=   -1 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000011; // iC=-1981 
// vC = 14'b0000000010000010; // vC=  130 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101011; // iC=-2133 
// vC = 14'b0000000010000111; // vC=  135 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b0000000000101100; // vC=   44 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100011; // iC=-1949 
// vC = 14'b0000000100010010; // vC=  274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b0000000001011110; // vC=   94 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100110; // iC=-2202 
// vC = 14'b0000000011010011; // vC=  211 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000000000111110; // vC=   62 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b0000000010011111; // vC=  159 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100101; // iC=-2203 
// vC = 14'b0000000001110011; // vC=  115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000010; // iC=-1918 
// vC = 14'b1111111110111110; // vC=  -66 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101101; // iC=-2195 
// vC = 14'b1111111111111100; // vC=   -4 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000000011001110; // vC=  206 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b0000000010010111; // vC=  151 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b1111111110100111; // vC=  -89 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000000000111111; // vC=   63 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000101; // iC=-2235 
// vC = 14'b1111111110101100; // vC=  -84 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110000; // iC=-2000 
// vC = 14'b0000000000110110; // vC=   54 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101100; // iC=-2196 
// vC = 14'b1111111101011111; // vC= -161 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001111; // iC=-1905 
// vC = 14'b1111111111010001; // vC=  -47 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001011; // iC=-2229 
// vC = 14'b0000000001001111; // vC=   79 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110011; // iC=-2125 
// vC = 14'b1111111110010101; // vC= -107 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010011; // iC=-2221 
// vC = 14'b1111111110011001; // vC= -103 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100001; // iC=-2207 
// vC = 14'b1111111110000001; // vC= -127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b0000000000110100; // vC=   52 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111000; // iC=-2120 
// vC = 14'b1111111101000001; // vC= -191 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110110; // iC=-2122 
// vC = 14'b1111111110100110; // vC=  -90 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b1111111111000001; // vC=  -63 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110000; // iC=-2000 
// vC = 14'b0000000000001010; // vC=   10 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b1111111011110111; // vC= -265 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b1111111111111101; // vC=   -3 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111000; // iC=-2120 
// vC = 14'b1111111111101110; // vC=  -18 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101000; // iC=-2200 
// vC = 14'b1111111101111110; // vC= -130 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011000; // iC=-2088 
// vC = 14'b1111111110111010; // vC=  -70 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110010; // iC=-1934 
// vC = 14'b1111111111100101; // vC=  -27 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b1111111011110000; // vC= -272 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101101; // iC=-2195 
// vC = 14'b1111111100011010; // vC= -230 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101001; // iC=-1879 
// vC = 14'b1111111110110100; // vC=  -76 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111010; // iC=-2118 
// vC = 14'b1111111100100111; // vC= -217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b1111111011101110; // vC= -274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010001; // iC=-2031 
// vC = 14'b1111111100101100; // vC= -212 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b1111111010011101; // vC= -355 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110010; // iC=-2062 
// vC = 14'b1111111011101101; // vC= -275 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b1111111110000111; // vC= -121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000100; // iC=-2044 
// vC = 14'b1111111001101101; // vC= -403 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b1111111101001001; // vC= -183 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b1111111101110111; // vC= -137 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b1111111010001000; // vC= -376 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100010; // iC=-1886 
// vC = 14'b1111111110010001; // vC= -111 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b1111111101001000; // vC= -184 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b1111111010111101; // vC= -323 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000010; // iC=-2046 
// vC = 14'b1111111011010100; // vC= -300 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b1111111100011101; // vC= -227 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000110; // iC=-1978 
// vC = 14'b1111111010100100; // vC= -348 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b1111111001001110; // vC= -434 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000110; // iC=-1978 
// vC = 14'b1111111011001000; // vC= -312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000110; // iC=-1850 
// vC = 14'b1111111010111010; // vC= -326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011111; // iC=-2017 
// vC = 14'b1111111010011011; // vC= -357 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b1111111001101011; // vC= -405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b1111111100011001; // vC= -231 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011111; // iC=-2145 
// vC = 14'b1111111011010011; // vC= -301 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110011; // iC=-1933 
// vC = 14'b1111111010011101; // vC= -355 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b1111111010100010; // vC= -350 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b1111111011011111; // vC= -289 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b1111111010001101; // vC= -371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b1111111011001101; // vC= -307 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b1111111001001011; // vC= -437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011000; // iC=-2088 
// vC = 14'b1111111011011111; // vC= -289 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011100; // iC=-1892 
// vC = 14'b1111111001001011; // vC= -437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b1111111010011110; // vC= -354 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001011; // iC=-1973 
// vC = 14'b1111111000010001; // vC= -495 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b1111111010111000; // vC= -328 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100010; // iC=-1886 
// vC = 14'b1111110110100010; // vC= -606 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100011; // iC=-2077 
// vC = 14'b1111111000011011; // vC= -485 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111100; // iC=-2116 
// vC = 14'b1111111001001110; // vC= -434 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b1111110110100101; // vC= -603 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010110; // iC=-2090 
// vC = 14'b1111111010000011; // vC= -381 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000011; // iC=-1789 
// vC = 14'b1111111000111010; // vC= -454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b1111111000010011; // vC= -493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000010; // iC=-1854 
// vC = 14'b1111110101011000; // vC= -680 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b1111110101001100; // vC= -692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001111; // iC=-1777 
// vC = 14'b1111111000010100; // vC= -492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011001; // iC=-1895 
// vC = 14'b1111110100111010; // vC= -710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b1111110110100111; // vC= -601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011000; // iC=-1832 
// vC = 14'b1111110101100010; // vC= -670 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110010; // iC=-1998 
// vC = 14'b1111110100011101; // vC= -739 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b1111110110011011; // vC= -613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011000; // iC=-2024 
// vC = 14'b1111110101001100; // vC= -692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010110; // iC=-1898 
// vC = 14'b1111110111000010; // vC= -574 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b1111110100100100; // vC= -732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101011; // iC=-2069 
// vC = 14'b1111110011101111; // vC= -785 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010100; // iC=-1900 
// vC = 14'b1111110111001010; // vC= -566 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b1111110011011101; // vC= -803 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b1111110111101010; // vC= -534 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b1111110101101110; // vC= -658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b1111110110011110; // vC= -610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101101; // iC=-1811 
// vC = 14'b1111110100010110; // vC= -746 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b1111110101001010; // vC= -694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b1111110101100101; // vC= -667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110010; // iC=-1742 
// vC = 14'b1111110010110001; // vC= -847 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100101; // iC=-1947 
// vC = 14'b1111110110100100; // vC= -604 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011011; // iC=-1765 
// vC = 14'b1111110110000001; // vC= -639 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b1111110100000110; // vC= -762 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100110; // iC=-1754 
// vC = 14'b1111110010011001; // vC= -871 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100010; // iC=-1758 
// vC = 14'b1111110110100000; // vC= -608 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101000; // iC=-2008 
// vC = 14'b1111110100000101; // vC= -763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b1111110100011100; // vC= -740 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b1111110101001100; // vC= -692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001001; // iC=-1783 
// vC = 14'b1111110100000110; // vC= -762 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100000; // iC=-1824 
// vC = 14'b1111110011110011; // vC= -781 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011101; // iC=-1763 
// vC = 14'b1111110001011101; // vC= -931 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011111; // iC=-1697 
// vC = 14'b1111110100111100; // vC= -708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110000; // iC=-1744 
// vC = 14'b1111110001000110; // vC= -954 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000001; // iC=-1727 
// vC = 14'b1111110001100100; // vC= -924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b1111110100100100; // vC= -732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110011; // iC=-1805 
// vC = 14'b1111110001101001; // vC= -919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b1111110101010000; // vC= -688 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b1111110100111010; // vC= -710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000101; // iC=-1915 
// vC = 14'b1111110000111101; // vC= -963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b1111110100000010; // vC= -766 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010000; // iC=-1648 
// vC = 14'b1111110000000010; // vC=-1022 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111110001011011; // vC= -933 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001110; // iC=-1906 
// vC = 14'b1111101111110101; // vC=-1035 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101001; // iC=-1687 
// vC = 14'b1111110100010001; // vC= -751 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110011; // iC=-1869 
// vC = 14'b1111110001111000; // vC= -904 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110011; // iC=-1869 
// vC = 14'b1111110010101000; // vC= -856 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000111; // iC=-1785 
// vC = 14'b1111110010000111; // vC= -889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010111; // iC=-1769 
// vC = 14'b1111101111111100; // vC=-1028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001000; // iC=-1720 
// vC = 14'b1111101111100111; // vC=-1049 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011011; // iC=-1765 
// vC = 14'b1111101111010010; // vC=-1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b1111101111010010; // vC=-1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011101; // iC=-1827 
// vC = 14'b1111110001010001; // vC= -943 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b1111110010111010; // vC= -838 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100110; // iC=-1754 
// vC = 14'b1111101110101110; // vC=-1106 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111010; // iC=-1734 
// vC = 14'b1111101110110011; // vC=-1101 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010101; // iC=-1707 
// vC = 14'b1111110001010111; // vC= -937 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110001; // iC=-1615 
// vC = 14'b1111101111101111; // vC=-1041 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101111; // iC=-1681 
// vC = 14'b1111110000011110; // vC= -994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010010; // iC=-1646 
// vC = 14'b1111110010100100; // vC= -860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111101; // iC=-1731 
// vC = 14'b1111110010110100; // vC= -844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101111; // iC=-1745 
// vC = 14'b1111101111011000; // vC=-1064 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111000; // iC=-1800 
// vC = 14'b1111110000101101; // vC= -979 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100111; // iC=-1817 
// vC = 14'b1111101101100011; // vC=-1181 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101010; // iC=-1558 
// vC = 14'b1111110001100101; // vC= -923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010000; // iC=-1776 
// vC = 14'b1111110010001111; // vC= -881 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011110; // iC=-1570 
// vC = 14'b1111110000010111; // vC=-1001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010011; // iC=-1837 
// vC = 14'b1111101110101110; // vC=-1106 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110001; // iC=-1679 
// vC = 14'b1111110001100111; // vC= -921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101010; // iC=-1814 
// vC = 14'b1111101101111010; // vC=-1158 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010001; // iC=-1711 
// vC = 14'b1111110001000111; // vC= -953 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000100; // iC=-1532 
// vC = 14'b1111101110101111; // vC=-1105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111101; // iC=-1731 
// vC = 14'b1111101110001010; // vC=-1142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001101; // iC=-1587 
// vC = 14'b1111101100111111; // vC=-1217 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011001; // iC=-1575 
// vC = 14'b1111101100010101; // vC=-1259 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110010; // iC=-1550 
// vC = 14'b1111110000001101; // vC=-1011 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010011; // iC=-1581 
// vC = 14'b1111101100011010; // vC=-1254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011110; // iC=-1634 
// vC = 14'b1111101111101100; // vC=-1044 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101110; // iC=-1746 
// vC = 14'b1111110000011010; // vC= -998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001111; // iC=-1649 
// vC = 14'b1111101111110010; // vC=-1038 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001001; // iC=-1719 
// vC = 14'b1111101101000011; // vC=-1213 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111001; // iC=-1735 
// vC = 14'b1111101011101010; // vC=-1302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011101; // iC=-1699 
// vC = 14'b1111101111101011; // vC=-1045 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110001; // iC=-1615 
// vC = 14'b1111101110001001; // vC=-1143 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100001; // iC=-1503 
// vC = 14'b1111110000001100; // vC=-1012 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000010; // iC=-1534 
// vC = 14'b1111101100111100; // vC=-1220 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111010; // iC=-1606 
// vC = 14'b1111101011010100; // vC=-1324 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110101; // iC=-1483 
// vC = 14'b1111101011010101; // vC=-1323 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101011; // iC=-1685 
// vC = 14'b1111101111010010; // vC=-1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010101; // iC=-1707 
// vC = 14'b1111101101110101; // vC=-1163 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100111; // iC=-1497 
// vC = 14'b1111101100010010; // vC=-1262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001101; // iC=-1715 
// vC = 14'b1111101111010110; // vC=-1066 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101010; // iC=-1558 
// vC = 14'b1111101101000110; // vC=-1210 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111101; // iC=-1667 
// vC = 14'b1111101100101001; // vC=-1239 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000011; // iC=-1661 
// vC = 14'b1111101011011001; // vC=-1319 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110011; // iC=-1485 
// vC = 14'b1111101110111010; // vC=-1094 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110111; // iC=-1545 
// vC = 14'b1111101101100000; // vC=-1184 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111011; // iC=-1477 
// vC = 14'b1111101100101010; // vC=-1238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010101; // iC=-1451 
// vC = 14'b1111101101100100; // vC=-1180 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111000; // iC=-1672 
// vC = 14'b1111101101110000; // vC=-1168 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110111; // iC=-1545 
// vC = 14'b1111101101111110; // vC=-1154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101111; // iC=-1617 
// vC = 14'b1111101101011010; // vC=-1190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011110; // iC=-1506 
// vC = 14'b1111101110011001; // vC=-1127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110101; // iC=-1419 
// vC = 14'b1111101100010000; // vC=-1264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101100; // iC=-1492 
// vC = 14'b1111101010001100; // vC=-1396 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100111; // iC=-1497 
// vC = 14'b1111101101110101; // vC=-1163 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101000; // iC=-1560 
// vC = 14'b1111101011010001; // vC=-1327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111011; // iC=-1413 
// vC = 14'b1111101100011110; // vC=-1250 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100011; // iC=-1501 
// vC = 14'b1111101001101000; // vC=-1432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010000; // iC=-1584 
// vC = 14'b1111101011111011; // vC=-1285 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011100; // iC=-1572 
// vC = 14'b1111101000101001; // vC=-1495 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111010; // iC=-1542 
// vC = 14'b1111101001000000; // vC=-1472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001010; // iC=-1334 
// vC = 14'b1111101010101101; // vC=-1363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000101; // iC=-1403 
// vC = 14'b1111101011101101; // vC=-1299 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101001; // iC=-1431 
// vC = 14'b1111101000010011; // vC=-1517 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101011; // iC=-1365 
// vC = 14'b1111101010010000; // vC=-1392 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000100; // iC=-1340 
// vC = 14'b1111101011111001; // vC=-1287 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010010; // iC=-1518 
// vC = 14'b1111101001010010; // vC=-1454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101110; // iC=-1298 
// vC = 14'b1111101001000010; // vC=-1470 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100101; // iC=-1435 
// vC = 14'b1111101100010011; // vC=-1261 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100101; // iC=-1499 
// vC = 14'b1111101000010110; // vC=-1514 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110000; // iC=-1424 
// vC = 14'b1111101001000011; // vC=-1469 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010011; // iC=-1453 
// vC = 14'b1111101100000110; // vC=-1274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101011; // iC=-1493 
// vC = 14'b1111101100000100; // vC=-1276 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101101; // iC=-1299 
// vC = 14'b1111101011001001; // vC=-1335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010101; // iC=-1515 
// vC = 14'b1111101010010110; // vC=-1386 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101110; // iC=-1554 
// vC = 14'b1111100111111011; // vC=-1541 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110111; // iC=-1289 
// vC = 14'b1111100111101011; // vC=-1557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100110; // iC=-1562 
// vC = 14'b1111100111110001; // vC=-1551 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011100; // iC=-1316 
// vC = 14'b1111101001010010; // vC=-1454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101101; // iC=-1235 
// vC = 14'b1111100111100100; // vC=-1564 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110011; // iC=-1293 
// vC = 14'b1111101000000000; // vC=-1536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011101; // iC=-1507 
// vC = 14'b1111100110110011; // vC=-1613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000000; // iC=-1536 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110001; // iC=-1423 
// vC = 14'b1111101001011011; // vC=-1445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000111; // iC=-1209 
// vC = 14'b1111101010010101; // vC=-1387 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011111; // iC=-1249 
// vC = 14'b1111100111101101; // vC=-1555 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100011; // iC=-1437 
// vC = 14'b1111101001000100; // vC=-1468 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010011; // iC=-1261 
// vC = 14'b1111100110110101; // vC=-1611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111000; // iC=-1224 
// vC = 14'b1111101010110101; // vC=-1355 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100110; // iC=-1242 
// vC = 14'b1111101001110000; // vC=-1424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101111; // iC=-1297 
// vC = 14'b1111101000101111; // vC=-1489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101010; // iC=-1430 
// vC = 14'b1111101010100101; // vC=-1371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011001; // iC=-1191 
// vC = 14'b1111101001010010; // vC=-1454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010001; // iC=-1263 
// vC = 14'b1111101000111100; // vC=-1476 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011001; // iC=-1383 
// vC = 14'b1111101001000110; // vC=-1466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001110; // iC=-1266 
// vC = 14'b1111100110101111; // vC=-1617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010100; // iC=-1388 
// vC = 14'b1111101010010010; // vC=-1390 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110110; // iC=-1226 
// vC = 14'b1111100101011010; // vC=-1702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100001; // iC=-1375 
// vC = 14'b1111100110101011; // vC=-1621 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111000; // iC=-1160 
// vC = 14'b1111101001100000; // vC=-1440 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111011; // iC=-1413 
// vC = 14'b1111100110100000; // vC=-1632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011111; // iC=-1313 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011001; // iC=-1191 
// vC = 14'b1111100111110101; // vC=-1547 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100100; // iC=-1372 
// vC = 14'b1111101001011111; // vC=-1441 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100000; // iC=-1376 
// vC = 14'b1111100101100111; // vC=-1689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111110; // iC=-1090 
// vC = 14'b1111100110100110; // vC=-1626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100011; // iC=-1309 
// vC = 14'b1111100110100001; // vC=-1631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100001; // iC=-1247 
// vC = 14'b1111100100011101; // vC=-1763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111100; // iC=-1220 
// vC = 14'b1111101000010100; // vC=-1516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000100; // iC=-1212 
// vC = 14'b1111100110100001; // vC=-1631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111110; // iC=-1154 
// vC = 14'b1111100101001100; // vC=-1716 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011010; // iC=-1318 
// vC = 14'b1111100101011011; // vC=-1701 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001110; // iC=-1266 
// vC = 14'b1111100110010101; // vC=-1643 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011101; // iC=-1315 
// vC = 14'b1111101000000000; // vC=-1536 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101111; // iC=-1105 
// vC = 14'b1111100100001101; // vC=-1779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010100; // iC=-1324 
// vC = 14'b1111100111100001; // vC=-1567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101000; // iC=-1240 
// vC = 14'b1111100011110111; // vC=-1801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001100; // iC=-1204 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110100; // iC=-1036 
// vC = 14'b1111100011110001; // vC=-1807 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111111; // iC=-1089 
// vC = 14'b1111100111101101; // vC=-1555 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011011; // iC=-1317 
// vC = 14'b1111100110011001; // vC=-1639 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111111; // iC=-1281 
// vC = 14'b1111100110010001; // vC=-1647 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100100; // iC=-1308 
// vC = 14'b1111100110010101; // vC=-1643 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000010; // iC=-1278 
// vC = 14'b1111100110000010; // vC=-1662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111010; // iC=-1030 
// vC = 14'b1111100011010111; // vC=-1833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111001; // iC=-1223 
// vC = 14'b1111100110111111; // vC=-1601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101001; // iC=-1047 
// vC = 14'b1111100100010010; // vC=-1774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101010; // iC=-1110 
// vC = 14'b1111100100110011; // vC=-1741 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001001; // iC=-1207 
// vC = 14'b1111100011100110; // vC=-1818 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001010; // iC=-1078 
// vC = 14'b1111100100100010; // vC=-1758 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111100; // iC=-1156 
// vC = 14'b1111100100100101; // vC=-1755 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b1111100110000000; // vC=-1664 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110110; // iC=-1034 
// vC = 14'b1111100110110000; // vC=-1616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011010; // iC=-1190 
// vC = 14'b1111100110011100; // vC=-1636 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010110; // iC=-1130 
// vC = 14'b1111100011101001; // vC=-1815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100111; // iC=-1177 
// vC = 14'b1111100010010111; // vC=-1897 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111010; // iC=-1158 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101110; // iC=-1042 
// vC = 14'b1111100101011001; // vC=-1703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001000; // iC=-1016 
// vC = 14'b1111100110010000; // vC=-1648 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111110; // iC= -962 
// vC = 14'b1111100010101001; // vC=-1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101011; // iC= -917 
// vC = 14'b1111100110111001; // vC=-1607 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010010; // iC=-1134 
// vC = 14'b1111100100110111; // vC=-1737 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000001; // iC= -959 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011010; // iC=-1062 
// vC = 14'b1111100110101101; // vC=-1619 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001100; // iC=-1076 
// vC = 14'b1111100010111110; // vC=-1858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000001; // iC=-1151 
// vC = 14'b1111100110001110; // vC=-1650 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100011; // iC=-1117 
// vC = 14'b1111100010000000; // vC=-1920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011001; // iC= -871 
// vC = 14'b1111100101011000; // vC=-1704 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000111; // iC=-1145 
// vC = 14'b1111100101011110; // vC=-1698 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010010; // iC=-1006 
// vC = 14'b1111100100011111; // vC=-1761 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011001; // iC= -935 
// vC = 14'b1111100110001001; // vC=-1655 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110100; // iC= -908 
// vC = 14'b1111100010100011; // vC=-1885 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110100; // iC= -844 
// vC = 14'b1111100001110100; // vC=-1932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001110; // iC=-1010 
// vC = 14'b1111100100011110; // vC=-1762 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010001; // iC= -943 
// vC = 14'b1111100010111010; // vC=-1862 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001100; // iC= -948 
// vC = 14'b1111100101001000; // vC=-1720 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100100; // iC= -860 
// vC = 14'b1111100101001001; // vC=-1719 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011111; // iC=-1057 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101111; // iC= -977 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000111; // iC=-1017 
// vC = 14'b1111100001111000; // vC=-1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111110; // iC= -898 
// vC = 14'b1111100001111100; // vC=-1924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110011; // iC=-1037 
// vC = 14'b1111100001010001; // vC=-1967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011000; // iC= -936 
// vC = 14'b1111100001110000; // vC=-1936 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000010; // iC= -894 
// vC = 14'b1111100100000011; // vC=-1789 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111000; // iC= -776 
// vC = 14'b1111100000101010; // vC=-2006 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000101; // iC= -891 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011001; // iC= -935 
// vC = 14'b1111100001101111; // vC=-1937 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000010; // iC= -766 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110010; // iC= -910 
// vC = 14'b1111100001001111; // vC=-1969 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111001; // iC= -711 
// vC = 14'b1111100001001010; // vC=-1974 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101010; // iC= -982 
// vC = 14'b1111100011101010; // vC=-1814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101110; // iC= -722 
// vC = 14'b1111100000101000; // vC=-2008 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101110; // iC= -850 
// vC = 14'b1111100000100101; // vC=-2011 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000011; // iC= -701 
// vC = 14'b1111100011110100; // vC=-1804 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100011; // iC= -669 
// vC = 14'b1111100010100010; // vC=-1886 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100000; // iC= -864 
// vC = 14'b1111100011000101; // vC=-1851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101101; // iC= -787 
// vC = 14'b1111100001101000; // vC=-1944 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110111; // iC= -841 
// vC = 14'b1111100011000111; // vC=-1849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110110; // iC= -778 
// vC = 14'b1111100001110111; // vC=-1929 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111110; // iC= -834 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011100; // iC= -932 
// vC = 14'b1111011111110011; // vC=-2061 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000000; // iC= -704 
// vC = 14'b1111011111101100; // vC=-2068 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101011; // iC= -917 
// vC = 14'b1111011111100101; // vC=-2075 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010001; // iC= -879 
// vC = 14'b1111100000000101; // vC=-2043 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110001; // iC= -719 
// vC = 14'b1111100011101000; // vC=-1816 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000011; // iC= -829 
// vC = 14'b1111100001110000; // vC=-1936 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100001; // iC= -735 
// vC = 14'b1111100001011011; // vC=-1957 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110101; // iC= -651 
// vC = 14'b1111011111011110; // vC=-2082 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101101; // iC= -787 
// vC = 14'b1111100001010101; // vC=-1963 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001100; // iC= -884 
// vC = 14'b1111011111100000; // vC=-2080 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010110; // iC= -874 
// vC = 14'b1111100000110000; // vC=-2000 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011010; // iC= -742 
// vC = 14'b1111011111010100; // vC=-2092 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110110; // iC= -714 
// vC = 14'b1111011111110001; // vC=-2063 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001101; // iC= -691 
// vC = 14'b1111100010001011; // vC=-1909 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000011; // iC= -765 
// vC = 14'b1111100011111110; // vC=-1794 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100011; // iC= -669 
// vC = 14'b1111100010000101; // vC=-1915 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101010; // iC= -662 
// vC = 14'b1111100001000010; // vC=-1982 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010110; // iC= -554 
// vC = 14'b1111100100000000; // vC=-1792 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011111; // iC= -801 
// vC = 14'b1111100000101010; // vC=-2006 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000101; // iC= -635 
// vC = 14'b1111100010001111; // vC=-1905 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001010; // iC= -566 
// vC = 14'b1111100001011101; // vC=-1955 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101010; // iC= -598 
// vC = 14'b1111100001000000; // vC=-1984 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000001001; // iC= -503 
// vC = 14'b1111011111111001; // vC=-2055 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110110; // iC= -650 
// vC = 14'b1111100001010000; // vC=-1968 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010100; // iC= -556 
// vC = 14'b1111011111111010; // vC=-2054 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101011; // iC= -597 
// vC = 14'b1111100001001101; // vC=-1971 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000000; // iC= -640 
// vC = 14'b1111011111101101; // vC=-2067 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011111; // iC= -545 
// vC = 14'b1111100011001011; // vC=-1845 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010111; // iC= -489 
// vC = 14'b1111100001101101; // vC=-1939 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010100; // iC= -684 
// vC = 14'b1111011110110000; // vC=-2128 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110010; // iC= -590 
// vC = 14'b1111100010110001; // vC=-1871 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010110; // iC= -554 
// vC = 14'b1111011111000110; // vC=-2106 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100101; // iC= -411 
// vC = 14'b1111100011000011; // vC=-1853 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000110; // iC= -442 
// vC = 14'b1111100000110100; // vC=-1996 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101101; // iC= -467 
// vC = 14'b1111100000001110; // vC=-2034 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101011; // iC= -533 
// vC = 14'b1111100011001000; // vC=-1848 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001001; // iC= -311 
// vC = 14'b1111100001100010; // vC=-1950 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011110; // iC= -418 
// vC = 14'b1111100010010100; // vC=-1900 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111010; // iC= -390 
// vC = 14'b1111100001010110; // vC=-1962 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100101; // iC= -411 
// vC = 14'b1111011111010011; // vC=-2093 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111111; // iC= -321 
// vC = 14'b1111011111101000; // vC=-2072 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110010; // iC= -398 
// vC = 14'b1111100001001100; // vC=-1972 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000000110; // iC= -506 
// vC = 14'b1111011110101011; // vC=-2133 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001001; // iC= -247 
// vC = 14'b1111100011001111; // vC=-1841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000011; // iC= -381 
// vC = 14'b1111100010101101; // vC=-1875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101111; // iC= -401 
// vC = 14'b1111011111011000; // vC=-2088 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001100; // iC= -372 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001111; // iC= -369 
// vC = 14'b1111100000101001; // vC=-2007 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011100; // iC= -228 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010000; // iC= -304 
// vC = 14'b1111011110111011; // vC=-2117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101001; // iC= -279 
// vC = 14'b1111011111100100; // vC=-2076 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101101; // iC= -211 
// vC = 14'b1111011110100011; // vC=-2141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010000; // iC= -304 
// vC = 14'b1111100000100101; // vC=-2011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011111; // iC= -289 
// vC = 14'b1111100010101111; // vC=-1873 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010100; // iC= -108 
// vC = 14'b1111011110010110; // vC=-2154 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100011; // iC= -221 
// vC = 14'b1111100001110001; // vC=-1935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100110; // iC=   38 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111001; // iC= -135 
// vC = 14'b1111100000101111; // vC=-2001 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011110; // iC=  -98 
// vC = 14'b1111011110001110; // vC=-2162 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010101; // iC=  -43 
// vC = 14'b1111100000001011; // vC=-2037 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000011111; // iC=   31 
// vC = 14'b1111100010000110; // vC=-1914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000100; // iC=  -60 
// vC = 14'b1111100000010010; // vC=-2030 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000011; // iC= -125 
// vC = 14'b1111011111101000; // vC=-2072 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110101; // iC=  117 
// vC = 14'b1111011111101101; // vC=-2067 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101101; // iC=  109 
// vC = 14'b1111100011000000; // vC=-1856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000100; // iC=    4 
// vC = 14'b1111011111100011; // vC=-2077 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001000001; // iC=   65 
// vC = 14'b1111011111010110; // vC=-2090 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011011111; // iC=  223 
// vC = 14'b1111100010101110; // vC=-1874 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000010; // iC=  194 
// vC = 14'b1111011110111110; // vC=-2114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000101010; // iC=   42 
// vC = 14'b1111100000000011; // vC=-2045 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110111; // iC=  119 
// vC = 14'b1111011111101111; // vC=-2065 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010110; // iC=  342 
// vC = 14'b1111011111000100; // vC=-2108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000101; // iC=  325 
// vC = 14'b1111100010100010; // vC=-1886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000111; // iC=  391 
// vC = 14'b1111011111011100; // vC=-2084 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010011; // iC=  275 
// vC = 14'b1111011111011100; // vC=-2084 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100010; // iC=  226 
// vC = 14'b1111100000001000; // vC=-2040 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100110; // iC=  486 
// vC = 14'b1111100000100010; // vC=-2014 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001010; // iC=  394 
// vC = 14'b1111011110110010; // vC=-2126 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100011; // iC=  355 
// vC = 14'b1111011111111111; // vC=-2049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010000; // iC=  336 
// vC = 14'b1111011110101010; // vC=-2134 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011000; // iC=  472 
// vC = 14'b1111100010100100; // vC=-1884 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010011; // iC=  339 
// vC = 14'b1111011111100001; // vC=-2079 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101111; // iC=  367 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110110101; // iC=  437 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000000; // iC=  512 
// vC = 14'b1111100001100011; // vC=-1949 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111111; // iC=  703 
// vC = 14'b1111011110100111; // vC=-2137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001011; // iC=  651 
// vC = 14'b1111100000101101; // vC=-2003 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011010; // iC=  602 
// vC = 14'b1111100001100101; // vC=-1947 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000000; // iC=  640 
// vC = 14'b1111100010011000; // vC=-1896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001011; // iC=  523 
// vC = 14'b1111100001111110; // vC=-1922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100110; // iC=  550 
// vC = 14'b1111100010110001; // vC=-1871 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011011; // iC=  603 
// vC = 14'b1111100010000010; // vC=-1918 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001011; // iC=  779 
// vC = 14'b1111100010101110; // vC=-1874 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111110; // iC=  638 
// vC = 14'b1111100011001011; // vC=-1845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100010; // iC=  738 
// vC = 14'b1111100010011111; // vC=-1889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011001; // iC=  729 
// vC = 14'b1111100001010111; // vC=-1961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110010; // iC=  754 
// vC = 14'b1111100001000000; // vC=-1984 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101011; // iC=  811 
// vC = 14'b1111100010001111; // vC=-1905 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111011; // iC=  763 
// vC = 14'b1111011111010111; // vC=-2089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110101; // iC=  757 
// vC = 14'b1111011111110011; // vC=-2061 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000011; // iC=  963 
// vC = 14'b1111100001011010; // vC=-1958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111101; // iC=  893 
// vC = 14'b1111100011011111; // vC=-1825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010100; // iC=  916 
// vC = 14'b1111100010110011; // vC=-1869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010000; // iC=  912 
// vC = 14'b1111100011000100; // vC=-1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000001; // iC= 1025 
// vC = 14'b1111100010110011; // vC=-1869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111000; // iC= 1080 
// vC = 14'b1111011111110101; // vC=-2059 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000000; // iC=  896 
// vC = 14'b1111100011001001; // vC=-1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110100; // iC=  948 
// vC = 14'b1111100011111100; // vC=-1796 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101011; // iC= 1067 
// vC = 14'b1111100100010011; // vC=-1773 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110110; // iC=  950 
// vC = 14'b1111100001011101; // vC=-1955 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010011; // iC= 1107 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001100; // iC=  972 
// vC = 14'b1111100011001110; // vC=-1842 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101101; // iC= 1133 
// vC = 14'b1111100011110110; // vC=-1802 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010011; // iC= 1043 
// vC = 14'b1111100000010101; // vC=-2027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000111; // iC= 1287 
// vC = 14'b1111100000111101; // vC=-1987 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101100; // iC= 1068 
// vC = 14'b1111100001011000; // vC=-1960 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011111; // iC= 1055 
// vC = 14'b1111100011001000; // vC=-1848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100011; // iC= 1379 
// vC = 14'b1111100011000100; // vC=-1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110010; // iC= 1138 
// vC = 14'b1111100101010001; // vC=-1711 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100000; // iC= 1248 
// vC = 14'b1111100001110101; // vC=-1931 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000011; // iC= 1283 
// vC = 14'b1111100100111010; // vC=-1734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101110; // iC= 1390 
// vC = 14'b1111100110000110; // vC=-1658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101001; // iC= 1385 
// vC = 14'b1111100011111011; // vC=-1797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010101; // iC= 1493 
// vC = 14'b1111100010111110; // vC=-1858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001110; // iC= 1358 
// vC = 14'b1111100110001110; // vC=-1650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111000; // iC= 1272 
// vC = 14'b1111100001101100; // vC=-1940 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010000; // iC= 1424 
// vC = 14'b1111100010000110; // vC=-1914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101100; // iC= 1516 
// vC = 14'b1111100011111100; // vC=-1796 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101001; // iC= 1385 
// vC = 14'b1111100011110001; // vC=-1807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000100; // iC= 1476 
// vC = 14'b1111100100000110; // vC=-1786 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001100; // iC= 1548 
// vC = 14'b1111100010111111; // vC=-1857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100100; // iC= 1444 
// vC = 14'b1111100110101000; // vC=-1624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011001; // iC= 1625 
// vC = 14'b1111100011111101; // vC=-1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110111; // iC= 1527 
// vC = 14'b1111100100100010; // vC=-1758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100000; // iC= 1440 
// vC = 14'b1111100011001001; // vC=-1847 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001100; // iC= 1548 
// vC = 14'b1111100100000010; // vC=-1790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000100; // iC= 1412 
// vC = 14'b1111100011100011; // vC=-1821 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100100; // iC= 1444 
// vC = 14'b1111100100001111; // vC=-1777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010111; // iC= 1559 
// vC = 14'b1111100110100010; // vC=-1630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001000; // iC= 1672 
// vC = 14'b1111100100011100; // vC=-1764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b1111100100010110; // vC=-1770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111000; // iC= 1528 
// vC = 14'b1111100011111011; // vC=-1797 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000001; // iC= 1793 
// vC = 14'b1111100100101001; // vC=-1751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000101; // iC= 1605 
// vC = 14'b1111100110001110; // vC=-1650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111011; // iC= 1531 
// vC = 14'b1111100110100010; // vC=-1630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001111; // iC= 1551 
// vC = 14'b1111100111001001; // vC=-1591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111101; // iC= 1597 
// vC = 14'b1111100111010101; // vC=-1579 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111100; // iC= 1660 
// vC = 14'b1111100100111000; // vC=-1736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010000; // iC= 1616 
// vC = 14'b1111100111011111; // vC=-1569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100000; // iC= 1568 
// vC = 14'b1111100111011111; // vC=-1569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b1111101000111100; // vC=-1476 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001101; // iC= 1677 
// vC = 14'b1111100110001111; // vC=-1649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100000; // iC= 1632 
// vC = 14'b1111100111100010; // vC=-1566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101010; // iC= 1770 
// vC = 14'b1111100101100010; // vC=-1694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000011; // iC= 1731 
// vC = 14'b1111100110101011; // vC=-1621 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100110; // iC= 1830 
// vC = 14'b1111101000110111; // vC=-1481 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000011; // iC= 1859 
// vC = 14'b1111101000110110; // vC=-1482 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b1111101001010110; // vC=-1450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010011; // iC= 1683 
// vC = 14'b1111101001111110; // vC=-1410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111000; // iC= 1976 
// vC = 14'b1111101001001101; // vC=-1459 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100010; // iC= 1762 
// vC = 14'b1111100111110010; // vC=-1550 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010011; // iC= 1747 
// vC = 14'b1111100110100111; // vC=-1625 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111101000111100; // vC=-1476 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b1111101001000001; // vC=-1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110010; // iC= 1778 
// vC = 14'b1111100111001111; // vC=-1585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000101; // iC= 1733 
// vC = 14'b1111100111001100; // vC=-1588 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b1111100111101000; // vC=-1560 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b1111100110100010; // vC=-1630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001000; // iC= 1928 
// vC = 14'b1111101010110000; // vC=-1360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010101; // iC= 1813 
// vC = 14'b1111100111000101; // vC=-1595 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000000; // iC= 1856 
// vC = 14'b1111101001111101; // vC=-1411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b1111101001100100; // vC=-1436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111100; // iC= 1852 
// vC = 14'b1111101010110000; // vC=-1360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100000; // iC= 2016 
// vC = 14'b1111100111100100; // vC=-1564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101010; // iC= 2090 
// vC = 14'b1111101010100110; // vC=-1370 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b1111100111100011; // vC=-1565 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111110; // iC= 1854 
// vC = 14'b1111101010110000; // vC=-1360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110111; // iC= 2039 
// vC = 14'b1111101001110000; // vC=-1424 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000110; // iC= 2118 
// vC = 14'b1111101011001010; // vC=-1334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b1111101100001001; // vC=-1271 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100011; // iC= 1891 
// vC = 14'b1111101010111111; // vC=-1345 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011000; // iC= 2136 
// vC = 14'b1111101100111011; // vC=-1221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011100; // iC= 2140 
// vC = 14'b1111101011001101; // vC=-1331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010001; // iC= 1873 
// vC = 14'b1111101011111111; // vC=-1281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b1111101101010111; // vC=-1193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b1111101001111100; // vC=-1412 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100010; // iC= 2082 
// vC = 14'b1111101101001101; // vC=-1203 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111101011011010; // vC=-1318 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011100; // iC= 2076 
// vC = 14'b1111101101011011; // vC=-1189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110011; // iC= 2099 
// vC = 14'b1111101101110100; // vC=-1164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b1111101110000010; // vC=-1150 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100110; // iC= 2022 
// vC = 14'b1111101010001001; // vC=-1399 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101100; // iC= 1900 
// vC = 14'b1111101110101100; // vC=-1108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100100; // iC= 2020 
// vC = 14'b1111101010010101; // vC=-1387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b1111101111001010; // vC=-1078 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111110; // iC= 1982 
// vC = 14'b1111101100100001; // vC=-1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110001; // iC= 2161 
// vC = 14'b1111101101000101; // vC=-1211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001111; // iC= 2063 
// vC = 14'b1111101010110000; // vC=-1360 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000111; // iC= 2183 
// vC = 14'b1111101101000101; // vC=-1211 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100011; // iC= 2147 
// vC = 14'b1111101100111011; // vC=-1221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111101100001101; // vC=-1267 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000100; // iC= 2180 
// vC = 14'b1111101110110111; // vC=-1097 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001000; // iC= 2120 
// vC = 14'b1111101101110010; // vC=-1166 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b1111101100010101; // vC=-1259 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000101; // iC= 2181 
// vC = 14'b1111101110110110; // vC=-1098 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111000; // iC= 2168 
// vC = 14'b1111101101101000; // vC=-1176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011011; // iC= 2139 
// vC = 14'b1111110000100010; // vC= -990 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001010; // iC= 2058 
// vC = 14'b1111101110100101; // vC=-1115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110110; // iC= 2102 
// vC = 14'b1111101110000001; // vC=-1151 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101110; // iC= 1966 
// vC = 14'b1111101110000000; // vC=-1152 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b1111101111110001; // vC=-1039 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100000; // iC= 2016 
// vC = 14'b1111101111111101; // vC=-1027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010010; // iC= 2002 
// vC = 14'b1111101100111010; // vC=-1222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011011; // iC= 2203 
// vC = 14'b1111101110101000; // vC=-1112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001111; // iC= 2191 
// vC = 14'b1111101101111111; // vC=-1153 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111100; // iC= 2172 
// vC = 14'b1111101110001010; // vC=-1142 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111101; // iC= 2045 
// vC = 14'b1111110000101011; // vC= -981 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b1111101110101001; // vC=-1111 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000011; // iC= 2179 
// vC = 14'b1111101101111010; // vC=-1158 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000001; // iC= 2177 
// vC = 14'b1111101111001011; // vC=-1077 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b1111101110101111; // vC=-1105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b1111110010110010; // vC= -846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111110010100111; // vC= -857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000000; // iC= 2176 
// vC = 14'b1111110000010101; // vC=-1003 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110010; // iC= 2162 
// vC = 14'b1111101110011011; // vC=-1125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110001; // iC= 2225 
// vC = 14'b1111110001101011; // vC= -917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111110010010111; // vC= -873 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b1111101111010110; // vC=-1066 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110111; // iC= 2039 
// vC = 14'b1111110001001111; // vC= -945 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010011; // iC= 2131 
// vC = 14'b1111101111011101; // vC=-1059 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b1111110011010000; // vC= -816 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110100; // iC= 2100 
// vC = 14'b1111110010111000; // vC= -840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101100; // iC= 2156 
// vC = 14'b1111110010000101; // vC= -891 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111110100100100; // vC= -732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100000; // iC= 2144 
// vC = 14'b1111110100000110; // vC= -762 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b1111110100100010; // vC= -734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b1111110011110101; // vC= -779 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111110011101010; // vC= -790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b1111110001111001; // vC= -903 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101001; // iC= 2217 
// vC = 14'b1111110000110011; // vC= -973 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b1111110001011011; // vC= -933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b1111110001010110; // vC= -938 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001011; // iC= 2251 
// vC = 14'b1111110101101101; // vC= -659 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b1111110101011010; // vC= -678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011110; // iC= 2142 
// vC = 14'b1111110001110101; // vC= -907 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100001; // iC= 2081 
// vC = 14'b1111110101011010; // vC= -678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001101; // iC= 2253 
// vC = 14'b1111110101100010; // vC= -670 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010101; // iC= 2069 
// vC = 14'b1111110100000100; // vC= -764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001001; // iC= 2249 
// vC = 14'b1111110110101000; // vC= -600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000101; // iC= 1989 
// vC = 14'b1111110010110111; // vC= -841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101001; // iC= 2153 
// vC = 14'b1111110011000010; // vC= -830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111110100000111; // vC= -761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111011; // iC= 2235 
// vC = 14'b1111110010101101; // vC= -851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000001; // iC= 2241 
// vC = 14'b1111110101101011; // vC= -661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010010; // iC= 2258 
// vC = 14'b1111110100001101; // vC= -755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100100; // iC= 2212 
// vC = 14'b1111110111110110; // vC= -522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111110; // iC= 2174 
// vC = 14'b1111110100001010; // vC= -758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111110101101111; // vC= -657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110000; // iC= 2160 
// vC = 14'b1111110110000111; // vC= -633 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110000; // iC= 2160 
// vC = 14'b1111110100111101; // vC= -707 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101101; // iC= 2157 
// vC = 14'b1111110101101101; // vC= -659 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011011; // iC= 2075 
// vC = 14'b1111111000100101; // vC= -475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000101; // iC= 2053 
// vC = 14'b1111110101101100; // vC= -660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b1111110011111101; // vC= -771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b1111110111110101; // vC= -523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b1111110101000101; // vC= -699 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b1111110111011000; // vC= -552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000100; // iC= 2180 
// vC = 14'b1111110111011010; // vC= -550 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111111; // iC= 2175 
// vC = 14'b1111110110101100; // vC= -596 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011111; // iC= 2079 
// vC = 14'b1111110101110000; // vC= -656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001100; // iC= 2252 
// vC = 14'b1111111000001010; // vC= -502 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b1111111000111110; // vC= -450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111011; // iC= 2235 
// vC = 14'b1111110111100110; // vC= -538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100111; // iC= 2087 
// vC = 14'b1111110110000000; // vC= -640 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010000; // iC= 2064 
// vC = 14'b1111111000001001; // vC= -503 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011011; // iC= 2075 
// vC = 14'b1111111000111101; // vC= -451 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111111010110010; // vC= -334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110001; // iC= 2097 
// vC = 14'b1111111000010101; // vC= -491 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b1111110111101001; // vC= -535 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111111001111110; // vC= -386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111000; // iC= 1976 
// vC = 14'b1111111001000010; // vC= -446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010110; // iC= 2134 
// vC = 14'b1111110111111100; // vC= -516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001101; // iC= 1997 
// vC = 14'b1111111000011110; // vC= -482 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001111; // iC= 2191 
// vC = 14'b1111110111111100; // vC= -516 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001000; // iC= 2184 
// vC = 14'b1111111011101011; // vC= -277 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100101; // iC= 2213 
// vC = 14'b1111111010110010; // vC= -334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100001; // iC= 2145 
// vC = 14'b1111111010000000; // vC= -384 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000100; // iC= 2180 
// vC = 14'b1111111100010010; // vC= -238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010101; // iC= 2197 
// vC = 14'b1111111000101100; // vC= -468 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111001; // iC= 2233 
// vC = 14'b1111111000010110; // vC= -490 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111111001001100; // vC= -436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011000; // iC= 2136 
// vC = 14'b1111111010110001; // vC= -335 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010110; // iC= 2070 
// vC = 14'b1111111100001001; // vC= -247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001000; // iC= 2248 
// vC = 14'b1111111010000000; // vC= -384 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b1111111001010110; // vC= -426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100100; // iC= 2212 
// vC = 14'b1111111001001111; // vC= -433 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b1111111101011011; // vC= -165 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001101; // iC= 1997 
// vC = 14'b1111111001000011; // vC= -445 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110100; // iC= 2036 
// vC = 14'b1111111010111001; // vC= -327 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000101; // iC= 2053 
// vC = 14'b1111111011100010; // vC= -286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b1111111010110000; // vC= -336 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100011; // iC= 2147 
// vC = 14'b1111111100110100; // vC= -204 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b1111111011110000; // vC= -272 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010001; // iC= 2257 
// vC = 14'b1111111010101001; // vC= -343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010001; // iC= 2257 
// vC = 14'b1111111010100111; // vC= -345 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000001; // iC= 2241 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011111; // iC= 2143 
// vC = 14'b1111111100000010; // vC= -254 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101100; // iC= 2092 
// vC = 14'b1111111100100011; // vC= -221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111111011000101; // vC= -315 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110010; // iC= 2162 
// vC = 14'b1111111111100101; // vC=  -27 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000000; // iC= 2176 
// vC = 14'b1111111100111111; // vC= -193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101000; // iC= 2152 
// vC = 14'b1111111111101110; // vC=  -18 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b1111111101111100; // vC= -132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010101; // iC= 2133 
// vC = 14'b1111111101001111; // vC= -177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000001; // iC= 2049 
// vC = 14'b1111111101010100; // vC= -172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110101; // iC= 2165 
// vC = 14'b1111111101000111; // vC= -185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100011; // iC= 1955 
// vC = 14'b1111111101011101; // vC= -163 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011100; // iC= 2076 
// vC = 14'b1111111101110101; // vC= -139 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011000000; // iC= 2240 
// vC = 14'b1111111101011100; // vC= -164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001010; // iC= 1994 
// vC = 14'b0000000000010110; // vC=   22 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b0000000000001001; // vC=    9 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111000; // iC= 2104 
// vC = 14'b0000000001001110; // vC=   78 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000010; // iC= 1922 
// vC = 14'b0000000000010010; // vC=   18 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b1111111101000010; // vC= -190 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b1111111111001000; // vC=  -56 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111111110000110; // vC= -122 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000000; // iC= 2048 
// vC = 14'b1111111111111111; // vC=   -1 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101100; // iC= 2220 
// vC = 14'b0000000001111110; // vC=  126 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111111110011100; // vC= -100 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000010; // iC= 1986 
// vC = 14'b1111111110011011; // vC= -101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b1111111110101100; // vC=  -84 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111111111001110; // vC=  -50 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b0000000000001111; // vC=   15 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110000; // iC= 2160 
// vC = 14'b1111111101111111; // vC= -129 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100111; // iC= 2023 
// vC = 14'b0000000010111010; // vC=  186 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000000; // iC= 2048 
// vC = 14'b0000000010100011; // vC=  163 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b1111111111010011; // vC=  -45 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111001; // iC= 2105 
// vC = 14'b0000000000101111; // vC=   47 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011100; // iC= 2140 
// vC = 14'b0000000000101110; // vC=   46 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b0000000010100100; // vC=  164 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111110; // iC= 2046 
// vC = 14'b0000000010101111; // vC=  175 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111100; // iC= 1980 
// vC = 14'b0000000010000000; // vC=  128 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001110; // iC= 2126 
// vC = 14'b0000000010110101; // vC=  181 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b0000000010110011; // vC=  179 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b0000000000011000; // vC=   24 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111110; // iC= 2174 
// vC = 14'b0000000100000110; // vC=  262 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101110; // iC= 1966 
// vC = 14'b1111111111111000; // vC=   -8 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010001; // iC= 2129 
// vC = 14'b0000000001101111; // vC=  111 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000101; // iC= 1925 
// vC = 14'b0000000100100111; // vC=  295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b0000000011000111; // vC=  199 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b0000000010111110; // vC=  190 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000010; // iC= 2178 
// vC = 14'b0000000100101111; // vC=  303 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b0000000010001001; // vC=  137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b0000000101001101; // vC=  333 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b0000000010101101; // vC=  173 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001001; // iC= 1993 
// vC = 14'b0000000101110010; // vC=  370 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b0000000001100000; // vC=   96 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b0000000001110011; // vC=  115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111000; // iC= 2104 
// vC = 14'b0000000001100101; // vC=  101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010010; // iC= 1874 
// vC = 14'b0000000110010101; // vC=  405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b0000000010010110; // vC=  150 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b0000000100110100; // vC=  308 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011010; // iC= 2138 
// vC = 14'b0000000010000100; // vC=  132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b0000000110010010; // vC=  402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001111; // iC= 2063 
// vC = 14'b0000000100001010; // vC=  266 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110011; // iC= 1971 
// vC = 14'b0000000011010111; // vC=  215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101110; // iC= 2158 
// vC = 14'b0000000100111001; // vC=  313 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011010; // iC= 2138 
// vC = 14'b0000000101011010; // vC=  346 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111100; // iC= 1980 
// vC = 14'b0000000111001111; // vC=  463 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b0000000101010111; // vC=  343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b0000000110000000; // vC=  384 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000000100010000; // vC=  272 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100011; // iC= 1955 
// vC = 14'b0000000111011101; // vC=  477 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b0000000011110111; // vC=  247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100001; // iC= 1953 
// vC = 14'b0000000111100111; // vC=  487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b0000000100001101; // vC=  269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111110; // iC= 1854 
// vC = 14'b0000000110011011; // vC=  411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111111; // iC= 1919 
// vC = 14'b0000000100011000; // vC=  280 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b0000001000010100; // vC=  532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b0000000101100001; // vC=  353 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b0000000110001001; // vC=  393 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000110; // iC= 1862 
// vC = 14'b0000000110010101; // vC=  405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010001; // iC= 1873 
// vC = 14'b0000000111111110; // vC=  510 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b0000001000010000; // vC=  528 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001101; // iC= 2125 
// vC = 14'b0000000101001110; // vC=  334 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011110; // iC= 2078 
// vC = 14'b0000000110111011; // vC=  443 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110001; // iC= 1905 
// vC = 14'b0000001001000110; // vC=  582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010110; // iC= 1814 
// vC = 14'b0000001000100110; // vC=  550 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110001; // iC= 2097 
// vC = 14'b0000001000000111; // vC=  519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101101; // iC= 2093 
// vC = 14'b0000001001001010; // vC=  586 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000010; // iC= 2050 
// vC = 14'b0000001010001010; // vC=  650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001100; // iC= 1804 
// vC = 14'b0000000111000111; // vC=  455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b0000000111000111; // vC=  455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b0000000110010000; // vC=  400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011111; // iC= 1887 
// vC = 14'b0000000111110101; // vC=  501 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100010; // iC= 2082 
// vC = 14'b0000000111100100; // vC=  484 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111100; // iC= 1980 
// vC = 14'b0000001001000110; // vC=  582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011100; // iC= 2012 
// vC = 14'b0000001011001001; // vC=  713 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010101; // iC= 1813 
// vC = 14'b0000001010010010; // vC=  658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010010; // iC= 2002 
// vC = 14'b0000001010110100; // vC=  692 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b0000001001011100; // vC=  604 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100111; // iC= 1895 
// vC = 14'b0000001000011000; // vC=  536 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101110; // iC= 1902 
// vC = 14'b0000000111010011; // vC=  467 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011001; // iC= 2009 
// vC = 14'b0000001001000111; // vC=  583 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111011; // iC= 1915 
// vC = 14'b0000001000101100; // vC=  556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b0000001010001010; // vC=  650 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111100; // iC= 1916 
// vC = 14'b0000001011011000; // vC=  728 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100100; // iC= 1828 
// vC = 14'b0000001001010011; // vC=  595 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b0000001000101101; // vC=  557 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b0000001010111001; // vC=  697 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111110; // iC= 1918 
// vC = 14'b0000001001011110; // vC=  606 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010101; // iC= 2005 
// vC = 14'b0000001011101010; // vC=  746 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b0000001101011110; // vC=  862 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b0000001001000110; // vC=  582 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110100; // iC= 1716 
// vC = 14'b0000001010100101; // vC=  677 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000101; // iC= 1733 
// vC = 14'b0000001001001101; // vC=  589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b0000001101111100; // vC=  892 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110010; // iC= 1842 
// vC = 14'b0000001010100101; // vC=  677 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011110; // iC= 2014 
// vC = 14'b0000001001001101; // vC=  589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b0000001010011000; // vC=  664 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100010; // iC= 2018 
// vC = 14'b0000001101001101; // vC=  845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000001; // iC= 1729 
// vC = 14'b0000001010001101; // vC=  653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011010; // iC= 1882 
// vC = 14'b0000001101000010; // vC=  834 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100001; // iC= 1761 
// vC = 14'b0000001011011111; // vC=  735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001000; // iC= 1928 
// vC = 14'b0000001010001100; // vC=  652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100011; // iC= 1955 
// vC = 14'b0000001011010110; // vC=  726 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101000; // iC= 1832 
// vC = 14'b0000001100000001; // vC=  769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010111; // iC= 1815 
// vC = 14'b0000001100000111; // vC=  775 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b0000001110111000; // vC=  952 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000101; // iC= 1797 
// vC = 14'b0000001110010010; // vC=  914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010101; // iC= 1749 
// vC = 14'b0000001011011100; // vC=  732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001110; // iC= 1870 
// vC = 14'b0000001100101010; // vC=  810 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010100; // iC= 1684 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b0000001101011111; // vC=  863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101010; // iC= 1706 
// vC = 14'b0000001100110010; // vC=  818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000010; // iC= 1794 
// vC = 14'b0000001011100001; // vC=  737 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100101; // iC= 1829 
// vC = 14'b0000001110111100; // vC=  956 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b0000001110111011; // vC=  955 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001110; // iC= 1742 
// vC = 14'b0000001110000000; // vC=  896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111111; // iC= 1727 
// vC = 14'b0000001111101010; // vC= 1002 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011100; // iC= 1628 
// vC = 14'b0000001100101111; // vC=  815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010110; // iC= 1622 
// vC = 14'b0000010000101001; // vC= 1065 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000101; // iC= 1797 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001101; // iC= 1869 
// vC = 14'b0000010000101110; // vC= 1070 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011100; // iC= 1756 
// vC = 14'b0000001110111011; // vC=  955 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010011; // iC= 1747 
// vC = 14'b0000001110011110; // vC=  926 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000100; // iC= 1796 
// vC = 14'b0000001100101100; // vC=  812 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101100; // iC= 1900 
// vC = 14'b0000001110011010; // vC=  922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110011; // iC= 1651 
// vC = 14'b0000010001100111; // vC= 1127 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011000; // iC= 1688 
// vC = 14'b0000010000110001; // vC= 1073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b0000001101101011; // vC=  875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101110; // iC= 1582 
// vC = 14'b0000001110010100; // vC=  916 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000100; // iC= 1604 
// vC = 14'b0000010001111111; // vC= 1151 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111000; // iC= 1592 
// vC = 14'b0000001101101110; // vC=  878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000100; // iC= 1604 
// vC = 14'b0000010001000011; // vC= 1091 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101010; // iC= 1706 
// vC = 14'b0000010010100110; // vC= 1190 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100110; // iC= 1702 
// vC = 14'b0000001111110011; // vC= 1011 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000011; // iC= 1859 
// vC = 14'b0000010000101000; // vC= 1064 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011110; // iC= 1694 
// vC = 14'b0000010000110001; // vC= 1073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000101; // iC= 1733 
// vC = 14'b0000001110100011; // vC=  931 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111101; // iC= 1789 
// vC = 14'b0000010011000101; // vC= 1221 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111010; // iC= 1658 
// vC = 14'b0000010000011011; // vC= 1051 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010101; // iC= 1685 
// vC = 14'b0000010000000110; // vC= 1030 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111001; // iC= 1785 
// vC = 14'b0000010000100010; // vC= 1058 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001100; // iC= 1740 
// vC = 14'b0000010001010111; // vC= 1111 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110100; // iC= 1588 
// vC = 14'b0000010000000011; // vC= 1027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110101; // iC= 1589 
// vC = 14'b0000001111010000; // vC=  976 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001010; // iC= 1738 
// vC = 14'b0000010000100110; // vC= 1062 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110000; // iC= 1776 
// vC = 14'b0000010010000101; // vC= 1157 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000010; // iC= 1602 
// vC = 14'b0000010010010011; // vC= 1171 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111110; // iC= 1726 
// vC = 14'b0000001111110001; // vC= 1009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001010; // iC= 1610 
// vC = 14'b0000010011111110; // vC= 1278 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101011; // iC= 1771 
// vC = 14'b0000010000011010; // vC= 1050 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110101; // iC= 1589 
// vC = 14'b0000010000101101; // vC= 1069 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110011; // iC= 1587 
// vC = 14'b0000010011010001; // vC= 1233 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011001; // iC= 1753 
// vC = 14'b0000010010010100; // vC= 1172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010001; // iC= 1489 
// vC = 14'b0000010000011000; // vC= 1048 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110100; // iC= 1652 
// vC = 14'b0000010000101000; // vC= 1064 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100001; // iC= 1569 
// vC = 14'b0000010001000100; // vC= 1092 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110010; // iC= 1714 
// vC = 14'b0000010001011110; // vC= 1118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000011; // iC= 1603 
// vC = 14'b0000010000110110; // vC= 1078 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001101; // iC= 1549 
// vC = 14'b0000010011001100; // vC= 1228 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100000; // iC= 1632 
// vC = 14'b0000010010101011; // vC= 1195 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100111; // iC= 1447 
// vC = 14'b0000010001101010; // vC= 1130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011100; // iC= 1756 
// vC = 14'b0000010100011111; // vC= 1311 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001010; // iC= 1482 
// vC = 14'b0000010001110101; // vC= 1141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110010; // iC= 1650 
// vC = 14'b0000010011001101; // vC= 1229 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010010; // iC= 1426 
// vC = 14'b0000010011010110; // vC= 1238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101000; // iC= 1576 
// vC = 14'b0000010001100011; // vC= 1123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001111; // iC= 1551 
// vC = 14'b0000010101110010; // vC= 1394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100111; // iC= 1447 
// vC = 14'b0000010011010111; // vC= 1239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100100; // iC= 1444 
// vC = 14'b0000010110100011; // vC= 1443 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011001; // iC= 1561 
// vC = 14'b0000010010011110; // vC= 1182 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001101; // iC= 1549 
// vC = 14'b0000010100111111; // vC= 1343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000101; // iC= 1413 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101001; // iC= 1449 
// vC = 14'b0000010100010101; // vC= 1301 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010010; // iC= 1490 
// vC = 14'b0000010111000101; // vC= 1477 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011111; // iC= 1567 
// vC = 14'b0000010101011110; // vC= 1374 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001010; // iC= 1418 
// vC = 14'b0000010110011101; // vC= 1437 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010010; // iC= 1362 
// vC = 14'b0000010110101010; // vC= 1450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101011; // iC= 1579 
// vC = 14'b0000010011111100; // vC= 1276 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001001; // iC= 1417 
// vC = 14'b0000010101001000; // vC= 1352 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110111; // iC= 1463 
// vC = 14'b0000010011100110; // vC= 1254 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000001; // iC= 1345 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111111; // iC= 1471 
// vC = 14'b0000010010111001; // vC= 1209 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000011; // iC= 1603 
// vC = 14'b0000010011000001; // vC= 1217 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101110; // iC= 1390 
// vC = 14'b0000010111101011; // vC= 1515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011010; // iC= 1434 
// vC = 14'b0000010100001100; // vC= 1292 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b0000010100111110; // vC= 1342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100110; // iC= 1574 
// vC = 14'b0000010101111010; // vC= 1402 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011110; // iC= 1374 
// vC = 14'b0000010111011101; // vC= 1501 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111111; // iC= 1535 
// vC = 14'b0000010100101001; // vC= 1321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b0000010110010110; // vC= 1430 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101011; // iC= 1515 
// vC = 14'b0000010101001011; // vC= 1355 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110101; // iC= 1333 
// vC = 14'b0000010110110110; // vC= 1462 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000101; // iC= 1605 
// vC = 14'b0000011000000100; // vC= 1540 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101110; // iC= 1390 
// vC = 14'b0000010100110011; // vC= 1331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100110; // iC= 1446 
// vC = 14'b0000010111001000; // vC= 1480 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101100; // iC= 1516 
// vC = 14'b0000011001000011; // vC= 1603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110011; // iC= 1459 
// vC = 14'b0000010100110001; // vC= 1329 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111010; // iC= 1274 
// vC = 14'b0000010111101011; // vC= 1515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111011; // iC= 1531 
// vC = 14'b0000010110111111; // vC= 1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111110; // iC= 1470 
// vC = 14'b0000010110000011; // vC= 1411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101101; // iC= 1517 
// vC = 14'b0000010111010100; // vC= 1492 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100011; // iC= 1251 
// vC = 14'b0000010101100011; // vC= 1379 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001111; // iC= 1423 
// vC = 14'b0000010101001101; // vC= 1357 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011011; // iC= 1243 
// vC = 14'b0000010101111000; // vC= 1400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111110; // iC= 1534 
// vC = 14'b0000010111101111; // vC= 1519 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101011100; // iC= 1372 
// vC = 14'b0000011000010100; // vC= 1556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100011; // iC= 1443 
// vC = 14'b0000010111101001; // vC= 1513 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100011; // iC= 1251 
// vC = 14'b0000011001010100; // vC= 1620 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110001; // iC= 1393 
// vC = 14'b0000011001010011; // vC= 1619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101011; // iC= 1451 
// vC = 14'b0000011000010111; // vC= 1559 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001010; // iC= 1226 
// vC = 14'b0000011000101000; // vC= 1576 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011000; // iC= 1496 
// vC = 14'b0000011001101101; // vC= 1645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011010; // iC= 1434 
// vC = 14'b0000011001111101; // vC= 1661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010001; // iC= 1169 
// vC = 14'b0000010110110000; // vC= 1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000010; // iC= 1474 
// vC = 14'b0000010101110111; // vC= 1399 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101101; // iC= 1325 
// vC = 14'b0000011010000110; // vC= 1670 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111111; // iC= 1215 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110011; // iC= 1395 
// vC = 14'b0000011001001001; // vC= 1609 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101111; // iC= 1199 
// vC = 14'b0000010110001011; // vC= 1419 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110011; // iC= 1331 
// vC = 14'b0000010111111101; // vC= 1533 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111111; // iC= 1215 
// vC = 14'b0000010111011011; // vC= 1499 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111111; // iC= 1407 
// vC = 14'b0000011001101111; // vC= 1647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101110; // iC= 1326 
// vC = 14'b0000011000010010; // vC= 1554 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100110; // iC= 1382 
// vC = 14'b0000010111100110; // vC= 1510 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101001; // iC= 1129 
// vC = 14'b0000011011010110; // vC= 1750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000010; // iC= 1410 
// vC = 14'b0000011010001010; // vC= 1674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111100; // iC= 1404 
// vC = 14'b0000011001100010; // vC= 1634 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111101; // iC= 1405 
// vC = 14'b0000010111001110; // vC= 1486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100010; // iC= 1314 
// vC = 14'b0000011000000001; // vC= 1537 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100110; // iC= 1126 
// vC = 14'b0000010111100010; // vC= 1506 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000110; // iC= 1094 
// vC = 14'b0000011011011000; // vC= 1752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100010; // iC= 1314 
// vC = 14'b0000010111100100; // vC= 1508 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101010; // iC= 1258 
// vC = 14'b0000011000001010; // vC= 1546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000001; // iC= 1345 
// vC = 14'b0000011010111101; // vC= 1725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000001; // iC= 1281 
// vC = 14'b0000010111101110; // vC= 1518 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001101; // iC= 1357 
// vC = 14'b0000011000100001; // vC= 1569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001010; // iC= 1226 
// vC = 14'b0000011010000010; // vC= 1666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000010; // iC= 1218 
// vC = 14'b0000011001000110; // vC= 1606 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011101; // iC= 1245 
// vC = 14'b0000010111111100; // vC= 1532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111110; // iC= 1022 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011111; // iC= 1119 
// vC = 14'b0000011000011100; // vC= 1564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110011; // iC= 1203 
// vC = 14'b0000011010100011; // vC= 1699 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110000; // iC= 1264 
// vC = 14'b0000011011010010; // vC= 1746 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101010; // iC= 1258 
// vC = 14'b0000011100011110; // vC= 1822 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010011; // iC= 1043 
// vC = 14'b0000011011100101; // vC= 1765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101110; // iC= 1006 
// vC = 14'b0000011010001100; // vC= 1676 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110011; // iC= 1139 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001111; // iC= 1231 
// vC = 14'b0000011001000110; // vC= 1606 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101101; // iC= 1197 
// vC = 14'b0000011000011110; // vC= 1566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100010; // iC= 1250 
// vC = 14'b0000011000101001; // vC= 1577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100011; // iC=  995 
// vC = 14'b0000011010001111; // vC= 1679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110111; // iC= 1207 
// vC = 14'b0000011100110000; // vC= 1840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111100; // iC= 1212 
// vC = 14'b0000011010000010; // vC= 1666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100111; // iC=  999 
// vC = 14'b0000011010111000; // vC= 1720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010001; // iC=  977 
// vC = 14'b0000011101010011; // vC= 1875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101111; // iC=  943 
// vC = 14'b0000011011011110; // vC= 1758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001011; // iC= 1163 
// vC = 14'b0000011010000100; // vC= 1668 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110000; // iC= 1136 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110100; // iC= 1076 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111111; // iC= 1215 
// vC = 14'b0000011101100010; // vC= 1890 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110000; // iC= 1200 
// vC = 14'b0000011001111100; // vC= 1660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100001; // iC= 1185 
// vC = 14'b0000011001011000; // vC= 1624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111100; // iC= 1148 
// vC = 14'b0000011101111101; // vC= 1917 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001001; // iC= 1033 
// vC = 14'b0000011010001011; // vC= 1675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011001; // iC=  985 
// vC = 14'b0000011010011110; // vC= 1694 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101011; // iC= 1067 
// vC = 14'b0000011101000001; // vC= 1857 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000010; // iC= 1154 
// vC = 14'b0000011010111010; // vC= 1722 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111010; // iC= 1082 
// vC = 14'b0000011011110100; // vC= 1780 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010101; // iC= 1045 
// vC = 14'b0000011010111000; // vC= 1720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001101; // iC=  909 
// vC = 14'b0000011011011110; // vC= 1758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101100; // iC= 1132 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110001; // iC=  945 
// vC = 14'b0000011011110111; // vC= 1783 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011111; // iC=  863 
// vC = 14'b0000011111000001; // vC= 1985 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100100; // iC= 1124 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011010; // iC=  986 
// vC = 14'b0000011101000111; // vC= 1863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010001; // iC= 1041 
// vC = 14'b0000011101101100; // vC= 1900 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001111; // iC= 1103 
// vC = 14'b0000011100110010; // vC= 1842 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111110; // iC= 1022 
// vC = 14'b0000011110100011; // vC= 1955 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010010; // iC=  914 
// vC = 14'b0000011010110110; // vC= 1718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100100; // iC=  996 
// vC = 14'b0000011011011110; // vC= 1758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000111; // iC= 1031 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110001; // iC=  945 
// vC = 14'b0000011111010011; // vC= 2003 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100100; // iC=  804 
// vC = 14'b0000011011001010; // vC= 1738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110010; // iC=  946 
// vC = 14'b0000011100010111; // vC= 1815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011101; // iC= 1053 
// vC = 14'b0000011110010111; // vC= 1943 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111100; // iC=  892 
// vC = 14'b0000011011101010; // vC= 1770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101011; // iC=  939 
// vC = 14'b0000011011100011; // vC= 1763 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010110; // iC= 1046 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001000; // iC= 1032 
// vC = 14'b0000011101011000; // vC= 1880 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110010; // iC=  818 
// vC = 14'b0000011011101110; // vC= 1774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000100; // iC=  964 
// vC = 14'b0000011101010101; // vC= 1877 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000000; // iC=  896 
// vC = 14'b0000011101111000; // vC= 1912 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110111010; // iC=  954 
// vC = 14'b0000011011101010; // vC= 1770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010001; // iC=  721 
// vC = 14'b0000011011100111; // vC= 1767 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001111; // iC=  911 
// vC = 14'b0000011110000001; // vC= 1921 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010111; // iC=  983 
// vC = 14'b0000011011011100; // vC= 1756 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011101; // iC=  989 
// vC = 14'b0000100000011100; // vC= 2076 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101100; // iC=  748 
// vC = 14'b0000011011100100; // vC= 1764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001010; // iC=  714 
// vC = 14'b0000011101111100; // vC= 1916 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110001; // iC=  753 
// vC = 14'b0000011101100111; // vC= 1895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010000; // iC=  656 
// vC = 14'b0000011111111000; // vC= 2040 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101001; // iC=  681 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100101000; // iC=  808 
// vC = 14'b0000011111111000; // vC= 2040 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110000; // iC=  624 
// vC = 14'b0000011100011000; // vC= 1816 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000110; // iC=  646 
// vC = 14'b0000100000011000; // vC= 2072 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011011; // iC=  795 
// vC = 14'b0000011100010110; // vC= 1814 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001011; // iC=  779 
// vC = 14'b0000011100010000; // vC= 1808 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001100; // iC=  780 
// vC = 14'b0000011100110111; // vC= 1847 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011101; // iC=  605 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001011; // iC=  779 
// vC = 14'b0000011110001010; // vC= 1930 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011110; // iC=  734 
// vC = 14'b0000011110010110; // vC= 1942 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100010; // iC=  866 
// vC = 14'b0000011100001100; // vC= 1804 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110110; // iC=  566 
// vC = 14'b0000011110111101; // vC= 1981 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111110; // iC=  702 
// vC = 14'b0000100000001010; // vC= 2058 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110011; // iC=  691 
// vC = 14'b0000011100101000; // vC= 1832 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011011; // iC=  795 
// vC = 14'b0000011101011100; // vC= 1884 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010110; // iC=  790 
// vC = 14'b0000011111100010; // vC= 2018 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100000; // iC=  800 
// vC = 14'b0000011110101101; // vC= 1965 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000101; // iC=  645 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001010; // iC=  522 
// vC = 14'b0000011110011000; // vC= 1944 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101101; // iC=  557 
// vC = 14'b0000011110101111; // vC= 1967 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011010; // iC=  666 
// vC = 14'b0000011111010010; // vC= 2002 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111111111; // iC=  511 
// vC = 14'b0000100001100101; // vC= 2149 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000111111; // iC=  575 
// vC = 14'b0000011111011010; // vC= 2010 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110100; // iC=  756 
// vC = 14'b0000011101111101; // vC= 1917 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101110; // iC=  558 
// vC = 14'b0000011101011100; // vC= 1884 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001111; // iC=  591 
// vC = 14'b0000011111100111; // vC= 2023 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110001; // iC=  689 
// vC = 14'b0000011110110011; // vC= 1971 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100010; // iC=  546 
// vC = 14'b0000100001001110; // vC= 2126 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100001; // iC=  609 
// vC = 14'b0000100000010011; // vC= 2067 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000000; // iC=  576 
// vC = 14'b0000100000010101; // vC= 2069 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000000; // iC=  448 
// vC = 14'b0000100000011001; // vC= 2073 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110000; // iC=  496 
// vC = 14'b0000011101010001; // vC= 1873 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001010; // iC=  650 
// vC = 14'b0000100001110011; // vC= 2163 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100000; // iC=  480 
// vC = 14'b0000011101101010; // vC= 1898 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010101; // iC=  341 
// vC = 14'b0000100000011011; // vC= 2075 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101011001; // iC=  345 
// vC = 14'b0000011111100010; // vC= 2018 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011001; // iC=  281 
// vC = 14'b0000100000000110; // vC= 2054 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100001; // iC=  545 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100101; // iC=  549 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000111; // iC=  327 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011001; // iC=  409 
// vC = 14'b0000011110001100; // vC= 1932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111111; // iC=  319 
// vC = 14'b0000011110110000; // vC= 1968 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111010; // iC=  378 
// vC = 14'b0000011110000011; // vC= 1923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101100; // iC=  172 
// vC = 14'b0000100010000101; // vC= 2181 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111100; // iC=  444 
// vC = 14'b0000100001110100; // vC= 2164 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110001000; // iC=  392 
// vC = 14'b0000100001110100; // vC= 2164 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110111; // iC=  183 
// vC = 14'b0000100000100100; // vC= 2084 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001001; // iC=  137 
// vC = 14'b0000011111001111; // vC= 1999 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111010; // iC=  122 
// vC = 14'b0000011111000000; // vC= 1984 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000010; // iC=  322 
// vC = 14'b0000100001001010; // vC= 2122 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001110; // iC=   78 
// vC = 14'b0000100001001010; // vC= 2122 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101111; // iC=  303 
// vC = 14'b0000100000110000; // vC= 2096 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000110111; // iC=   55 
// vC = 14'b0000100001111001; // vC= 2169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111101; // iC=  253 
// vC = 14'b0000011110001001; // vC= 1929 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111110001; // iC=  -15 
// vC = 14'b0000011101111100; // vC= 1916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100010; // iC=  226 
// vC = 14'b0000011110111011; // vC= 1979 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001010001; // iC=   81 
// vC = 14'b0000100010000101; // vC= 2181 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111011; // iC=  -69 
// vC = 14'b0000100000100010; // vC= 2082 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000110111; // iC=   55 
// vC = 14'b0000011111000111; // vC= 1991 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000000011; // iC=    3 
// vC = 14'b0000011110101011; // vC= 1963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000111100; // iC=   60 
// vC = 14'b0000100010000000; // vC= 2176 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011101; // iC=  -99 
// vC = 14'b0000100010000101; // vC= 2181 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110110010; // iC=  -78 
// vC = 14'b0000011101101001; // vC= 1897 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011111; // iC=  -97 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101100; // iC=  -20 
// vC = 14'b0000011110110001; // vC= 1969 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111101; // iC= -131 
// vC = 14'b0000011101110100; // vC= 1908 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010001; // iC=  -47 
// vC = 14'b0000011111010101; // vC= 2005 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010011; // iC= -237 
// vC = 14'b0000011110101111; // vC= 1967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000000; // iC=  -64 
// vC = 14'b0000011111010010; // vC= 2002 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101000100; // iC= -188 
// vC = 14'b0000100001100110; // vC= 2150 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001000; // iC= -184 
// vC = 14'b0000011111001111; // vC= 1999 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100111; // iC= -345 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100001; // iC= -223 
// vC = 14'b0000011110110000; // vC= 1968 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111110; // iC= -386 
// vC = 14'b0000011101011100; // vC= 1884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110101; // iC= -459 
// vC = 14'b0000100000101000; // vC= 2088 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111111; // iC= -449 
// vC = 14'b0000011111011111; // vC= 2015 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000100; // iC= -252 
// vC = 14'b0000100000101001; // vC= 2089 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001110; // iC= -434 
// vC = 14'b0000011101010100; // vC= 1876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000110011; // iC= -461 
// vC = 14'b0000011110111010; // vC= 1978 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001101; // iC= -563 
// vC = 14'b0000011101001101; // vC= 1869 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011001; // iC= -551 
// vC = 14'b0000011101011110; // vC= 1886 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000010; // iC= -446 
// vC = 14'b0000011110101110; // vC= 1966 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101110; // iC= -466 
// vC = 14'b0000011110111001; // vC= 1977 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100110; // iC= -474 
// vC = 14'b0000011110101111; // vC= 1967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100001; // iC= -479 
// vC = 14'b0000011100110101; // vC= 1845 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100010; // iC= -606 
// vC = 14'b0000011110100011; // vC= 1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101001; // iC= -727 
// vC = 14'b0000011110100011; // vC= 1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010101; // iC= -747 
// vC = 14'b0000011101101000; // vC= 1896 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111100; // iC= -644 
// vC = 14'b0000011111001010; // vC= 1994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011101; // iC= -547 
// vC = 14'b0000011100011011; // vC= 1819 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101010; // iC= -662 
// vC = 14'b0000011101110000; // vC= 1904 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011001; // iC= -615 
// vC = 14'b0000011110110010; // vC= 1970 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000011; // iC= -573 
// vC = 14'b0000011100110111; // vC= 1847 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110111; // iC= -649 
// vC = 14'b0000100001000001; // vC= 2113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111101; // iC= -707 
// vC = 14'b0000011100011101; // vC= 1821 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110100; // iC= -780 
// vC = 14'b0000011111010010; // vC= 2002 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101110; // iC= -786 
// vC = 14'b0000011101100010; // vC= 1890 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001001; // iC= -951 
// vC = 14'b0000011100100001; // vC= 1825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100111111; // iC= -705 
// vC = 14'b0000011101101101; // vC= 1901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110100; // iC= -844 
// vC = 14'b0000011110001100; // vC= 1932 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110000; // iC= -912 
// vC = 14'b0000011110100000; // vC= 1952 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111011; // iC= -773 
// vC = 14'b0000011110101111; // vC= 1967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111100; // iC= -964 
// vC = 14'b0000011101101100; // vC= 1900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000010; // iC= -830 
// vC = 14'b0000011110000011; // vC= 1923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b0000011110011001; // vC= 1945 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b0000011100001110; // vC= 1806 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110001; // iC=-1167 
// vC = 14'b0000011100001001; // vC= 1801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100111; // iC=-1049 
// vC = 14'b0000011101000110; // vC= 1862 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101010; // iC=-1238 
// vC = 14'b0000011111011100; // vC= 2012 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100111; // iC=-1049 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001000; // iC=-1016 
// vC = 14'b0000011100110001; // vC= 1841 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001011; // iC=-1141 
// vC = 14'b0000011110111000; // vC= 1976 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001000; // iC=-1272 
// vC = 14'b0000011100110110; // vC= 1846 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110101; // iC=-1099 
// vC = 14'b0000011110010101; // vC= 1941 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001100; // iC=-1140 
// vC = 14'b0000011010111111; // vC= 1727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111111; // iC=-1281 
// vC = 14'b0000011110000001; // vC= 1921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101100; // iC=-1300 
// vC = 14'b0000011100001101; // vC= 1805 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001100; // iC=-1268 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110000; // iC=-1232 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100111; // iC=-1369 
// vC = 14'b0000011100001101; // vC= 1805 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011000; // iC=-1384 
// vC = 14'b0000011010110010; // vC= 1714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101001; // iC=-1239 
// vC = 14'b0000011010010100; // vC= 1684 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011111; // iC=-1377 
// vC = 14'b0000011101100111; // vC= 1895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101100; // iC=-1364 
// vC = 14'b0000011110011111; // vC= 1951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111001; // iC=-1479 
// vC = 14'b0000011101100111; // vC= 1895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001011; // iC=-1269 
// vC = 14'b0000011101011011; // vC= 1883 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110100; // iC=-1356 
// vC = 14'b0000011110100011; // vC= 1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001010; // iC=-1590 
// vC = 14'b0000011101001101; // vC= 1869 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100111; // iC=-1369 
// vC = 14'b0000011100111110; // vC= 1854 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000001; // iC=-1407 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001000; // iC=-1336 
// vC = 14'b0000011100011000; // vC= 1816 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001101; // iC=-1651 
// vC = 14'b0000011101111001; // vC= 1913 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100111; // iC=-1497 
// vC = 14'b0000011001000000; // vC= 1600 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110011; // iC=-1613 
// vC = 14'b0000011011100101; // vC= 1765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110100; // iC=-1612 
// vC = 14'b0000011001000010; // vC= 1602 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010101; // iC=-1707 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100000; // iC=-1504 
// vC = 14'b0000011000101110; // vC= 1582 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000010; // iC=-1470 
// vC = 14'b0000011011100101; // vC= 1765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000101; // iC=-1595 
// vC = 14'b0000011011000111; // vC= 1735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011001; // iC=-1703 
// vC = 14'b0000011100101101; // vC= 1837 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010000; // iC=-1648 
// vC = 14'b0000011010000111; // vC= 1671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110000; // iC=-1680 
// vC = 14'b0000011001101011; // vC= 1643 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110011; // iC=-1613 
// vC = 14'b0000011001001011; // vC= 1611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110101; // iC=-1675 
// vC = 14'b0000010111110011; // vC= 1523 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101001; // iC=-1559 
// vC = 14'b0000011100000101; // vC= 1797 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111011; // iC=-1541 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000001; // iC=-1855 
// vC = 14'b0000011011000101; // vC= 1733 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101011; // iC=-1621 
// vC = 14'b0000011010101011; // vC= 1707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011011; // iC=-1701 
// vC = 14'b0000011011010011; // vC= 1747 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110111; // iC=-1865 
// vC = 14'b0000011010111011; // vC= 1723 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010111; // iC=-1641 
// vC = 14'b0000011001101001; // vC= 1641 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101101; // iC=-1619 
// vC = 14'b0000010111110011; // vC= 1523 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110100; // iC=-1804 
// vC = 14'b0000011010110010; // vC= 1714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011000; // iC=-1768 
// vC = 14'b0000011010101001; // vC= 1705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111000; // iC=-1736 
// vC = 14'b0000011010101011; // vC= 1707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101101; // iC=-1811 
// vC = 14'b0000010110100010; // vC= 1442 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b0000011011000001; // vC= 1729 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000010110000101; // vC= 1413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b0000011011000000; // vC= 1728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000010; // iC=-1726 
// vC = 14'b0000010110000001; // vC= 1409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000110; // iC=-1786 
// vC = 14'b0000011001010000; // vC= 1616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b0000011010010011; // vC= 1683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b0000010111111000; // vC= 1528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011001; // iC=-1767 
// vC = 14'b0000011001110110; // vC= 1654 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011010; // iC=-2022 
// vC = 14'b0000011001011100; // vC= 1628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b0000011000101000; // vC= 1576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001110; // iC=-1906 
// vC = 14'b0000011001110111; // vC= 1655 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b0000011000100011; // vC= 1571 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100110; // iC=-1818 
// vC = 14'b0000011000101000; // vC= 1576 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111101; // iC=-1859 
// vC = 14'b0000010111111011; // vC= 1531 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b0000010101011110; // vC= 1374 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001110; // iC=-2034 
// vC = 14'b0000011000011111; // vC= 1567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011010; // iC=-1894 
// vC = 14'b0000010111111001; // vC= 1529 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000100; // iC=-1916 
// vC = 14'b0000010110110011; // vC= 1459 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000000; // iC=-1920 
// vC = 14'b0000010110000110; // vC= 1414 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000010101101010; // vC= 1386 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100110; // iC=-1818 
// vC = 14'b0000011000011100; // vC= 1564 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110010; // iC=-1870 
// vC = 14'b0000010110011100; // vC= 1436 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100110; // iC=-1882 
// vC = 14'b0000010100001100; // vC= 1292 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b0000010011101110; // vC= 1262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010010; // iC=-2094 
// vC = 14'b0000010101011101; // vC= 1373 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b0000010100010110; // vC= 1302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b0000010111010000; // vC= 1488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000010011111000; // vC= 1272 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b0000010100001110; // vC= 1294 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b0000010110111100; // vC= 1468 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000010010101100; // vC= 1196 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b0000010011000110; // vC= 1222 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000010; // iC=-1918 
// vC = 14'b0000010110000110; // vC= 1414 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b0000010001110000; // vC= 1136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100101; // iC=-2075 
// vC = 14'b0000010110001011; // vC= 1419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000110; // iC=-2106 
// vC = 14'b0000010101110001; // vC= 1393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101001; // iC=-2071 
// vC = 14'b0000010101101001; // vC= 1385 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b0000010001100001; // vC= 1121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010100; // iC=-1964 
// vC = 14'b0000010101010011; // vC= 1363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100101; // iC=-2011 
// vC = 14'b0000010100000100; // vC= 1284 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b0000010000111110; // vC= 1086 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011001; // iC=-2087 
// vC = 14'b0000010000110110; // vC= 1078 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101010; // iC=-2134 
// vC = 14'b0000010100011010; // vC= 1306 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b0000010011110100; // vC= 1268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111111; // iC=-1985 
// vC = 14'b0000010000111101; // vC= 1085 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110011; // iC=-1997 
// vC = 14'b0000010011010111; // vC= 1239 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100001; // iC=-2143 
// vC = 14'b0000010010101001; // vC= 1193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b0000010010101001; // vC= 1193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000001; // iC=-1983 
// vC = 14'b0000010000000100; // vC= 1028 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b0000001111100000; // vC=  992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110100; // iC=-2124 
// vC = 14'b0000010010101111; // vC= 1199 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b0000010000101101; // vC= 1069 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000111; // iC=-1977 
// vC = 14'b0000010000000001; // vC= 1025 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b0000001111011001; // vC=  985 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000010010101011; // vC= 1195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b0000010011000111; // vC= 1223 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000010000011100; // vC= 1052 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b0000010000111011; // vC= 1083 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010011; // iC=-2221 
// vC = 14'b0000010010110000; // vC= 1200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b0000010000000001; // vC= 1025 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000001110010100; // vC=  916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010011; // iC=-2221 
// vC = 14'b0000010010011011; // vC= 1179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b0000001111101111; // vC= 1007 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001001; // iC=-2103 
// vC = 14'b0000010000000001; // vC= 1025 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010100; // iC=-2092 
// vC = 14'b0000001110001001; // vC=  905 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b0000001111100111; // vC=  999 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101001; // iC=-2007 
// vC = 14'b0000001101010000; // vC=  848 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101111; // iC=-1937 
// vC = 14'b0000001101100001; // vC=  865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b0000001111010111; // vC=  983 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b0000001110111001; // vC=  953 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110001; // iC=-1999 
// vC = 14'b0000001110101001; // vC=  937 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b0000010000101110; // vC= 1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010101; // iC=-2091 
// vC = 14'b0000010000011110; // vC= 1054 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001111; // iC=-2097 
// vC = 14'b0000010000101110; // vC= 1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000001101011010; // vC=  858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011101; // iC=-2211 
// vC = 14'b0000001111111100; // vC= 1020 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000001110010111; // vC=  919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011101; // iC=-2019 
// vC = 14'b0000001011011000; // vC=  728 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001101; // iC=-2035 
// vC = 14'b0000001100101011; // vC=  811 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010000; // iC=-2160 
// vC = 14'b0000001101100000; // vC=  864 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b0000001011110101; // vC=  757 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b0000001100100011; // vC=  803 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110000; // iC=-2256 
// vC = 14'b0000001101011101; // vC=  861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101010; // iC=-2134 
// vC = 14'b0000001100100111; // vC=  807 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111100; // iC=-2116 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b0000001100010010; // vC=  786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100000; // iC=-1952 
// vC = 14'b0000001011000110; // vC=  710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000000; // iC=-2176 
// vC = 14'b0000001101101000; // vC=  872 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b0000001101000111; // vC=  839 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000111; // iC=-1977 
// vC = 14'b0000001011101111; // vC=  751 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001001; // iC=-2167 
// vC = 14'b0000001010011111; // vC=  671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001010; // iC=-2230 
// vC = 14'b0000001100100111; // vC=  807 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b0000001001100111; // vC=  615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b0000001101101000; // vC=  872 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100000; // iC=-2080 
// vC = 14'b0000001100000110; // vC=  774 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100000; // iC=-1952 
// vC = 14'b0000001100101011; // vC=  811 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000001100111001; // vC=  825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000001; // iC=-2175 
// vC = 14'b0000001001111001; // vC=  633 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100100111; // iC=-2265 
// vC = 14'b0000001010000011; // vC=  643 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010110; // iC=-2026 
// vC = 14'b0000001001110100; // vC=  628 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000001; // iC=-1983 
// vC = 14'b0000001011010101; // vC=  725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111110; // iC=-2242 
// vC = 14'b0000000111110110; // vC=  502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b0000001000101010; // vC=  554 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111100; // iC=-2180 
// vC = 14'b0000001100010100; // vC=  788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000001011011110; // vC=  734 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b0000000111011000; // vC=  472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011000; // iC=-2152 
// vC = 14'b0000001001101101; // vC=  621 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001111; // iC=-2161 
// vC = 14'b0000001000100110; // vC=  550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111011; // iC=-2245 
// vC = 14'b0000000111111010; // vC=  506 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011000; // iC=-2216 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010001; // iC=-2223 
// vC = 14'b0000001001110111; // vC=  631 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b0000001010111101; // vC=  701 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100111; // iC=-2009 
// vC = 14'b0000001000110001; // vC=  561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100011; // iC=-2141 
// vC = 14'b0000000110010001; // vC=  401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b0000001001000001; // vC=  577 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000110; // iC=-2042 
// vC = 14'b0000001000001011; // vC=  523 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011001; // iC=-2087 
// vC = 14'b0000000111011100; // vC=  476 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000100; // iC=-2172 
// vC = 14'b0000000111001000; // vC=  456 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010111; // iC=-2025 
// vC = 14'b0000000111100000; // vC=  480 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b0000001000101000; // vC=  552 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100000; // iC=-2208 
// vC = 14'b0000001000010001; // vC=  529 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101011; // iC=-2133 
// vC = 14'b0000001000000100; // vC=  516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011101; // iC=-2083 
// vC = 14'b0000000111111110; // vC=  510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100110; // iC=-2074 
// vC = 14'b0000000110001110; // vC=  398 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011101; // iC=-2211 
// vC = 14'b0000000110010100; // vC=  404 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011101; // iC=-2147 
// vC = 14'b0000000110111101; // vC=  445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011001; // iC=-2151 
// vC = 14'b0000001000000100; // vC=  516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b0000000111011010; // vC=  474 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b0000000110100101; // vC=  421 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111111; // iC=-2049 
// vC = 14'b0000000101100010; // vC=  354 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011011; // iC=-2085 
// vC = 14'b0000001000011001; // vC=  537 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111010; // iC=-2246 
// vC = 14'b0000000110011111; // vC=  415 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b0000000110010010; // vC=  402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000000110101111; // vC=  431 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100011101; // iC=-2275 
// vC = 14'b0000000101010101; // vC=  341 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000001000000010; // vC=  514 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000001; // iC=-2175 
// vC = 14'b0000000011010100; // vC=  212 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010011; // iC=-2093 
// vC = 14'b0000000110110111; // vC=  439 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101110; // iC=-2130 
// vC = 14'b0000000011010010; // vC=  210 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b0000000011001010; // vC=  202 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001111; // iC=-2097 
// vC = 14'b0000000010010011; // vC=  147 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111111; // iC=-2049 
// vC = 14'b0000000110101000; // vC=  424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010100; // iC=-2156 
// vC = 14'b0000000011101000; // vC=  232 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010000; // iC=-1968 
// vC = 14'b0000000100110101; // vC=  309 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000010; // iC=-2174 
// vC = 14'b0000000110010100; // vC=  404 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001000; // iC=-2232 
// vC = 14'b0000000010101000; // vC=  168 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b0000000100111101; // vC=  317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b0000000101010100; // vC=  340 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000000011100000; // vC=  224 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111000; // iC=-2056 
// vC = 14'b0000000010001101; // vC=  141 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010010; // iC=-2222 
// vC = 14'b0000000100100011; // vC=  291 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110010; // iC=-2254 
// vC = 14'b0000000101000110; // vC=  326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b0000000001110110; // vC=  118 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101010; // iC=-2070 
// vC = 14'b0000000010001000; // vC=  136 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011011; // iC=-2213 
// vC = 14'b0000000100111110; // vC=  318 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010110; // iC=-2154 
// vC = 14'b0000000011001011; // vC=  203 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b0000000010101001; // vC=  169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000111; // iC=-2105 
// vC = 14'b0000000010011000; // vC=  152 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000000010000000; // vC=  128 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000100; // iC=-1980 
// vC = 14'b0000000100000101; // vC=  261 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100101; // iC=-2075 
// vC = 14'b0000000001111100; // vC=  124 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111111; // iC=-2049 
// vC = 14'b0000000000011100; // vC=   28 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b0000000001010110; // vC=   86 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b0000000010100001; // vC=  161 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111000; // iC=-2184 
// vC = 14'b0000000010111001; // vC=  185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b0000000011011000; // vC=  216 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000110; // iC=-2106 
// vC = 14'b0000000011100000; // vC=  224 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b1111111111001101; // vC=  -51 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100111; // iC=-2073 
// vC = 14'b0000000011001001; // vC=  201 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b1111111110100110; // vC=  -90 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000011; // iC=-2045 
// vC = 14'b1111111111000101; // vC=  -59 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b1111111101111011; // vC= -133 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010001; // iC=-2223 
// vC = 14'b0000000000101011; // vC=   43 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101001; // iC=-2007 
// vC = 14'b1111111101101000; // vC= -152 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000011; // iC=-2237 
// vC = 14'b1111111110011001; // vC= -103 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011110; // iC=-2210 
// vC = 14'b0000000001100010; // vC=   98 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b0000000001111101; // vC=  125 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b1111111111010011; // vC=  -45 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011101; // iC=-2211 
// vC = 14'b1111111110111001; // vC=  -71 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011110; // iC=-2210 
// vC = 14'b1111111101101110; // vC= -146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000100; // iC=-1916 
// vC = 14'b1111111111111010; // vC=   -6 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b1111111110001011; // vC= -117 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b1111111111010011; // vC=  -45 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011111; // iC=-2081 
// vC = 14'b1111111111010101; // vC=  -43 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000110; // iC=-2170 
// vC = 14'b1111111110000111; // vC= -121 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111000; // iC=-2120 
// vC = 14'b1111111101001101; // vC= -179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b1111111111100100; // vC=  -28 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b1111111110110111; // vC=  -73 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b1111111101100011; // vC= -157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b1111111011111010; // vC= -262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000101; // iC=-2107 
// vC = 14'b1111111011011000; // vC= -296 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010001; // iC=-2031 
// vC = 14'b1111111111011111; // vC=  -33 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001010; // iC=-2166 
// vC = 14'b1111111101011011; // vC= -165 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101100; // iC=-2196 
// vC = 14'b1111111101001101; // vC= -179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100110; // iC=-2138 
// vC = 14'b1111111010111101; // vC= -323 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010111; // iC=-2025 
// vC = 14'b1111111100100000; // vC= -224 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b1111111101110110; // vC= -138 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b1111111100101011; // vC= -213 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011110; // iC=-2146 
// vC = 14'b1111111101101010; // vC= -150 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b1111111100000100; // vC= -252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100011; // iC=-2141 
// vC = 14'b1111111110011110; // vC=  -98 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101101; // iC=-2067 
// vC = 14'b1111111100101100; // vC= -212 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b1111111110100100; // vC=  -92 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100001; // iC=-2143 
// vC = 14'b1111111011100001; // vC= -287 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000001; // iC=-1983 
// vC = 14'b1111111011001000; // vC= -312 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b1111111110001000; // vC= -120 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111001; // iC=-1991 
// vC = 14'b1111111011011101; // vC= -291 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100101; // iC=-2011 
// vC = 14'b1111111100000100; // vC= -252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b1111111011000111; // vC= -313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001101; // iC=-1907 
// vC = 14'b1111111011111010; // vC= -262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110000; // iC=-2128 
// vC = 14'b1111111010010100; // vC= -364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100000; // iC=-2080 
// vC = 14'b1111111001100111; // vC= -409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b1111111010011000; // vC= -360 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110010; // iC=-1870 
// vC = 14'b1111111000001011; // vC= -501 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010101; // iC=-2091 
// vC = 14'b1111111100010010; // vC= -238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100111; // iC=-1881 
// vC = 14'b1111111000010100; // vC= -492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b1111111011110011; // vC= -269 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000000; // iC=-1856 
// vC = 14'b1111111011110101; // vC= -267 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b1111111000111110; // vC= -450 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000001; // iC=-1919 
// vC = 14'b1111111011101011; // vC= -277 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b1111111010011001; // vC= -359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110011; // iC=-1933 
// vC = 14'b1111110111100000; // vC= -544 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b1111111010011001; // vC= -359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b1111111001111001; // vC= -391 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b1111111001011100; // vC= -420 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b1111111010111001; // vC= -327 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b1111111001101111; // vC= -401 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110001; // iC=-2127 
// vC = 14'b1111111001101110; // vC= -402 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b1111111001110100; // vC= -396 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b1111111011000000; // vC= -320 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101100; // iC=-1876 
// vC = 14'b1111111000111010; // vC= -454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010110; // iC=-2090 
// vC = 14'b1111110110010110; // vC= -618 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001011; // iC=-1973 
// vC = 14'b1111111000100110; // vC= -474 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b1111110101101010; // vC= -662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011101; // iC=-1827 
// vC = 14'b1111111000100010; // vC= -478 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100111; // iC=-2073 
// vC = 14'b1111111010001111; // vC= -369 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001101; // iC=-2099 
// vC = 14'b1111111001111011; // vC= -389 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b1111110111011000; // vC= -552 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100011; // iC=-1821 
// vC = 14'b1111111000111101; // vC= -451 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101110; // iC=-1810 
// vC = 14'b1111111001101011; // vC= -405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010011; // iC=-2093 
// vC = 14'b1111110111001000; // vC= -568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001001; // iC=-2039 
// vC = 14'b1111111000100011; // vC= -477 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b1111110101111111; // vC= -641 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b1111110111110011; // vC= -525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101001; // iC=-2071 
// vC = 14'b1111110101010110; // vC= -682 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b1111111000011000; // vC= -488 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011100; // iC=-1956 
// vC = 14'b1111111000100100; // vC= -476 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b1111110101011001; // vC= -679 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101101; // iC=-1939 
// vC = 14'b1111110011110001; // vC= -783 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111011; // iC=-1861 
// vC = 14'b1111110101110101; // vC= -651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b1111111000010111; // vC= -489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110001; // iC=-1807 
// vC = 14'b1111110100111110; // vC= -706 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001100; // iC=-1908 
// vC = 14'b1111110110100110; // vC= -602 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b1111110111100001; // vC= -543 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101010; // iC=-1750 
// vC = 14'b1111110110010010; // vC= -622 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b1111110101001101; // vC= -691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111110011010001; // vC= -815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100111; // iC=-2009 
// vC = 14'b1111110101110010; // vC= -654 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101000; // iC=-1752 
// vC = 14'b1111110011001100; // vC= -820 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111001; // iC=-1735 
// vC = 14'b1111110100110101; // vC= -715 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b1111110100101100; // vC= -724 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010111; // iC=-1705 
// vC = 14'b1111110011000001; // vC= -831 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111111; // iC=-1729 
// vC = 14'b1111110010000111; // vC= -889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b1111110110110001; // vC= -591 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b1111110100011001; // vC= -743 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011111; // iC=-1889 
// vC = 14'b1111110110011100; // vC= -612 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000000; // iC=-1856 
// vC = 14'b1111110110010010; // vC= -622 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110001; // iC=-1743 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001100; // iC=-1780 
// vC = 14'b1111110101001001; // vC= -695 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001000; // iC=-1720 
// vC = 14'b1111110100001101; // vC= -755 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001101; // iC=-1907 
// vC = 14'b1111110001011110; // vC= -930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110001; // iC=-1743 
// vC = 14'b1111110101010101; // vC= -683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b1111110010101101; // vC= -851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111101; // iC=-1859 
// vC = 14'b1111110011101000; // vC= -792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b1111110101011011; // vC= -677 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b1111110101000101; // vC= -699 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101010; // iC=-1750 
// vC = 14'b1111110000111001; // vC= -967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000110; // iC=-1850 
// vC = 14'b1111110001101011; // vC= -917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111001; // iC=-1927 
// vC = 14'b1111110001111101; // vC= -899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010110; // iC=-1898 
// vC = 14'b1111110100110100; // vC= -716 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000111; // iC=-1657 
// vC = 14'b1111110000001011; // vC=-1013 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111100; // iC=-1860 
// vC = 14'b1111110010110111; // vC= -841 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010110; // iC=-1770 
// vC = 14'b1111110011100010; // vC= -798 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010101; // iC=-1835 
// vC = 14'b1111110010010011; // vC= -877 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010001; // iC=-1647 
// vC = 14'b1111110011000110; // vC= -826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010111; // iC=-1641 
// vC = 14'b1111110000100000; // vC= -992 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101001; // iC=-1815 
// vC = 14'b1111110011101101; // vC= -787 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010111; // iC=-1769 
// vC = 14'b1111101110111110; // vC=-1090 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111101; // iC=-1667 
// vC = 14'b1111110001101000; // vC= -920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100011; // iC=-1693 
// vC = 14'b1111110011010000; // vC= -816 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b1111110000111011; // vC= -965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000010; // iC=-1598 
// vC = 14'b1111110000101111; // vC= -977 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100101; // iC=-1755 
// vC = 14'b1111101111111011; // vC=-1029 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110010; // iC=-1614 
// vC = 14'b1111110001000000; // vC= -960 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001010; // iC=-1590 
// vC = 14'b1111110001001001; // vC= -951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010000; // iC=-1776 
// vC = 14'b1111101111111010; // vC=-1030 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101111; // iC=-1809 
// vC = 14'b1111110010110001; // vC= -847 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111100; // iC=-1860 
// vC = 14'b1111110000110100; // vC= -972 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110011; // iC=-1741 
// vC = 14'b1111110010100001; // vC= -863 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011111; // iC=-1569 
// vC = 14'b1111101111011110; // vC=-1058 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100001; // iC=-1823 
// vC = 14'b1111110001000111; // vC= -953 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100000; // iC=-1696 
// vC = 14'b1111110000110101; // vC= -971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111001; // iC=-1671 
// vC = 14'b1111110001010011; // vC= -941 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111001; // iC=-1671 
// vC = 14'b1111110001100010; // vC= -926 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100111; // iC=-1625 
// vC = 14'b1111101111001111; // vC=-1073 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100101; // iC=-1627 
// vC = 14'b1111101101001110; // vC=-1202 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000000; // iC=-1536 
// vC = 14'b1111110001000101; // vC= -955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111000; // iC=-1736 
// vC = 14'b1111110001011011; // vC= -933 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101100; // iC=-1748 
// vC = 14'b1111110000101000; // vC= -984 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011010; // iC=-1766 
// vC = 14'b1111110000001010; // vC=-1014 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011110; // iC=-1826 
// vC = 14'b1111101100001101; // vC=-1267 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000111; // iC=-1721 
// vC = 14'b1111101111010010; // vC=-1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100011; // iC=-1821 
// vC = 14'b1111110000001010; // vC=-1014 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100001; // iC=-1631 
// vC = 14'b1111101011111100; // vC=-1284 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010100; // iC=-1772 
// vC = 14'b1111101101101011; // vC=-1173 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110001; // iC=-1551 
// vC = 14'b1111101110111110; // vC=-1090 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011101; // iC=-1635 
// vC = 14'b1111101100001010; // vC=-1270 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010000; // iC=-1776 
// vC = 14'b1111101101111000; // vC=-1160 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001100; // iC=-1524 
// vC = 14'b1111101101110011; // vC=-1165 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101111; // iC=-1489 
// vC = 14'b1111101101000001; // vC=-1215 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011110; // iC=-1634 
// vC = 14'b1111101111000010; // vC=-1086 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000000; // iC=-1536 
// vC = 14'b1111101111100100; // vC=-1052 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101001; // iC=-1751 
// vC = 14'b1111101101100011; // vC=-1181 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011100; // iC=-1764 
// vC = 14'b1111101110011001; // vC=-1127 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001110; // iC=-1522 
// vC = 14'b1111101110100100; // vC=-1116 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000010; // iC=-1470 
// vC = 14'b1111101010110101; // vC=-1355 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000111; // iC=-1721 
// vC = 14'b1111101101110000; // vC=-1168 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010110; // iC=-1642 
// vC = 14'b1111101110011010; // vC=-1126 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000010; // iC=-1726 
// vC = 14'b1111101110101110; // vC=-1106 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011101; // iC=-1507 
// vC = 14'b1111101010001101; // vC=-1395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001110; // iC=-1714 
// vC = 14'b1111101110101101; // vC=-1107 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100011; // iC=-1693 
// vC = 14'b1111101110110001; // vC=-1103 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010011; // iC=-1517 
// vC = 14'b1111101100001101; // vC=-1267 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101001; // iC=-1431 
// vC = 14'b1111101011000110; // vC=-1338 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110111; // iC=-1545 
// vC = 14'b1111101100101110; // vC=-1234 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001001; // iC=-1655 
// vC = 14'b1111101100000000; // vC=-1280 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110110; // iC=-1610 
// vC = 14'b1111101100001001; // vC=-1271 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010101; // iC=-1707 
// vC = 14'b1111101010000100; // vC=-1404 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011010; // iC=-1574 
// vC = 14'b1111101001101100; // vC=-1428 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111110; // iC=-1410 
// vC = 14'b1111101001101000; // vC=-1432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000010; // iC=-1598 
// vC = 14'b1111101011111101; // vC=-1283 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111001; // iC=-1415 
// vC = 14'b1111101010101010; // vC=-1366 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100101; // iC=-1371 
// vC = 14'b1111101010010001; // vC=-1391 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110010; // iC=-1486 
// vC = 14'b1111101101010010; // vC=-1198 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000110; // iC=-1530 
// vC = 14'b1111101100001001; // vC=-1271 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101101; // iC=-1555 
// vC = 14'b1111101100101000; // vC=-1240 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101111; // iC=-1617 
// vC = 14'b1111101101001001; // vC=-1207 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111111; // iC=-1537 
// vC = 14'b1111101101011011; // vC=-1189 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110001; // iC=-1423 
// vC = 14'b1111101000111111; // vC=-1473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011101; // iC=-1379 
// vC = 14'b1111101101010000; // vC=-1200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100101; // iC=-1499 
// vC = 14'b1111101010110010; // vC=-1358 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001000; // iC=-1400 
// vC = 14'b1111101100111001; // vC=-1223 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111111; // iC=-1345 
// vC = 14'b1111101001100001; // vC=-1439 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000010; // iC=-1534 
// vC = 14'b1111101000100111; // vC=-1497 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011011; // iC=-1509 
// vC = 14'b1111101000011011; // vC=-1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110011; // iC=-1421 
// vC = 14'b1111101000110100; // vC=-1484 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000111; // iC=-1337 
// vC = 14'b1111101000111110; // vC=-1474 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000000; // iC=-1344 
// vC = 14'b1111100111101001; // vC=-1559 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010111; // iC=-1449 
// vC = 14'b1111101010101001; // vC=-1367 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010001; // iC=-1583 
// vC = 14'b1111101001111111; // vC=-1409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110010; // iC=-1486 
// vC = 14'b1111101001001010; // vC=-1462 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101101; // iC=-1299 
// vC = 14'b1111101010000011; // vC=-1405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101001; // iC=-1303 
// vC = 14'b1111101011110111; // vC=-1289 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001011; // iC=-1397 
// vC = 14'b1111101011111001; // vC=-1287 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011001; // iC=-1255 
// vC = 14'b1111100111001100; // vC=-1588 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110111; // iC=-1417 
// vC = 14'b1111101000010010; // vC=-1518 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101010; // iC=-1430 
// vC = 14'b1111100110111111; // vC=-1601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111000; // iC=-1480 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111111; // iC=-1281 
// vC = 14'b1111100110111000; // vC=-1608 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011110; // iC=-1378 
// vC = 14'b1111100111110101; // vC=-1547 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111000; // iC=-1352 
// vC = 14'b1111101001110101; // vC=-1419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100101; // iC=-1371 
// vC = 14'b1111100110101101; // vC=-1619 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010111; // iC=-1385 
// vC = 14'b1111101010000010; // vC=-1406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010111; // iC=-1385 
// vC = 14'b1111101010011111; // vC=-1377 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110111; // iC=-1289 
// vC = 14'b1111100110110011; // vC=-1613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111001; // iC=-1223 
// vC = 14'b1111101001111000; // vC=-1416 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011000; // iC=-1320 
// vC = 14'b1111101001100101; // vC=-1435 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000110100; // iC=-1484 
// vC = 14'b1111101000110101; // vC=-1483 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000111; // iC=-1273 
// vC = 14'b1111101001101101; // vC=-1427 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101011; // iC=-1493 
// vC = 14'b1111100111110010; // vC=-1550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000010; // iC=-1342 
// vC = 14'b1111100111000011; // vC=-1597 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000000; // iC=-1280 
// vC = 14'b1111101001000101; // vC=-1467 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010001; // iC=-1327 
// vC = 14'b1111101000001010; // vC=-1526 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100001; // iC=-1375 
// vC = 14'b1111101010001010; // vC=-1398 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100011; // iC=-1181 
// vC = 14'b1111100111000001; // vC=-1599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001100; // iC=-1460 
// vC = 14'b1111101000011100; // vC=-1508 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011111; // iC=-1249 
// vC = 14'b1111100111100111; // vC=-1561 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001000; // iC=-1272 
// vC = 14'b1111100111101010; // vC=-1558 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110111; // iC=-1225 
// vC = 14'b1111100110000111; // vC=-1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110110; // iC=-1354 
// vC = 14'b1111100111100010; // vC=-1566 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101101; // iC=-1363 
// vC = 14'b1111100101111000; // vC=-1672 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101010; // iC=-1238 
// vC = 14'b1111100101000001; // vC=-1727 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111001; // iC=-1159 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011001; // iC=-1127 
// vC = 14'b1111100110011010; // vC=-1638 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001100; // iC=-1396 
// vC = 14'b1111101001000001; // vC=-1471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000100; // iC=-1404 
// vC = 14'b1111100101111000; // vC=-1672 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100101; // iC=-1307 
// vC = 14'b1111100110110000; // vC=-1616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101010; // iC=-1366 
// vC = 14'b1111101000111110; // vC=-1474 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110100; // iC=-1356 
// vC = 14'b1111100110011111; // vC=-1633 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111100; // iC=-1284 
// vC = 14'b1111100111001011; // vC=-1589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111110; // iC=-1282 
// vC = 14'b1111100111111011; // vC=-1541 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011000; // iC=-1256 
// vC = 14'b1111100111010101; // vC=-1579 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000111; // iC=-1273 
// vC = 14'b1111100111111111; // vC=-1537 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000110; // iC=-1274 
// vC = 14'b1111100110101001; // vC=-1623 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000101; // iC=-1147 
// vC = 14'b1111100110001100; // vC=-1652 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110100; // iC=-1228 
// vC = 14'b1111100110100000; // vC=-1632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011010; // iC=-1126 
// vC = 14'b1111100101111100; // vC=-1668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111111; // iC=-1089 
// vC = 14'b1111100111010001; // vC=-1583 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110011; // iC=-1101 
// vC = 14'b1111100110000000; // vC=-1664 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111011; // iC=-1221 
// vC = 14'b1111101000001011; // vC=-1525 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011110; // iC=-1314 
// vC = 14'b1111100100100100; // vC=-1756 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111010; // iC=-1094 
// vC = 14'b1111100110110001; // vC=-1615 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010011; // iC=-1197 
// vC = 14'b1111100111001111; // vC=-1585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110011; // iC=-1229 
// vC = 14'b1111100010111100; // vC=-1860 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110110; // iC=-1226 
// vC = 14'b1111100100010001; // vC=-1775 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010000; // iC=-1264 
// vC = 14'b1111100111011101; // vC=-1571 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010101; // iC=-1067 
// vC = 14'b1111100110101111; // vC=-1617 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101001; // iC= -983 
// vC = 14'b1111100101011100; // vC=-1700 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010000; // iC=-1136 
// vC = 14'b1111100101010100; // vC=-1708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110111; // iC=-1161 
// vC = 14'b1111100111000111; // vC=-1593 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101111001; // iC=-1159 
// vC = 14'b1111100011011101; // vC=-1827 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011111; // iC= -993 
// vC = 14'b1111100110001110; // vC=-1650 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010000; // iC= -944 
// vC = 14'b1111100110000111; // vC=-1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001000; // iC= -952 
// vC = 14'b1111100010101000; // vC=-1880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101011; // iC= -917 
// vC = 14'b1111100110100000; // vC=-1632 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010011; // iC=-1133 
// vC = 14'b1111100110101100; // vC=-1620 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010010; // iC= -942 
// vC = 14'b1111100110000001; // vC=-1663 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000000; // iC= -896 
// vC = 14'b1111100110011100; // vC=-1636 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000010; // iC=-1086 
// vC = 14'b1111100100111101; // vC=-1731 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011010; // iC=-1190 
// vC = 14'b1111100010101011; // vC=-1877 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000011; // iC=-1149 
// vC = 14'b1111100010100111; // vC=-1881 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100100; // iC=-1180 
// vC = 14'b1111100100001001; // vC=-1783 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000011; // iC=-1149 
// vC = 14'b1111100010011111; // vC=-1889 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110110; // iC=-1098 
// vC = 14'b1111100110001101; // vC=-1651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001110; // iC= -882 
// vC = 14'b1111100001101110; // vC=-1938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001001; // iC=-1079 
// vC = 14'b1111100011000101; // vC=-1851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010000; // iC= -944 
// vC = 14'b1111100101001101; // vC=-1715 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010100; // iC= -876 
// vC = 14'b1111100101100111; // vC=-1689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100011; // iC=-1053 
// vC = 14'b1111100101000110; // vC=-1722 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110000; // iC=-1040 
// vC = 14'b1111100100011011; // vC=-1765 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000111; // iC=-1081 
// vC = 14'b1111100001101110; // vC=-1938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110011101; // iC=-1123 
// vC = 14'b1111100011101010; // vC=-1814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010100; // iC= -876 
// vC = 14'b1111100011101010; // vC=-1814 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001100; // iC= -948 
// vC = 14'b1111100101101100; // vC=-1684 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010100; // iC=-1068 
// vC = 14'b1111100101110010; // vC=-1678 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001101; // iC=-1075 
// vC = 14'b1111100011011011; // vC=-1829 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000010; // iC= -958 
// vC = 14'b1111100011010100; // vC=-1836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010110; // iC= -938 
// vC = 14'b1111100101011111; // vC=-1697 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011111; // iC=-1057 
// vC = 14'b1111100001111111; // vC=-1921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001011011; // iC= -933 
// vC = 14'b1111100000100110; // vC=-2010 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110111; // iC= -905 
// vC = 14'b1111100100000001; // vC=-1791 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011100; // iC=-1060 
// vC = 14'b1111100000100111; // vC=-2009 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100001; // iC= -735 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110011; // iC=-1037 
// vC = 14'b1111100011110001; // vC=-1807 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110110; // iC=-1034 
// vC = 14'b1111100100001110; // vC=-1778 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001001101; // iC= -947 
// vC = 14'b1111100100000000; // vC=-1792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110101; // iC= -907 
// vC = 14'b1111100000001100; // vC=-2036 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000010; // iC= -958 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000011; // iC= -829 
// vC = 14'b1111100100010001; // vC=-1775 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111101; // iC= -771 
// vC = 14'b1111100100101111; // vC=-1745 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100011; // iC= -861 
// vC = 14'b1111100001101110; // vC=-1938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111000; // iC= -776 
// vC = 14'b1111100001110001; // vC=-1935 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111011; // iC= -837 
// vC = 14'b1111100000100101; // vC=-2011 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111000; // iC= -904 
// vC = 14'b1111011111110000; // vC=-2064 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100100; // iC= -796 
// vC = 14'b1111100001011001; // vC=-1959 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101010; // iC= -790 
// vC = 14'b1111100001010101; // vC=-1963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011111; // iC= -737 
// vC = 14'b1111011111101000; // vC=-2072 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110011; // iC= -845 
// vC = 14'b1111100011000011; // vC=-1853 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101001; // iC= -663 
// vC = 14'b1111100000110101; // vC=-1995 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110101; // iC= -715 
// vC = 14'b1111100001000010; // vC=-1982 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000010; // iC= -766 
// vC = 14'b1111100100011100; // vC=-1764 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100110; // iC= -730 
// vC = 14'b1111100011100001; // vC=-1823 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100000011; // iC= -765 
// vC = 14'b1111011111011000; // vC=-2088 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100110; // iC= -666 
// vC = 14'b1111100000100010; // vC=-2014 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100010; // iC= -862 
// vC = 14'b1111100100010010; // vC=-1774 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110011; // iC= -653 
// vC = 14'b1111100001110110; // vC=-1930 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001010; // iC= -758 
// vC = 14'b1111100000110111; // vC=-1993 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100101; // iC= -795 
// vC = 14'b1111100001110111; // vC=-1929 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001110; // iC= -818 
// vC = 14'b1111100011100100; // vC=-1820 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110101; // iC= -651 
// vC = 14'b1111100001110000; // vC=-1936 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010011; // iC= -749 
// vC = 14'b1111011111011111; // vC=-2081 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110011; // iC= -653 
// vC = 14'b1111011111101000; // vC=-2072 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001001; // iC= -567 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001111; // iC= -561 
// vC = 14'b1111100001010011; // vC=-1965 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001100; // iC= -756 
// vC = 14'b1111011111000100; // vC=-2108 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111100; // iC= -644 
// vC = 14'b1111100011011001; // vC=-1831 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110101; // iC= -779 
// vC = 14'b1111011111000010; // vC=-2110 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101001; // iC= -727 
// vC = 14'b1111100010000011; // vC=-1917 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100010; // iC= -734 
// vC = 14'b1111100010001100; // vC=-1908 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000010; // iC= -574 
// vC = 14'b1111100000100011; // vC=-2013 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001101; // iC= -563 
// vC = 14'b1111011111101010; // vC=-2070 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111110; // iC= -514 
// vC = 14'b1111100000001110; // vC=-2034 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010111; // iC= -745 
// vC = 14'b1111100001010110; // vC=-1962 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111100; // iC= -580 
// vC = 14'b1111100010000110; // vC=-1914 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010100; // iC= -684 
// vC = 14'b1111100000110110; // vC=-1994 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100011; // iC= -669 
// vC = 14'b1111100000000010; // vC=-2046 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000000100; // iC= -508 
// vC = 14'b1111100000111010; // vC=-1990 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100010; // iC= -606 
// vC = 14'b1111100011010111; // vC=-1833 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110000001; // iC= -639 
// vC = 14'b1111100000011110; // vC=-2018 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111101; // iC= -451 
// vC = 14'b1111100001011000; // vC=-1960 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101011; // iC= -533 
// vC = 14'b1111100011000000; // vC=-1856 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001101001; // iC= -407 
// vC = 14'b1111011110100010; // vC=-2142 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100010; // iC= -414 
// vC = 14'b1111100001011011; // vC=-1957 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111000; // iC= -584 
// vC = 14'b1111100000110101; // vC=-1995 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000011; // iC= -573 
// vC = 14'b1111011111010101; // vC=-2091 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111010000; // iC= -560 
// vC = 14'b1111011110001010; // vC=-2166 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111101; // iC= -451 
// vC = 14'b1111011111011010; // vC=-2086 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001011000; // iC= -424 
// vC = 14'b1111011111101010; // vC=-2070 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111101; // iC= -451 
// vC = 14'b1111100010111100; // vC=-1860 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110011; // iC= -333 
// vC = 14'b1111100001110101; // vC=-1931 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100010; // iC= -478 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010100010; // iC= -350 
// vC = 14'b1111100010001100; // vC=-1908 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010101111; // iC= -337 
// vC = 14'b1111100001101100; // vC=-1940 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010101; // iC= -299 
// vC = 14'b1111100001010101; // vC=-1963 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101010; // iC= -214 
// vC = 14'b1111100001100100; // vC=-1948 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001100110; // iC= -410 
// vC = 14'b1111100010011000; // vC=-1896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101101; // iC= -275 
// vC = 14'b1111100001111010; // vC=-1926 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000111; // iC= -121 
// vC = 14'b1111011111000011; // vC=-2109 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100010; // iC= -222 
// vC = 14'b1111100000100011; // vC=-2013 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100100111; // iC= -217 
// vC = 14'b1111011110000111; // vC=-2169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101010; // iC= -150 
// vC = 14'b1111011110101110; // vC=-2130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101010; // iC= -214 
// vC = 14'b1111100010000110; // vC=-1914 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001101; // iC= -243 
// vC = 14'b1111100000100100; // vC=-2012 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001110; // iC=   14 
// vC = 14'b1111011111101110; // vC=-2066 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110110001; // iC=  -79 
// vC = 14'b1111011110100101; // vC=-2139 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111000; // iC= -200 
// vC = 14'b1111100010001001; // vC=-1911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101101; // iC= -211 
// vC = 14'b1111011111111001; // vC=-2055 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100100; // iC=   36 
// vC = 14'b1111011111011101; // vC=-2083 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100101001; // iC= -215 
// vC = 14'b1111100000110100; // vC=-1996 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110010111; // iC= -105 
// vC = 14'b1111100000011110; // vC=-2018 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000110101; // iC=   53 
// vC = 14'b1111100010111110; // vC=-1858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011101; // iC=   93 
// vC = 14'b1111100000010110; // vC=-2026 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111101; // iC=  -67 
// vC = 14'b1111011110010110; // vC=-2154 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100001; // iC=   97 
// vC = 14'b1111100000101111; // vC=-2001 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101011; // iC=  -21 
// vC = 14'b1111100000100100; // vC=-2012 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101111; // iC=  -17 
// vC = 14'b1111100010110111; // vC=-1865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001000011; // iC=   67 
// vC = 14'b1111011111100001; // vC=-2079 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111110; // iC=  190 
// vC = 14'b1111011110010001; // vC=-2159 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100101; // iC=  165 
// vC = 14'b1111100010011110; // vC=-1890 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111001; // iC=  185 
// vC = 14'b1111011110000010; // vC=-2174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010010; // iC=  338 
// vC = 14'b1111011111001110; // vC=-2098 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111001; // iC=  185 
// vC = 14'b1111100001011000; // vC=-1960 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101101; // iC=  109 
// vC = 14'b1111100010001001; // vC=-1911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100101; // iC=  293 
// vC = 14'b1111100000110100; // vC=-1996 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010101000; // iC=  168 
// vC = 14'b1111100000011000; // vC=-2024 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010100; // iC=  212 
// vC = 14'b1111100000000001; // vC=-2047 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100001100; // iC=  268 
// vC = 14'b1111011110110111; // vC=-2121 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100100; // iC=  420 
// vC = 14'b1111011111101100; // vC=-2068 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101010; // iC=  362 
// vC = 14'b1111011111000110; // vC=-2106 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011101011; // iC=  235 
// vC = 14'b1111011110010100; // vC=-2156 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010001; // iC=  273 
// vC = 14'b1111011110111010; // vC=-2118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100111; // iC=  359 
// vC = 14'b1111100010000111; // vC=-1913 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000101; // iC=  517 
// vC = 14'b1111011110111010; // vC=-2118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010101; // iC=  405 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110010; // iC=  626 
// vC = 14'b1111011111010100; // vC=-2092 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110010; // iC=  498 
// vC = 14'b1111100000101101; // vC=-2003 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010111100; // iC=  700 
// vC = 14'b1111011111101010; // vC=-2070 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110110; // iC=  566 
// vC = 14'b1111100000111000; // vC=-1992 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010111; // iC=  727 
// vC = 14'b1111100010011111; // vC=-1889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100000; // iC=  672 
// vC = 14'b1111011111010100; // vC=-2092 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000100; // iC=  708 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010110111; // iC=  695 
// vC = 14'b1111100000111010; // vC=-1990 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100110; // iC=  806 
// vC = 14'b1111011111111100; // vC=-2052 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111111; // iC=  831 
// vC = 14'b1111011111000111; // vC=-2105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101110; // iC=  750 
// vC = 14'b1111100010010000; // vC=-1904 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011001; // iC=  793 
// vC = 14'b1111100010000000; // vC=-1920 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011100; // iC=  668 
// vC = 14'b1111100010000001; // vC=-1919 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101101; // iC=  941 
// vC = 14'b1111011111111101; // vC=-2051 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011000; // iC=  792 
// vC = 14'b1111011111011101; // vC=-2083 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110010; // iC=  818 
// vC = 14'b1111100000100100; // vC=-2012 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011101; // iC=  861 
// vC = 14'b1111100100000100; // vC=-1788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100111; // iC=  807 
// vC = 14'b1111100001101101; // vC=-1939 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100011; // iC=  931 
// vC = 14'b1111100010110101; // vC=-1867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000010; // iC=  962 
// vC = 14'b1111100011001101; // vC=-1843 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111010; // iC=  826 
// vC = 14'b1111100011110000; // vC=-1808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110110001; // iC=  945 
// vC = 14'b1111100001011011; // vC=-1957 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111010; // iC=  826 
// vC = 14'b1111100011011010; // vC=-1830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000010; // iC=  962 
// vC = 14'b1111100010100101; // vC=-1883 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010111; // iC= 1111 
// vC = 14'b1111100011101111; // vC=-1809 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011010; // iC=  986 
// vC = 14'b1111100010000001; // vC=-1919 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100011; // iC= 1059 
// vC = 14'b1111100000010001; // vC=-2031 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001110; // iC= 1230 
// vC = 14'b1111100001100111; // vC=-1945 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011101; // iC= 1181 
// vC = 14'b1111100000011001; // vC=-2023 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110110; // iC= 1078 
// vC = 14'b1111100000001010; // vC=-2038 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011100; // iC= 1180 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011000; // iC= 1112 
// vC = 14'b1111100001111111; // vC=-1921 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100111; // iC= 1191 
// vC = 14'b1111100001100101; // vC=-1947 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000100; // iC= 1220 
// vC = 14'b1111100000111101; // vC=-1987 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110010; // iC= 1074 
// vC = 14'b1111100100011100; // vC=-1764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001110; // iC= 1166 
// vC = 14'b1111100011000110; // vC=-1850 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011100; // iC= 1244 
// vC = 14'b1111100001000111; // vC=-1977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001000; // iC= 1288 
// vC = 14'b1111100101011101; // vC=-1699 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110110; // iC= 1462 
// vC = 14'b1111100010101110; // vC=-1874 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000010; // iC= 1410 
// vC = 14'b1111100100100010; // vC=-1758 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111101; // iC= 1213 
// vC = 14'b1111100001011000; // vC=-1960 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101101; // iC= 1261 
// vC = 14'b1111100110000100; // vC=-1660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111110; // iC= 1278 
// vC = 14'b1111100010011000; // vC=-1896 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000000; // iC= 1344 
// vC = 14'b1111100010010110; // vC=-1898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011110; // iC= 1246 
// vC = 14'b1111100011101111; // vC=-1809 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101100; // iC= 1516 
// vC = 14'b1111100100100110; // vC=-1754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100100; // iC= 1380 
// vC = 14'b1111100100010000; // vC=-1776 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000010101; // iC= 1557 
// vC = 14'b1111100100000001; // vC=-1791 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001111; // iC= 1423 
// vC = 14'b1111100011000100; // vC=-1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000001; // iC= 1473 
// vC = 14'b1111100100000011; // vC=-1789 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011010; // iC= 1562 
// vC = 14'b1111100100011101; // vC=-1763 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111100; // iC= 1404 
// vC = 14'b1111100110000101; // vC=-1659 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001011; // iC= 1419 
// vC = 14'b1111100101110101; // vC=-1675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011010; // iC= 1498 
// vC = 14'b1111100010101100; // vC=-1876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000110; // iC= 1606 
// vC = 14'b1111100011010000; // vC=-1840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101010; // iC= 1450 
// vC = 14'b1111100010110110; // vC=-1866 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101101; // iC= 1453 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011100; // iC= 1756 
// vC = 14'b1111100100101001; // vC=-1751 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100011; // iC= 1507 
// vC = 14'b1111100101100011; // vC=-1693 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110111; // iC= 1783 
// vC = 14'b1111100100011111; // vC=-1761 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011100; // iC= 1692 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111100; // iC= 1532 
// vC = 14'b1111100100010000; // vC=-1776 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101111; // iC= 1583 
// vC = 14'b1111100101101000; // vC=-1688 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100100; // iC= 1764 
// vC = 14'b1111101000001001; // vC=-1527 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111111; // iC= 1855 
// vC = 14'b1111100110111110; // vC=-1602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110000; // iC= 1776 
// vC = 14'b1111100100110100; // vC=-1740 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011011; // iC= 1755 
// vC = 14'b1111100100010110; // vC=-1770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100111; // iC= 1895 
// vC = 14'b1111100101111011; // vC=-1669 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110010; // iC= 1906 
// vC = 14'b1111100101000001; // vC=-1727 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110110; // iC= 1846 
// vC = 14'b1111100111000001; // vC=-1599 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100010; // iC= 1762 
// vC = 14'b1111100110101001; // vC=-1623 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101101; // iC= 1645 
// vC = 14'b1111101000101011; // vC=-1493 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100001; // iC= 1825 
// vC = 14'b1111101001101000; // vC=-1432 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b1111101000001101; // vC=-1523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010001; // iC= 1873 
// vC = 14'b1111101000001111; // vC=-1521 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000010; // iC= 1858 
// vC = 14'b1111101001100010; // vC=-1438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110000; // iC= 1840 
// vC = 14'b1111100101001001; // vC=-1719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b1111100110010111; // vC=-1641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b1111100110010110; // vC=-1642 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b1111101001111110; // vC=-1410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101111; // iC= 1775 
// vC = 14'b1111100111010111; // vC=-1577 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010011; // iC= 1875 
// vC = 14'b1111101001000011; // vC=-1469 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110111; // iC= 1719 
// vC = 14'b1111100110001111; // vC=-1649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b1111100110110011; // vC=-1613 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b1111100111000000; // vC=-1600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b1111101001111110; // vC=-1410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111010; // iC= 1786 
// vC = 14'b1111101010110111; // vC=-1353 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b1111101001010000; // vC=-1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111100111100100; // vC=-1564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b1111101010011000; // vC=-1384 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110011; // iC= 1779 
// vC = 14'b1111101000011010; // vC=-1510 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000110; // iC= 1798 
// vC = 14'b1111100111101110; // vC=-1554 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000001; // iC= 2049 
// vC = 14'b1111101001111110; // vC=-1410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100010; // iC= 2082 
// vC = 14'b1111101001111111; // vC=-1409 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101111; // iC= 1839 
// vC = 14'b1111101011010001; // vC=-1327 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b1111101010000001; // vC=-1407 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110001; // iC= 1841 
// vC = 14'b1111101011010000; // vC=-1328 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100000; // iC= 1888 
// vC = 14'b1111101011111111; // vC=-1281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b1111101100100101; // vC=-1243 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111101011110001; // vC=-1295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101010; // iC= 1898 
// vC = 14'b1111101001110010; // vC=-1422 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b1111101010010010; // vC=-1390 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011100; // iC= 1820 
// vC = 14'b1111101001100010; // vC=-1438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001100; // iC= 1868 
// vC = 14'b1111101001101010; // vC=-1430 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b1111101101011100; // vC=-1188 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011100; // iC= 2140 
// vC = 14'b1111101001010000; // vC=-1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b1111101011110111; // vC=-1289 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111100; // iC= 1916 
// vC = 14'b1111101001111001; // vC=-1415 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b1111101100100001; // vC=-1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010101; // iC= 2005 
// vC = 14'b1111101010110011; // vC=-1357 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b1111101110000111; // vC=-1145 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001100; // iC= 2060 
// vC = 14'b1111101011101001; // vC=-1303 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b1111101100100001; // vC=-1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000010; // iC= 1922 
// vC = 14'b1111101101011001; // vC=-1191 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001101; // iC= 1997 
// vC = 14'b1111101101100111; // vC=-1177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111001; // iC= 2169 
// vC = 14'b1111101100101001; // vC=-1239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b1111101100100001; // vC=-1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b1111101011001011; // vC=-1333 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b1111101011111010; // vC=-1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111000; // iC= 1912 
// vC = 14'b1111101100110000; // vC=-1232 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010000; // iC= 2192 
// vC = 14'b1111101100000100; // vC=-1276 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111101111010001; // vC=-1071 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011111; // iC= 2015 
// vC = 14'b1111101110110110; // vC=-1098 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111101011101000; // vC=-1304 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110111; // iC= 2167 
// vC = 14'b1111101100101010; // vC=-1238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b1111101100000100; // vC=-1276 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111101111010101; // vC=-1067 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011000; // iC= 2200 
// vC = 14'b1111101111101010; // vC=-1046 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b1111101100100001; // vC=-1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b1111110000010010; // vC=-1006 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b1111110000011010; // vC= -998 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b1111101101111101; // vC=-1155 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101000; // iC= 2152 
// vC = 14'b1111101111011010; // vC=-1062 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111010; // iC= 2106 
// vC = 14'b1111101110011100; // vC=-1124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101011; // iC= 1963 
// vC = 14'b1111110001011011; // vC= -933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010000; // iC= 2192 
// vC = 14'b1111101101101100; // vC=-1172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111110; // iC= 1918 
// vC = 14'b1111101101110110; // vC=-1162 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100000; // iC= 2080 
// vC = 14'b1111110000100100; // vC= -988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b1111110001100100; // vC= -924 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b1111101111000010; // vC=-1086 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000011; // iC= 1923 
// vC = 14'b1111101110111110; // vC=-1090 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000001; // iC= 2177 
// vC = 14'b1111110010110101; // vC= -843 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111110000000010; // vC=-1022 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101110; // iC= 2222 
// vC = 14'b1111110011011001; // vC= -807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011011; // iC= 2075 
// vC = 14'b1111110010111001; // vC= -839 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101110; // iC= 2222 
// vC = 14'b1111110010010101; // vC= -875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001000; // iC= 1992 
// vC = 14'b1111110010100001; // vC= -863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111101111010011; // vC=-1069 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b1111101111111101; // vC=-1027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100110; // iC= 2150 
// vC = 14'b1111110011101000; // vC= -792 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011111; // iC= 2207 
// vC = 14'b1111101111111010; // vC=-1030 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111100; // iC= 2044 
// vC = 14'b1111110001111111; // vC= -897 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011111; // iC= 2143 
// vC = 14'b1111110011101010; // vC= -790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b1111110011111100; // vC= -772 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011000; // iC= 1944 
// vC = 14'b1111110001010101; // vC= -939 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111110101000110; // vC= -698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100100; // iC= 2084 
// vC = 14'b1111110101001101; // vC= -691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b1111110100011110; // vC= -738 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b1111110010111000; // vC= -840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111100; // iC= 2236 
// vC = 14'b1111110001100111; // vC= -921 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001101; // iC= 2061 
// vC = 14'b1111110101000010; // vC= -702 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111110001101101; // vC= -915 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100110; // iC= 2022 
// vC = 14'b1111110001111000; // vC= -904 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b1111110100010100; // vC= -748 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111111; // iC= 2175 
// vC = 14'b1111110101110000; // vC= -656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111011; // iC= 2107 
// vC = 14'b1111110011110000; // vC= -784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111110; // iC= 1982 
// vC = 14'b1111110011010001; // vC= -815 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b1111110110100110; // vC= -602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001011; // iC= 2251 
// vC = 14'b1111110101101000; // vC= -664 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b1111110110110101; // vC= -587 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b1111110101101100; // vC= -660 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101101; // iC= 2221 
// vC = 14'b1111110101111011; // vC= -645 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101101; // iC= 2093 
// vC = 14'b1111110101100111; // vC= -665 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011100; // iC= 2140 
// vC = 14'b1111110110010000; // vC= -624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b1111110110000110; // vC= -634 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b1111110101101111; // vC= -657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011110; // iC= 1950 
// vC = 14'b1111110111101010; // vC= -534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100111; // iC= 2023 
// vC = 14'b1111110011110100; // vC= -780 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111100; // iC= 2108 
// vC = 14'b1111110110111100; // vC= -580 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111111; // iC= 2239 
// vC = 14'b1111110111101110; // vC= -530 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111110; // iC= 2046 
// vC = 14'b1111111000100101; // vC= -475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000100; // iC= 2180 
// vC = 14'b1111111000111000; // vC= -456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101010; // iC= 2090 
// vC = 14'b1111110100110000; // vC= -720 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b1111110100010100; // vC= -748 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010010; // iC= 2002 
// vC = 14'b1111110110110111; // vC= -585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100111; // iC= 2151 
// vC = 14'b1111110111001110; // vC= -562 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001011; // iC= 2123 
// vC = 14'b1111110111100000; // vC= -544 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b1111110111111000; // vC= -520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b1111111001010000; // vC= -432 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b1111111000000010; // vC= -510 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b1111110101100000; // vC= -672 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111011; // iC= 2235 
// vC = 14'b1111111001100110; // vC= -410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110000; // iC= 2032 
// vC = 14'b1111110111100001; // vC= -543 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b1111111001110110; // vC= -394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011011; // iC= 2011 
// vC = 14'b1111110110011001; // vC= -615 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010001; // iC= 2001 
// vC = 14'b1111110111000100; // vC= -572 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010000; // iC= 2256 
// vC = 14'b1111111001001111; // vC= -433 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111111011000010; // vC= -318 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b1111111010100110; // vC= -346 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b1111110111101100; // vC= -532 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010011; // iC= 2195 
// vC = 14'b1111111000000001; // vC= -511 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010101; // iC= 1941 
// vC = 14'b1111110110110001; // vC= -591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100111; // iC= 2023 
// vC = 14'b1111111001000000; // vC= -448 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011110; // iC= 2014 
// vC = 14'b1111110111010000; // vC= -560 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110001; // iC= 2161 
// vC = 14'b1111111010111111; // vC= -321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111101; // iC= 2045 
// vC = 14'b1111111001000100; // vC= -444 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b1111111001000010; // vC= -446 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b1111111000010001; // vC= -495 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100011; // iC= 2147 
// vC = 14'b1111111100101110; // vC= -210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010110; // iC= 2262 
// vC = 14'b1111111100011100; // vC= -228 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b1111111001101111; // vC= -401 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110000; // iC= 2160 
// vC = 14'b1111111100101011; // vC= -213 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010111; // iC= 1943 
// vC = 14'b1111111001100110; // vC= -410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011100; // iC= 2012 
// vC = 14'b1111111001001001; // vC= -439 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101011; // iC= 1963 
// vC = 14'b1111111011001011; // vC= -309 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b1111111101101101; // vC= -147 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010100111; // iC= 2215 
// vC = 14'b1111111101001110; // vC= -178 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b1111111100101110; // vC= -210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100011; // iC= 1955 
// vC = 14'b1111111100110001; // vC= -207 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b1111111011110101; // vC= -267 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b1111111010101010; // vC= -342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100110; // iC= 2022 
// vC = 14'b1111111010101000; // vC= -344 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111100; // iC= 2108 
// vC = 14'b1111111100010110; // vC= -234 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b1111111011001100; // vC= -308 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111111101001100; // vC= -180 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111010; // iC= 2106 
// vC = 14'b1111111011110111; // vC= -265 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010001; // iC= 2193 
// vC = 14'b1111111100101000; // vC= -216 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110110; // iC= 2102 
// vC = 14'b1111111010100101; // vC= -347 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010000; // iC= 2192 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101111; // iC= 1967 
// vC = 14'b1111111110011000; // vC= -104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000110; // iC= 2182 
// vC = 14'b1111111101101110; // vC= -146 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111110; // iC= 1982 
// vC = 14'b1111111111111000; // vC=   -8 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b1111111100010111; // vC= -233 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001000; // iC= 2184 
// vC = 14'b1111111011010001; // vC= -303 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001011; // iC= 1995 
// vC = 14'b1111111110001101; // vC= -115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111111; // iC= 2111 
// vC = 14'b1111111110001110; // vC= -114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010110; // iC= 2006 
// vC = 14'b1111111111100101; // vC=  -27 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101010; // iC= 2218 
// vC = 14'b1111111101010111; // vC= -169 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b1111111100100111; // vC= -217 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110100; // iC= 2228 
// vC = 14'b1111111110111010; // vC=  -70 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111100; // iC= 2172 
// vC = 14'b1111111110000110; // vC= -122 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010101; // iC= 2133 
// vC = 14'b1111111111001100; // vC=  -52 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100110; // iC= 2022 
// vC = 14'b0000000000100010; // vC=   34 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111110; // iC= 2110 
// vC = 14'b1111111100111010; // vC= -198 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111010; // iC= 2170 
// vC = 14'b1111111111011001; // vC=  -39 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b1111111110011110; // vC=  -98 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101011; // iC= 2155 
// vC = 14'b1111111101001011; // vC= -181 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001001; // iC= 2121 
// vC = 14'b0000000000100010; // vC=   34 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b0000000010000011; // vC=  131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000000; // iC= 2176 
// vC = 14'b0000000000100101; // vC=   37 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110011; // iC= 1971 
// vC = 14'b0000000000111011; // vC=   59 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b1111111110111110; // vC=  -66 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b0000000000000010; // vC=    2 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111100; // iC= 1916 
// vC = 14'b0000000001101010; // vC=  106 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010000; // iC= 2128 
// vC = 14'b0000000011000110; // vC=  198 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001010; // iC= 2122 
// vC = 14'b1111111110111010; // vC=  -70 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001010; // iC= 1994 
// vC = 14'b0000000001110101; // vC=  117 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b1111111111000001; // vC=  -63 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111111; // iC= 2175 
// vC = 14'b0000000010000111; // vC=  135 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000101; // iC= 2053 
// vC = 14'b0000000001010110; // vC=   86 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b0000000010010100; // vC=  148 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110101; // iC= 1909 
// vC = 14'b0000000011101100; // vC=  236 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001101; // iC= 2189 
// vC = 14'b0000000100001101; // vC=  269 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100010; // iC= 1890 
// vC = 14'b0000000011101011; // vC=  235 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011111; // iC= 1887 
// vC = 14'b0000000010011111; // vC=  159 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b0000000011000001; // vC=  193 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010000; // iC= 2064 
// vC = 14'b0000000011101110; // vC=  238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110111; // iC= 2103 
// vC = 14'b0000000011100010; // vC=  226 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b0000000000010111; // vC=   23 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101011; // iC= 1899 
// vC = 14'b0000000011010001; // vC=  209 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110000; // iC= 2096 
// vC = 14'b0000000011110010; // vC=  242 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000100; // iC= 1924 
// vC = 14'b0000000001000011; // vC=   67 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110001; // iC= 1905 
// vC = 14'b0000000001101000; // vC=  104 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101000; // iC= 2088 
// vC = 14'b0000000001100000; // vC=   96 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b0000000101000101; // vC=  325 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011101; // iC= 2141 
// vC = 14'b0000000110000101; // vC=  389 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000000; // iC= 1984 
// vC = 14'b0000000101000010; // vC=  322 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b0000000011001011; // vC=  203 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110101; // iC= 2037 
// vC = 14'b0000000100100010; // vC=  290 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010100; // iC= 2068 
// vC = 14'b0000000001101001; // vC=  105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011001; // iC= 2073 
// vC = 14'b0000000101000000; // vC=  320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b0000000110011001; // vC=  409 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101001; // iC= 2153 
// vC = 14'b0000000011010111; // vC=  215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010100; // iC= 2004 
// vC = 14'b0000000110011001; // vC=  409 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b0000000011010110; // vC=  214 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b0000000100000000; // vC=  256 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100111; // iC= 2087 
// vC = 14'b0000000111011011; // vC=  475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111101; // iC= 1981 
// vC = 14'b0000000101000000; // vC=  320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111011; // iC= 1979 
// vC = 14'b0000000100011100; // vC=  284 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b0000000100101000; // vC=  296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100001; // iC= 2017 
// vC = 14'b0000000101100010; // vC=  354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010110; // iC= 2070 
// vC = 14'b0000000111111000; // vC=  504 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b0000000100010110; // vC=  278 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101001; // iC= 1897 
// vC = 14'b0000000110010000; // vC=  400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b0000000101111010; // vC=  378 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b0000000011110011; // vC=  243 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001011; // iC= 1867 
// vC = 14'b0000000111011111; // vC=  479 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b0000000111111101; // vC=  509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b0000000111001001; // vC=  457 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001111; // iC= 1935 
// vC = 14'b0000001000001010; // vC=  522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101000; // iC= 1832 
// vC = 14'b0000000101010011; // vC=  339 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010110; // iC= 2070 
// vC = 14'b0000000111101110; // vC=  494 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110000; // iC= 2096 
// vC = 14'b0000000101010111; // vC=  343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b0000000111110011; // vC=  499 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101101; // iC= 1837 
// vC = 14'b0000001001101000; // vC=  616 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b0000000101101110; // vC=  366 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101010; // iC= 1898 
// vC = 14'b0000000101011101; // vC=  349 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010101; // iC= 1877 
// vC = 14'b0000001010010011; // vC=  659 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100001; // iC= 1825 
// vC = 14'b0000001001111100; // vC=  636 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000010; // iC= 2114 
// vC = 14'b0000001001110100; // vC=  628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010001; // iC= 1937 
// vC = 14'b0000000110001001; // vC=  393 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b0000000110101010; // vC=  426 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100000; // iC= 1824 
// vC = 14'b0000000110100001; // vC=  417 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b0000000111111001; // vC=  505 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000100; // iC= 1796 
// vC = 14'b0000001000111101; // vC=  573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b0000001001110110; // vC=  630 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111101; // iC= 2045 
// vC = 14'b0000001011001101; // vC=  717 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100011; // iC= 1827 
// vC = 14'b0000001000101000; // vC=  552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000000; // iC= 1792 
// vC = 14'b0000000111011000; // vC=  472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b0000001010100010; // vC=  674 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110110; // iC= 1910 
// vC = 14'b0000001011000010; // vC=  706 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111001; // iC= 1849 
// vC = 14'b0000001000001001; // vC=  521 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110011; // iC= 1907 
// vC = 14'b0000001000010101; // vC=  533 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000111; // iC= 1991 
// vC = 14'b0000001010010101; // vC=  661 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011001; // iC= 1881 
// vC = 14'b0000001001011011; // vC=  603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010010; // iC= 1746 
// vC = 14'b0000001100000000; // vC=  768 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b0000001100110100; // vC=  820 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101001; // iC= 2025 
// vC = 14'b0000001011111111; // vC=  767 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011110; // iC= 1822 
// vC = 14'b0000001011001111; // vC=  719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000011; // iC= 1923 
// vC = 14'b0000001000110011; // vC=  563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000110; // iC= 1926 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010111; // iC= 2007 
// vC = 14'b0000001001111010; // vC=  634 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b0000001011101110; // vC=  750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100110; // iC= 1894 
// vC = 14'b0000001100000010; // vC=  770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110011; // iC= 1779 
// vC = 14'b0000001001011010; // vC=  602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010001; // iC= 1873 
// vC = 14'b0000001001010101; // vC=  597 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111001; // iC= 1849 
// vC = 14'b0000001101110011; // vC=  883 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010110; // iC= 1750 
// vC = 14'b0000001100001110; // vC=  782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011001; // iC= 1817 
// vC = 14'b0000001101001101; // vC=  845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100001; // iC= 1697 
// vC = 14'b0000001100111110; // vC=  830 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000001; // iC= 1857 
// vC = 14'b0000001101001000; // vC=  840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001010; // iC= 1866 
// vC = 14'b0000001101111000; // vC=  888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b0000001011110010; // vC=  754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001110; // iC= 1934 
// vC = 14'b0000001011011011; // vC=  731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100001; // iC= 1889 
// vC = 14'b0000001010001101; // vC=  653 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111111; // iC= 1983 
// vC = 14'b0000001111000001; // vC=  961 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b0000001101001011; // vC=  843 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010011; // iC= 1875 
// vC = 14'b0000001100000010; // vC=  770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b0000001110000010; // vC=  898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001000; // iC= 1864 
// vC = 14'b0000001101111010; // vC=  890 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b0000001100000010; // vC=  770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011000; // iC= 1816 
// vC = 14'b0000001110100100; // vC=  932 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001100; // iC= 1676 
// vC = 14'b0000001101101010; // vC=  874 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110001; // iC= 1905 
// vC = 14'b0000001111100001; // vC=  993 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b0000001110010011; // vC=  915 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101110; // iC= 1838 
// vC = 14'b0000001110110011; // vC=  947 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111100; // iC= 1724 
// vC = 14'b0000010000001110; // vC= 1038 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100011; // iC= 1699 
// vC = 14'b0000001100110110; // vC=  822 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111010; // iC= 1786 
// vC = 14'b0000001110110100; // vC=  948 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001100; // iC= 1932 
// vC = 14'b0000001111111100; // vC= 1020 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100111; // iC= 1831 
// vC = 14'b0000010000011010; // vC= 1050 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001011; // iC= 1931 
// vC = 14'b0000001111100010; // vC=  994 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101101; // iC= 1709 
// vC = 14'b0000001110111010; // vC=  954 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010010; // iC= 1618 
// vC = 14'b0000001101011100; // vC=  860 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100011; // iC= 1699 
// vC = 14'b0000001111111001; // vC= 1017 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101100; // iC= 1644 
// vC = 14'b0000001110100101; // vC=  933 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101101000; // iC= 1896 
// vC = 14'b0000001110101111; // vC=  943 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101111; // iC= 1775 
// vC = 14'b0000001110000011; // vC=  899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111001; // iC= 1913 
// vC = 14'b0000001110001111; // vC=  911 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101110; // iC= 1646 
// vC = 14'b0000001101110010; // vC=  882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001110; // iC= 1806 
// vC = 14'b0000001111100110; // vC=  998 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111110; // iC= 1790 
// vC = 14'b0000010001111101; // vC= 1149 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000000; // iC= 1664 
// vC = 14'b0000010001111101; // vC= 1149 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011000; // iC= 1624 
// vC = 14'b0000001111011110; // vC=  990 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100101; // iC= 1765 
// vC = 14'b0000010000011101; // vC= 1053 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111111; // iC= 1855 
// vC = 14'b0000001111010011; // vC=  979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010100; // iC= 1684 
// vC = 14'b0000010000011001; // vC= 1049 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b0000001110100111; // vC=  935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011101110; // iC= 1774 
// vC = 14'b0000010001010100; // vC= 1108 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111011; // iC= 1659 
// vC = 14'b0000010010000110; // vC= 1158 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001001; // iC= 1801 
// vC = 14'b0000001111011010; // vC=  986 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101011; // iC= 1579 
// vC = 14'b0000001111111011; // vC= 1019 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100101; // iC= 1765 
// vC = 14'b0000001111011000; // vC=  984 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001110; // iC= 1550 
// vC = 14'b0000010010010110; // vC= 1174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001111; // iC= 1551 
// vC = 14'b0000010000101000; // vC= 1064 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100001; // iC= 1697 
// vC = 14'b0000010001000111; // vC= 1095 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101100; // iC= 1580 
// vC = 14'b0000010010010100; // vC= 1172 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100010; // iC= 1826 
// vC = 14'b0000010011101101; // vC= 1261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100010; // iC= 1570 
// vC = 14'b0000010001010110; // vC= 1110 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000111; // iC= 1799 
// vC = 14'b0000010010101101; // vC= 1197 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011101; // iC= 1821 
// vC = 14'b0000010100000110; // vC= 1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111011; // iC= 1595 
// vC = 14'b0000010011000110; // vC= 1222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000111; // iC= 1799 
// vC = 14'b0000010100011100; // vC= 1308 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010011; // iC= 1747 
// vC = 14'b0000010000100000; // vC= 1056 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111001; // iC= 1593 
// vC = 14'b0000010001000001; // vC= 1089 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001001; // iC= 1673 
// vC = 14'b0000010100011001; // vC= 1305 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101100; // iC= 1708 
// vC = 14'b0000010011011100; // vC= 1244 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001011; // iC= 1739 
// vC = 14'b0000010010110000; // vC= 1200 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000011; // iC= 1667 
// vC = 14'b0000010011010111; // vC= 1239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011011; // iC= 1499 
// vC = 14'b0000010010101010; // vC= 1194 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001010; // iC= 1610 
// vC = 14'b0000010010110111; // vC= 1207 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011000; // iC= 1560 
// vC = 14'b0000010011111011; // vC= 1275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001111; // iC= 1679 
// vC = 14'b0000010001101011; // vC= 1131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110100; // iC= 1460 
// vC = 14'b0000010100101011; // vC= 1323 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110110111; // iC= 1463 
// vC = 14'b0000010001100000; // vC= 1120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001110; // iC= 1614 
// vC = 14'b0000010101110111; // vC= 1399 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001101; // iC= 1485 
// vC = 14'b0000010100010011; // vC= 1299 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110100; // iC= 1588 
// vC = 14'b0000010001100100; // vC= 1124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010010; // iC= 1490 
// vC = 14'b0000010010000001; // vC= 1153 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100110; // iC= 1510 
// vC = 14'b0000010100001001; // vC= 1289 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100110; // iC= 1510 
// vC = 14'b0000010011010111; // vC= 1239 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101010; // iC= 1578 
// vC = 14'b0000010001101111; // vC= 1135 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011001; // iC= 1497 
// vC = 14'b0000010101101110; // vC= 1390 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011101; // iC= 1501 
// vC = 14'b0000010100001111; // vC= 1295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111011; // iC= 1659 
// vC = 14'b0000010110001111; // vC= 1423 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010110; // iC= 1430 
// vC = 14'b0000010110111010; // vC= 1466 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110010; // iC= 1586 
// vC = 14'b0000010110010011; // vC= 1427 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000111; // iC= 1671 
// vC = 14'b0000010011010101; // vC= 1237 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100000; // iC= 1632 
// vC = 14'b0000010100011111; // vC= 1311 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010100; // iC= 1492 
// vC = 14'b0000010101011000; // vC= 1368 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011110; // iC= 1630 
// vC = 14'b0000010111010001; // vC= 1489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100000; // iC= 1568 
// vC = 14'b0000010111011100; // vC= 1500 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101101; // iC= 1517 
// vC = 14'b0000010111011101; // vC= 1501 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101111; // iC= 1647 
// vC = 14'b0000010110100010; // vC= 1442 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111100; // iC= 1596 
// vC = 14'b0000010111111010; // vC= 1530 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011000; // iC= 1496 
// vC = 14'b0000010101001110; // vC= 1358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101110; // iC= 1454 
// vC = 14'b0000010110010111; // vC= 1431 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111110; // iC= 1342 
// vC = 14'b0000010100000110; // vC= 1286 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101101; // iC= 1517 
// vC = 14'b0000010110000001; // vC= 1409 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110000; // iC= 1328 
// vC = 14'b0000010110111100; // vC= 1468 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011101; // iC= 1309 
// vC = 14'b0000010111001111; // vC= 1487 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100101; // iC= 1509 
// vC = 14'b0000010111100111; // vC= 1511 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001101; // iC= 1421 
// vC = 14'b0000010101101110; // vC= 1390 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100100; // iC= 1508 
// vC = 14'b0000010111011001; // vC= 1497 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101101; // iC= 1517 
// vC = 14'b0000011000100111; // vC= 1575 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101011; // iC= 1387 
// vC = 14'b0000010111011110; // vC= 1502 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111110; // iC= 1342 
// vC = 14'b0000010101011101; // vC= 1373 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111100010; // iC= 1506 
// vC = 14'b0000010101000011; // vC= 1347 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111101; // iC= 1277 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110011; // iC= 1331 
// vC = 14'b0000010101010111; // vC= 1367 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110101; // iC= 1333 
// vC = 14'b0000010110101100; // vC= 1452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010000; // iC= 1424 
// vC = 14'b0000010100111000; // vC= 1336 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110100; // iC= 1268 
// vC = 14'b0000011001010010; // vC= 1618 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010001; // iC= 1489 
// vC = 14'b0000010111001001; // vC= 1481 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110100; // iC= 1268 
// vC = 14'b0000011000100001; // vC= 1569 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111110; // iC= 1278 
// vC = 14'b0000010111011101; // vC= 1501 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110110; // iC= 1334 
// vC = 14'b0000010111001110; // vC= 1486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011011; // iC= 1499 
// vC = 14'b0000010111011100; // vC= 1500 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110100; // iC= 1268 
// vC = 14'b0000010111110011; // vC= 1523 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000101; // iC= 1285 
// vC = 14'b0000010101001111; // vC= 1359 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000100; // iC= 1348 
// vC = 14'b0000010101101101; // vC= 1389 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001010; // iC= 1418 
// vC = 14'b0000010101110011; // vC= 1395 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110000; // iC= 1392 
// vC = 14'b0000010110001110; // vC= 1422 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000011; // iC= 1475 
// vC = 14'b0000011001101000; // vC= 1640 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111010; // iC= 1274 
// vC = 14'b0000010110011110; // vC= 1438 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100000; // iC= 1312 
// vC = 14'b0000011001010101; // vC= 1621 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100011; // iC= 1443 
// vC = 14'b0000011001100000; // vC= 1632 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100101; // iC= 1445 
// vC = 14'b0000011010111010; // vC= 1722 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001000; // iC= 1288 
// vC = 14'b0000010110011100; // vC= 1436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000110; // iC= 1286 
// vC = 14'b0000010110100000; // vC= 1440 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000111; // iC= 1351 
// vC = 14'b0000011001010011; // vC= 1619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100000; // iC= 1440 
// vC = 14'b0000010111110110; // vC= 1526 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100100; // iC= 1380 
// vC = 14'b0000011001100111; // vC= 1639 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010100; // iC= 1364 
// vC = 14'b0000011000100100; // vC= 1572 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111011; // iC= 1147 
// vC = 14'b0000011011000111; // vC= 1735 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010001011; // iC= 1163 
// vC = 14'b0000011000010100; // vC= 1556 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100010; // iC= 1378 
// vC = 14'b0000011010110110; // vC= 1718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100110; // iC= 1254 
// vC = 14'b0000011011101110; // vC= 1774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001101; // iC= 1357 
// vC = 14'b0000011000000101; // vC= 1541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101000110; // iC= 1350 
// vC = 14'b0000011010110001; // vC= 1713 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101110; // iC= 1198 
// vC = 14'b0000010111111011; // vC= 1531 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001010; // iC= 1354 
// vC = 14'b0000011001001100; // vC= 1612 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110110; // iC= 1398 
// vC = 14'b0000011010001100; // vC= 1676 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000011; // iC= 1155 
// vC = 14'b0000011010000110; // vC= 1670 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010101; // iC= 1109 
// vC = 14'b0000010111101001; // vC= 1513 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101110; // iC= 1134 
// vC = 14'b0000010111100101; // vC= 1509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101100; // iC= 1324 
// vC = 14'b0000011000111000; // vC= 1592 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000111; // iC= 1095 
// vC = 14'b0000011010110100; // vC= 1716 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110101; // iC= 1333 
// vC = 14'b0000011011100111; // vC= 1767 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010011; // iC= 1299 
// vC = 14'b0000011000000001; // vC= 1537 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011011; // iC= 1115 
// vC = 14'b0000011000110101; // vC= 1589 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111000; // iC= 1080 
// vC = 14'b0000011001001000; // vC= 1608 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111001; // iC= 1273 
// vC = 14'b0000011000000100; // vC= 1540 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111111; // iC= 1023 
// vC = 14'b0000011001101110; // vC= 1646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010110001; // iC= 1201 
// vC = 14'b0000011010000010; // vC= 1666 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111000; // iC= 1208 
// vC = 14'b0000011100100011; // vC= 1827 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100010; // iC= 1058 
// vC = 14'b0000011100000111; // vC= 1799 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111101; // iC= 1021 
// vC = 14'b0000011000001101; // vC= 1549 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010111; // iC= 1111 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011000; // iC=  984 
// vC = 14'b0000011011010001; // vC= 1745 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001111; // iC= 1295 
// vC = 14'b0000011000100101; // vC= 1573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011000; // iC=  984 
// vC = 14'b0000011001011000; // vC= 1624 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010111001; // iC= 1209 
// vC = 14'b0000011100101001; // vC= 1833 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110110; // iC= 1014 
// vC = 14'b0000011010011010; // vC= 1690 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100000; // iC= 1248 
// vC = 14'b0000011010100100; // vC= 1700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001000; // iC= 1224 
// vC = 14'b0000011100111101; // vC= 1853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011111; // iC= 1119 
// vC = 14'b0000011001111111; // vC= 1663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011001100; // iC= 1228 
// vC = 14'b0000011011000110; // vC= 1734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001101; // iC= 1037 
// vC = 14'b0000011101110101; // vC= 1909 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011110; // iC=  926 
// vC = 14'b0000011010100101; // vC= 1701 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110001; // iC= 1009 
// vC = 14'b0000011100000000; // vC= 1792 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011010; // iC= 1050 
// vC = 14'b0000011101000111; // vC= 1863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000100; // iC= 1028 
// vC = 14'b0000011101000111; // vC= 1863 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000011; // iC= 1091 
// vC = 14'b0000011001100101; // vC= 1637 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011010; // iC= 1114 
// vC = 14'b0000011010001110; // vC= 1678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100101; // iC= 1061 
// vC = 14'b0000011010111010; // vC= 1722 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101010; // iC= 1194 
// vC = 14'b0000011011110110; // vC= 1782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100110; // iC= 1190 
// vC = 14'b0000011101001110; // vC= 1870 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001111100; // iC= 1148 
// vC = 14'b0000011011000110; // vC= 1734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100111; // iC=  935 
// vC = 14'b0000011101111100; // vC= 1916 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001000001; // iC= 1089 
// vC = 14'b0000011011011010; // vC= 1754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110001; // iC=  881 
// vC = 14'b0000011110110000; // vC= 1968 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010001; // iC= 1041 
// vC = 14'b0000011010010111; // vC= 1687 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001010; // iC=  842 
// vC = 14'b0000011110000101; // vC= 1925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010110; // iC=  918 
// vC = 14'b0000011011010000; // vC= 1744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000110; // iC=  966 
// vC = 14'b0000011111001011; // vC= 1995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011011; // iC= 1051 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010111; // iC=  983 
// vC = 14'b0000011101100111; // vC= 1895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100001; // iC=  865 
// vC = 14'b0000011011110001; // vC= 1777 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111110; // iC=  830 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110100; // iC=  820 
// vC = 14'b0000011111010001; // vC= 2001 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101011110; // iC=  862 
// vC = 14'b0000011110111100; // vC= 1980 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001001; // iC=  969 
// vC = 14'b0000011110100100; // vC= 1956 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001111; // iC=  847 
// vC = 14'b0000011100011100; // vC= 1820 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011110; // iC=  990 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101011; // iC= 1003 
// vC = 14'b0000011100100001; // vC= 1825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011101; // iC=  989 
// vC = 14'b0000011111101010; // vC= 2026 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111001110; // iC=  974 
// vC = 14'b0000011100100000; // vC= 1824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011000; // iC=  984 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011001; // iC= 1049 
// vC = 14'b0000011110101011; // vC= 1963 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000100; // iC=  900 
// vC = 14'b0000011011111100; // vC= 1788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111110; // iC=  894 
// vC = 14'b0000011101010100; // vC= 1876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001101; // iC=  909 
// vC = 14'b0000011100101110; // vC= 1838 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110110; // iC=  886 
// vC = 14'b0000011111100101; // vC= 2021 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111000; // iC=  824 
// vC = 14'b0000011101110100; // vC= 1908 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111010; // iC=  890 
// vC = 14'b0000011110000101; // vC= 1925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001010; // iC=  842 
// vC = 14'b0000011100110001; // vC= 1841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010001; // iC=  721 
// vC = 14'b0000011110001110; // vC= 1934 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010100; // iC=  852 
// vC = 14'b0000011011101010; // vC= 1770 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011011; // iC=  667 
// vC = 14'b0000011110100001; // vC= 1953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001010; // iC=  778 
// vC = 14'b0000100000010011; // vC= 2067 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001101; // iC=  909 
// vC = 14'b0000011011110001; // vC= 1777 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100101; // iC=  741 
// vC = 14'b0000011111111010; // vC= 2042 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000100; // iC=  772 
// vC = 14'b0000100000010111; // vC= 2071 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010010001; // iC=  657 
// vC = 14'b0000011110111100; // vC= 1980 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010001; // iC=  785 
// vC = 14'b0000100000000110; // vC= 2054 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011001; // iC=  729 
// vC = 14'b0000011101011011; // vC= 1883 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100111; // iC=  743 
// vC = 14'b0000011110010110; // vC= 1942 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000010; // iC=  706 
// vC = 14'b0000100000010000; // vC= 2064 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100101; // iC=  741 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100110000; // iC=  816 
// vC = 14'b0000100000011011; // vC= 2075 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100110; // iC=  742 
// vC = 14'b0000011100001110; // vC= 1806 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010001; // iC=  593 
// vC = 14'b0000011100001010; // vC= 1802 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010001; // iC=  721 
// vC = 14'b0000011111101011; // vC= 2027 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110111; // iC=  759 
// vC = 14'b0000011100011000; // vC= 1816 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101000; // iC=  680 
// vC = 14'b0000011100010010; // vC= 1810 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100101; // iC=  613 
// vC = 14'b0000011110100011; // vC= 1955 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101000; // iC=  744 
// vC = 14'b0000011111001111; // vC= 1999 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100010; // iC=  546 
// vC = 14'b0000011101100011; // vC= 1891 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001001; // iC=  841 
// vC = 14'b0000100001011011; // vC= 2139 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100100100; // iC=  804 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000101010; // iC=  554 
// vC = 14'b0000100001001010; // vC= 2122 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000011110; // iC=  542 
// vC = 14'b0000011111101111; // vC= 2031 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000000000; // iC=  512 
// vC = 14'b0000011110001111; // vC= 1935 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101100; // iC=  620 
// vC = 14'b0000011100110101; // vC= 1845 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100100; // iC=  740 
// vC = 14'b0000011110100100; // vC= 1956 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111010011; // iC=  467 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100001; // iC=  609 
// vC = 14'b0000011110000111; // vC= 1927 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000001110; // iC=  526 
// vC = 14'b0000011111100011; // vC= 2019 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110100110; // iC=  422 
// vC = 14'b0000011101100001; // vC= 1889 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010100; // iC=  596 
// vC = 14'b0000011101000000; // vC= 1856 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011001; // iC=  409 
// vC = 14'b0000011111010110; // vC= 2006 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100010; // iC=  610 
// vC = 14'b0000100000000110; // vC= 2054 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001001; // iC=  649 
// vC = 14'b0000100000100010; // vC= 2082 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001010110; // iC=  598 
// vC = 14'b0000011110010101; // vC= 1941 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101000; // iC=  424 
// vC = 14'b0000011101110010; // vC= 1906 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100100; // iC=  484 
// vC = 14'b0000100000110011; // vC= 2099 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110001; // iC=  561 
// vC = 14'b0000011110001100; // vC= 1932 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000101; // iC=  581 
// vC = 14'b0000011110001110; // vC= 1934 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111110; // iC=  382 
// vC = 14'b0000100000101000; // vC= 2088 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100000; // iC=  480 
// vC = 14'b0000011101100001; // vC= 1889 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010011; // iC=  531 
// vC = 14'b0000100000111010; // vC= 2106 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000100; // iC=  324 
// vC = 14'b0000011101010100; // vC= 1876 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100010; // iC=  226 
// vC = 14'b0000011110001110; // vC= 1934 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001111; // iC=  207 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110111; // iC=  375 
// vC = 14'b0000100010000000; // vC= 2176 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000101; // iC=  453 
// vC = 14'b0000011101111001; // vC= 1913 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011000110; // iC=  198 
// vC = 14'b0000011101100100; // vC= 1892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011101; // iC=  413 
// vC = 14'b0000011101111110; // vC= 1918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110000; // iC=  240 
// vC = 14'b0000011111000011; // vC= 1987 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111101; // iC=  253 
// vC = 14'b0000011110101101; // vC= 1965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101010001; // iC=  337 
// vC = 14'b0000100000011100; // vC= 2076 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011001; // iC=   89 
// vC = 14'b0000100001011110; // vC= 2142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101111; // iC=  111 
// vC = 14'b0000011110011101; // vC= 1949 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011110010; // iC=  242 
// vC = 14'b0000011110001110; // vC= 1934 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001001001; // iC=   73 
// vC = 14'b0000011101010010; // vC= 1874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010100001; // iC=  161 
// vC = 14'b0000011101110101; // vC= 1909 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011010010; // iC=  210 
// vC = 14'b0000100000000000; // vC= 2048 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010001; // iC=  273 
// vC = 14'b0000100000001110; // vC= 2062 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010010; // iC=  -46 
// vC = 14'b0000100000110111; // vC= 2103 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111110; // iC=  126 
// vC = 14'b0000011111001011; // vC= 1995 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101001; // iC=  105 
// vC = 14'b0000011110001000; // vC= 1928 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110000; // iC=  176 
// vC = 14'b0000011111100000; // vC= 2016 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100100; // iC=   36 
// vC = 14'b0000100001001101; // vC= 2125 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111110110; // iC=  -10 
// vC = 14'b0000011101100110; // vC= 1894 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000001010; // iC=   10 
// vC = 14'b0000011110000110; // vC= 1926 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111100; // iC=  124 
// vC = 14'b0000011111100101; // vC= 2021 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101101110; // iC= -146 
// vC = 14'b0000100001000001; // vC= 2113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111101111; // iC=  -17 
// vC = 14'b0000100000111001; // vC= 2105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110101110; // iC=  -82 
// vC = 14'b0000011111010101; // vC= 2005 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111110; // iC= -194 
// vC = 14'b0000100001101011; // vC= 2155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011111101; // iC= -259 
// vC = 14'b0000100000011100; // vC= 2076 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100111011; // iC= -197 
// vC = 14'b0000100001101001; // vC= 2153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001011; // iC= -309 
// vC = 14'b0000100010000111; // vC= 2183 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000110; // iC= -250 
// vC = 14'b0000011110001011; // vC= 1931 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111100; // iC= -388 
// vC = 14'b0000011110110100; // vC= 1972 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011001011; // iC= -309 
// vC = 14'b0000011101011001; // vC= 1881 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010100; // iC= -364 
// vC = 14'b0000100000110001; // vC= 2097 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011110; // iC= -226 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011101010; // iC= -278 
// vC = 14'b0000011110110011; // vC= 1971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011101; // iC= -227 
// vC = 14'b0000100001010101; // vC= 2133 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110100; // iC= -396 
// vC = 14'b0000100000011111; // vC= 2079 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010100; // iC= -300 
// vC = 14'b0000011101101001; // vC= 1897 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111011; // iC= -581 
// vC = 14'b0000100000111100; // vC= 2108 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100111; // iC= -537 
// vC = 14'b0000011101100111; // vC= 1895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001000111; // iC= -441 
// vC = 14'b0000011101010101; // vC= 1877 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111111011; // iC= -517 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110100100; // iC= -604 
// vC = 14'b0000100001010110; // vC= 2134 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011000; // iC= -616 
// vC = 14'b0000100000101111; // vC= 2095 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010010; // iC= -686 
// vC = 14'b0000100001000110; // vC= 2118 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101011; // iC= -725 
// vC = 14'b0000100000010100; // vC= 2068 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111000000; // iC= -576 
// vC = 14'b0000011110100011; // vC= 1955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111110000; // iC= -528 
// vC = 14'b0000011100110111; // vC= 1847 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001011; // iC= -629 
// vC = 14'b0000011111011111; // vC= 2015 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111011001; // iC= -551 
// vC = 14'b0000011111101000; // vC= 2024 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111001; // iC= -839 
// vC = 14'b0000100000000011; // vC= 2051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001000; // iC= -696 
// vC = 14'b0000011111011100; // vC= 2012 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010010101; // iC= -875 
// vC = 14'b0000011100010111; // vC= 1815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101011; // iC= -917 
// vC = 14'b0000100000010110; // vC= 2070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100011; // iC= -861 
// vC = 14'b0000100000010111; // vC= 2071 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001000; // iC= -696 
// vC = 14'b0000100000111101; // vC= 2109 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011101; // iC= -867 
// vC = 14'b0000011101001001; // vC= 1865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010010; // iC=-1006 
// vC = 14'b0000100000110010; // vC= 2098 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111000; // iC= -904 
// vC = 14'b0000011111000011; // vC= 1987 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001100100; // iC= -924 
// vC = 14'b0000011111010000; // vC= 2000 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011011; // iC= -869 
// vC = 14'b0000011111001001; // vC= 1993 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011010; // iC= -870 
// vC = 14'b0000011101110111; // vC= 1911 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001011; // iC= -821 
// vC = 14'b0000100000001110; // vC= 2062 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010100; // iC=-1004 
// vC = 14'b0000011101100010; // vC= 1890 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000100; // iC=-1084 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111111010; // iC=-1030 
// vC = 14'b0000011011110011; // vC= 1779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011100; // iC=-1060 
// vC = 14'b0000011111010110; // vC= 2006 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011010; // iC=-1062 
// vC = 14'b0000011111101101; // vC= 2029 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000100; // iC=-1084 
// vC = 14'b0000011011111101; // vC= 1789 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111010; // iC=-1094 
// vC = 14'b0000011110011010; // vC= 1946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101101111; // iC=-1169 
// vC = 14'b0000011101111000; // vC= 1912 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010110; // iC=-1130 
// vC = 14'b0000011110010111; // vC= 1943 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000111; // iC=-1273 
// vC = 14'b0000011110110000; // vC= 1968 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001100; // iC=-1332 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110001; // iC=-1167 
// vC = 14'b0000011101010111; // vC= 1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011111; // iC=-1377 
// vC = 14'b0000011011101001; // vC= 1769 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100011; // iC=-1373 
// vC = 14'b0000011010110100; // vC= 1716 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001111; // iC=-1329 
// vC = 14'b0000011111000111; // vC= 1991 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100101; // iC=-1371 
// vC = 14'b0000011101010001; // vC= 1873 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111101; // iC=-1219 
// vC = 14'b0000011110011001; // vC= 1945 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010110; // iC=-1258 
// vC = 14'b0000011011101000; // vC= 1768 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101101; // iC=-1427 
// vC = 14'b0000011101001011; // vC= 1867 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000111; // iC=-1209 
// vC = 14'b0000011010111000; // vC= 1720 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000010; // iC=-1278 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110111; // iC=-1353 
// vC = 14'b0000011110000001; // vC= 1921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101101; // iC=-1363 
// vC = 14'b0000011010011110; // vC= 1694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010000; // iC=-1328 
// vC = 14'b0000011010101111; // vC= 1711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110101; // iC=-1547 
// vC = 14'b0000011110010101; // vC= 1941 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010111; // iC=-1513 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111111; // iC=-1345 
// vC = 14'b0000011001101001; // vC= 1641 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101111; // iC=-1361 
// vC = 14'b0000011101100111; // vC= 1895 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101001; // iC=-1623 
// vC = 14'b0000011001001010; // vC= 1610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000110; // iC=-1658 
// vC = 14'b0000011100011111; // vC= 1823 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001101; // iC=-1459 
// vC = 14'b0000011010011011; // vC= 1691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011100; // iC=-1444 
// vC = 14'b0000011011101011; // vC= 1771 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101010; // iC=-1430 
// vC = 14'b0000011011101111; // vC= 1775 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111111; // iC=-1473 
// vC = 14'b0000011010000110; // vC= 1670 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110101; // iC=-1675 
// vC = 14'b0000011011111001; // vC= 1785 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100001; // iC=-1759 
// vC = 14'b0000011011111010; // vC= 1786 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010011; // iC=-1517 
// vC = 14'b0000011001110010; // vC= 1650 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000001; // iC=-1663 
// vC = 14'b0000011100111011; // vC= 1851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101111; // iC=-1617 
// vC = 14'b0000011100000111; // vC= 1799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010101; // iC=-1515 
// vC = 14'b0000011010001010; // vC= 1674 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111110; // iC=-1794 
// vC = 14'b0000011010111001; // vC= 1721 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010100; // iC=-1644 
// vC = 14'b0000011010110001; // vC= 1713 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010111; // iC=-1641 
// vC = 14'b0000011001001101; // vC= 1613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011111; // iC=-1633 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111110; // iC=-1602 
// vC = 14'b0000011011101010; // vC= 1770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111010; // iC=-1670 
// vC = 14'b0000011011111101; // vC= 1789 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001111; // iC=-1841 
// vC = 14'b0000011000010110; // vC= 1558 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000101; // iC=-1851 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010011; // iC=-1709 
// vC = 14'b0000011000110000; // vC= 1584 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011011; // iC=-1701 
// vC = 14'b0000010110101011; // vC= 1451 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000111; // iC=-1721 
// vC = 14'b0000011010011111; // vC= 1695 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001111; // iC=-1649 
// vC = 14'b0000011001110110; // vC= 1654 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101010; // iC=-1814 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011000; // iC=-1896 
// vC = 14'b0000010111010010; // vC= 1490 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111100; // iC=-1988 
// vC = 14'b0000010110111000; // vC= 1464 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101111; // iC=-1937 
// vC = 14'b0000010111110001; // vC= 1521 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b0000010111101010; // vC= 1514 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b0000010111100101; // vC= 1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001001; // iC=-1847 
// vC = 14'b0000010101011110; // vC= 1374 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100101; // iC=-1755 
// vC = 14'b0000010110101011; // vC= 1451 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b0000011000011111; // vC= 1567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100101; // iC=-1883 
// vC = 14'b0000010110110100; // vC= 1460 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b0000010101110011; // vC= 1395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000101; // iC=-1787 
// vC = 14'b0000011001011010; // vC= 1626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b0000011000010101; // vC= 1557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010110; // iC=-1834 
// vC = 14'b0000010111100101; // vC= 1509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011110; // iC=-2082 
// vC = 14'b0000011001001110; // vC= 1614 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b0000010100101101; // vC= 1325 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000011000000101; // vC= 1541 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b0000010101000111; // vC= 1351 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000010; // iC=-2046 
// vC = 14'b0000010111101110; // vC= 1518 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b0000010110101010; // vC= 1450 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011011; // iC=-1829 
// vC = 14'b0000010101001111; // vC= 1359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b0000010111000110; // vC= 1478 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000011; // iC=-1981 
// vC = 14'b0000010100110111; // vC= 1335 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000101; // iC=-1851 
// vC = 14'b0000010011011110; // vC= 1246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000001; // iC=-1855 
// vC = 14'b0000010011110000; // vC= 1264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b0000010101001111; // vC= 1359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011101; // iC=-2147 
// vC = 14'b0000010110100001; // vC= 1441 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000010101110010; // vC= 1394 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010100; // iC=-1836 
// vC = 14'b0000010110011010; // vC= 1434 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010110; // iC=-2154 
// vC = 14'b0000010010111001; // vC= 1209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000011; // iC=-1981 
// vC = 14'b0000010110111100; // vC= 1468 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000100; // iC=-2044 
// vC = 14'b0000010010110000; // vC= 1200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b0000010100011100; // vC= 1308 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b0000010100100011; // vC= 1315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000010110011000; // vC= 1432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b0000010001111010; // vC= 1146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101110; // iC=-2130 
// vC = 14'b0000010101001001; // vC= 1353 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100000; // iC=-2016 
// vC = 14'b0000010001011101; // vC= 1117 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b0000010001010111; // vC= 1111 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010011; // iC=-2093 
// vC = 14'b0000010001001000; // vC= 1096 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111101; // iC=-2179 
// vC = 14'b0000010001001111; // vC= 1103 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b0000010011001001; // vC= 1225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011110; // iC=-2146 
// vC = 14'b0000010001010110; // vC= 1110 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111101; // iC=-1923 
// vC = 14'b0000010100010100; // vC= 1300 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b0000010100100100; // vC= 1316 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101001; // iC=-2135 
// vC = 14'b0000010000101010; // vC= 1066 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011110; // iC=-2146 
// vC = 14'b0000010000001101; // vC= 1037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b0000010010010010; // vC= 1170 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110111; // iC=-2121 
// vC = 14'b0000010100001010; // vC= 1290 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110000; // iC=-2064 
// vC = 14'b0000010000011001; // vC= 1049 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110011; // iC=-1997 
// vC = 14'b0000010000101001; // vC= 1065 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111001; // iC=-2183 
// vC = 14'b0000010010101101; // vC= 1197 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110111; // iC=-2121 
// vC = 14'b0000001111001001; // vC=  969 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000010; // iC=-2046 
// vC = 14'b0000010011100111; // vC= 1255 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100011; // iC=-2141 
// vC = 14'b0000010011001101; // vC= 1229 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000101; // iC=-2107 
// vC = 14'b0000010010001110; // vC= 1166 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b0000010000000111; // vC= 1031 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000010000100110; // vC= 1062 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000001; // iC=-1983 
// vC = 14'b0000010000011111; // vC= 1055 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001100; // iC=-1908 
// vC = 14'b0000001110011001; // vC=  921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100000; // iC=-1952 
// vC = 14'b0000010010110110; // vC= 1206 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000010; // iC=-2046 
// vC = 14'b0000010000100111; // vC= 1063 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111100; // iC=-1988 
// vC = 14'b0000010001000011; // vC= 1091 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b0000010001011110; // vC= 1118 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b0000001111110010; // vC= 1010 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b0000001111001111; // vC=  975 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b0000010000001110; // vC= 1038 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100111; // iC=-1945 
// vC = 14'b0000001110011110; // vC=  926 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100100; // iC=-2204 
// vC = 14'b0000001111001001; // vC=  969 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100110; // iC=-2074 
// vC = 14'b0000010000000000; // vC= 1024 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101111; // iC=-2129 
// vC = 14'b0000001101110111; // vC=  887 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b0000001101110010; // vC=  882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b0000010000011011; // vC= 1051 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110000; // iC=-2128 
// vC = 14'b0000001110000100; // vC=  900 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000001100001100; // vC=  780 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010000; // iC=-2032 
// vC = 14'b0000010000100110; // vC= 1062 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100111; // iC=-2073 
// vC = 14'b0000010000101010; // vC= 1066 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b0000001101111110; // vC=  894 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100011; // iC=-2205 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100010; // iC=-2206 
// vC = 14'b0000001011101001; // vC=  745 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000111; // iC=-2233 
// vC = 14'b0000001100001000; // vC=  776 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000010; // iC=-2110 
// vC = 14'b0000001100111011; // vC=  827 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100111; // iC=-2201 
// vC = 14'b0000001100110001; // vC=  817 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b0000001100100111; // vC=  807 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b0000001110010110; // vC=  918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000101; // iC=-2235 
// vC = 14'b0000001011100010; // vC=  738 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b0000001110111010; // vC=  954 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000001; // iC=-2047 
// vC = 14'b0000001100100001; // vC=  801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000100; // iC=-2172 
// vC = 14'b0000001100011101; // vC=  797 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000001101110100; // vC=  884 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111010; // iC=-2246 
// vC = 14'b0000001100100001; // vC=  801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110101; // iC=-2251 
// vC = 14'b0000001001111010; // vC=  634 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011100; // iC=-2212 
// vC = 14'b0000001011100011; // vC=  739 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010010; // iC=-2158 
// vC = 14'b0000001110001110; // vC=  910 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b0000001100111101; // vC=  829 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000001011011100; // vC=  732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101000; // iC=-2136 
// vC = 14'b0000001100001101; // vC=  781 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101001; // iC=-2199 
// vC = 14'b0000001011001000; // vC=  712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b0000001000101011; // vC=  555 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b0000001000010111; // vC=  535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011101; // iC=-2083 
// vC = 14'b0000001010001101; // vC=  653 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b0000001000110111; // vC=  567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110000; // iC=-2192 
// vC = 14'b0000001000110111; // vC=  567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100100100; // iC=-2268 
// vC = 14'b0000001001101000; // vC=  616 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100011; // iC=-2205 
// vC = 14'b0000001000010000; // vC=  528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101111; // iC=-2257 
// vC = 14'b0000001011001001; // vC=  713 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000101; // iC=-2235 
// vC = 14'b0000001011011111; // vC=  735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010001; // iC=-2095 
// vC = 14'b0000001001011111; // vC=  607 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b0000000110111101; // vC=  445 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b0000001000010000; // vC=  528 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110001; // iC=-2127 
// vC = 14'b0000001011101001; // vC=  745 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100111; // iC=-2137 
// vC = 14'b0000001010110111; // vC=  695 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101111; // iC=-2257 
// vC = 14'b0000000110101111; // vC=  431 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100001; // iC=-2079 
// vC = 14'b0000000111001000; // vC=  456 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010101; // iC=-2219 
// vC = 14'b0000001001100011; // vC=  611 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b0000000101111101; // vC=  381 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110100; // iC=-2124 
// vC = 14'b0000000110001001; // vC=  393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b0000001001100010; // vC=  610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001100; // iC=-2228 
// vC = 14'b0000001001110010; // vC=  626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011011; // iC=-2021 
// vC = 14'b0000000110011001; // vC=  409 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b0000001001011001; // vC=  601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110100; // iC=-2188 
// vC = 14'b0000000110001001; // vC=  393 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b0000000111101100; // vC=  492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b0000000111000011; // vC=  451 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b0000000110100001; // vC=  417 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100001; // iC=-2207 
// vC = 14'b0000000111100111; // vC=  487 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110011; // iC=-2125 
// vC = 14'b0000000101110011; // vC=  371 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100010; // iC=-2142 
// vC = 14'b0000001000111110; // vC=  574 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001111; // iC=-2097 
// vC = 14'b0000000111111101; // vC=  509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110110; // iC=-2250 
// vC = 14'b0000001000001110; // vC=  526 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100011; // iC=-2077 
// vC = 14'b0000000111111000; // vC=  504 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000010; // iC=-2174 
// vC = 14'b0000000100001100; // vC=  268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b0000000101100101; // vC=  357 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011000; // iC=-2216 
// vC = 14'b0000000111101010; // vC=  490 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101101; // iC=-2195 
// vC = 14'b0000001000000000; // vC=  512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000000101101001; // vC=  361 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000000100010100; // vC=  276 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110010; // iC=-1998 
// vC = 14'b0000000110110010; // vC=  434 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100010; // iC=-2078 
// vC = 14'b0000000011110000; // vC=  240 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111110; // iC=-2178 
// vC = 14'b0000000100001000; // vC=  264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110111; // iC=-1993 
// vC = 14'b0000000100010111; // vC=  279 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001100; // iC=-2164 
// vC = 14'b0000000100011010; // vC=  282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110110; // iC=-1994 
// vC = 14'b0000000101000110; // vC=  326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110000; // iC=-2192 
// vC = 14'b0000000010110010; // vC=  178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011001; // iC=-1959 
// vC = 14'b0000000010011101; // vC=  157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101110; // iC=-2066 
// vC = 14'b0000000100001101; // vC=  269 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b0000000011101100; // vC=  236 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000000101110010; // vC=  370 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110110; // iC=-2122 
// vC = 14'b0000000100110101; // vC=  309 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000000; // iC=-2176 
// vC = 14'b0000000101011110; // vC=  350 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001111; // iC=-2161 
// vC = 14'b0000000001010001; // vC=   81 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b0000000100111010; // vC=  314 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011101; // iC=-2083 
// vC = 14'b0000000100100010; // vC=  290 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010001; // iC=-2159 
// vC = 14'b0000000011100010; // vC=  226 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011110; // iC=-1954 
// vC = 14'b0000000010011010; // vC=  154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011001; // iC=-2215 
// vC = 14'b0000000011111001; // vC=  249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001001; // iC=-2231 
// vC = 14'b0000000000011111; // vC=   31 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b0000000001000111; // vC=   71 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000000001010110; // vC=   86 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b1111111111110000; // vC=  -16 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110111; // iC=-2121 
// vC = 14'b0000000000101101; // vC=   45 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110111; // iC=-2185 
// vC = 14'b0000000010101111; // vC=  175 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b0000000000111001; // vC=   57 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011001; // iC=-2151 
// vC = 14'b0000000100000111; // vC=  263 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010101; // iC=-2027 
// vC = 14'b0000000011010010; // vC=  210 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000101; // iC=-2171 
// vC = 14'b0000000010111110; // vC=  190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011010; // iC=-2214 
// vC = 14'b0000000001000011; // vC=   67 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000000001000001; // vC=   65 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110000; // iC=-2064 
// vC = 14'b0000000000100000; // vC=   32 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000010; // iC=-2046 
// vC = 14'b0000000001001000; // vC=   72 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001010; // iC=-2038 
// vC = 14'b0000000011001110; // vC=  206 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001100; // iC=-2228 
// vC = 14'b0000000010100010; // vC=  162 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111011; // iC=-1989 
// vC = 14'b1111111110110010; // vC=  -78 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100101; // iC=-2203 
// vC = 14'b0000000001100100; // vC=  100 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011111; // iC=-2081 
// vC = 14'b1111111110111010; // vC=  -70 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011011; // iC=-2149 
// vC = 14'b0000000001100000; // vC=   96 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100100; // iC=-2204 
// vC = 14'b1111111110011111; // vC=  -97 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010111; // iC=-1961 
// vC = 14'b1111111111000000; // vC=  -64 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010001; // iC=-2159 
// vC = 14'b1111111101110100; // vC= -140 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b1111111100111111; // vC= -193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010100; // iC=-2028 
// vC = 14'b1111111111011110; // vC=  -34 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110110; // iC=-1930 
// vC = 14'b0000000000010100; // vC=   20 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100101; // iC=-2139 
// vC = 14'b1111111110010010; // vC= -110 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100100; // iC=-2140 
// vC = 14'b1111111111010000; // vC=  -48 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101000; // iC=-2200 
// vC = 14'b0000000000110101; // vC=   53 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000110; // iC=-1978 
// vC = 14'b1111111110111111; // vC=  -65 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101101; // iC=-2195 
// vC = 14'b0000000000111001; // vC=   57 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111101; // iC=-1923 
// vC = 14'b1111111101001010; // vC= -182 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b1111111111111011; // vC=   -5 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b1111111011100001; // vC= -287 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111000; // iC=-2120 
// vC = 14'b1111111100111010; // vC= -198 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011110; // iC=-2018 
// vC = 14'b1111111111001011; // vC=  -53 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110000; // iC=-2128 
// vC = 14'b1111111101000010; // vC= -190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011101; // iC=-2147 
// vC = 14'b1111111100111111; // vC= -193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111000; // iC=-2184 
// vC = 14'b1111111101110100; // vC= -140 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001000; // iC=-2040 
// vC = 14'b1111111101010101; // vC= -171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b1111111101011000; // vC= -168 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b1111111010111111; // vC= -321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100111; // iC=-2073 
// vC = 14'b1111111101100101; // vC= -155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011000; // iC=-2088 
// vC = 14'b1111111011100000; // vC= -288 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b1111111011011110; // vC= -290 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010010; // iC=-2158 
// vC = 14'b1111111100111110; // vC= -194 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110001; // iC=-2063 
// vC = 14'b1111111100000010; // vC= -254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b1111111110011000; // vC= -104 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000110; // iC=-2170 
// vC = 14'b1111111100001101; // vC= -243 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b1111111010111010; // vC= -326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000101; // iC=-1979 
// vC = 14'b1111111100110100; // vC= -204 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001100; // iC=-2036 
// vC = 14'b1111111011110100; // vC= -268 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b1111111100101110; // vC= -210 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b1111111101001101; // vC= -179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010101; // iC=-2091 
// vC = 14'b1111111100010101; // vC= -235 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111111; // iC=-2113 
// vC = 14'b1111111000111111; // vC= -449 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111110; // iC=-1922 
// vC = 14'b1111111100100011; // vC= -221 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101010; // iC=-2006 
// vC = 14'b1111111001101100; // vC= -404 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111101; // iC=-1923 
// vC = 14'b1111111001010000; // vC= -432 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110000; // iC=-2128 
// vC = 14'b1111111011010000; // vC= -304 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b1111111000110101; // vC= -459 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000010; // iC=-1918 
// vC = 14'b1111111000010111; // vC= -489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b1111111010001111; // vC= -369 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100011; // iC=-2141 
// vC = 14'b1111111011101010; // vC= -278 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111000; // iC=-1928 
// vC = 14'b1111111010000100; // vC= -380 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101110; // iC=-2130 
// vC = 14'b1111111100000010; // vC= -254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010001; // iC=-1839 
// vC = 14'b1111111000000110; // vC= -506 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110101; // iC=-2123 
// vC = 14'b1111111010010000; // vC= -368 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100101; // iC=-2011 
// vC = 14'b1111111010101011; // vC= -341 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011001; // iC=-2023 
// vC = 14'b1111110111010010; // vC= -558 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001110; // iC=-2098 
// vC = 14'b1111111010111111; // vC= -321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001110; // iC=-1906 
// vC = 14'b1111111010011000; // vC= -360 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b1111111010001001; // vC= -375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b1111110110100110; // vC= -602 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101110; // iC=-1874 
// vC = 14'b1111110110111111; // vC= -577 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111100; // iC=-1796 
// vC = 14'b1111110110110001; // vC= -591 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b1111110111011010; // vC= -550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b1111111001111100; // vC= -388 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b1111111000000000; // vC= -512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b1111110101101001; // vC= -663 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b1111111001001010; // vC= -438 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b1111110101011011; // vC= -677 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b1111111000101110; // vC= -466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b1111110110010001; // vC= -623 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b1111110110110000; // vC= -592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000111; // iC=-1913 
// vC = 14'b1111111000100111; // vC= -473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b1111110110001111; // vC= -625 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000001; // iC=-1983 
// vC = 14'b1111111000010011; // vC= -493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111110; // iC=-1858 
// vC = 14'b1111110101001011; // vC= -693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b1111110101111001; // vC= -647 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110011; // iC=-1805 
// vC = 14'b1111110100011101; // vC= -739 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110010; // iC=-1998 
// vC = 14'b1111110111101011; // vC= -533 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b1111110110000000; // vC= -640 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111000; // iC=-1800 
// vC = 14'b1111110111110001; // vC= -527 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110110; // iC=-1994 
// vC = 14'b1111110101010011; // vC= -685 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b1111110101010101; // vC= -683 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b1111110111111000; // vC= -520 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101101; // iC=-2003 
// vC = 14'b1111110100001011; // vC= -757 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011000; // iC=-1768 
// vC = 14'b1111110100000110; // vC= -762 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110101; // iC=-1867 
// vC = 14'b1111110010111101; // vC= -835 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000011; // iC=-1789 
// vC = 14'b1111110110100111; // vC= -601 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101000; // iC=-1880 
// vC = 14'b1111110011111101; // vC= -771 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000100; // iC=-1852 
// vC = 14'b1111110011000111; // vC= -825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b1111110100011001; // vC= -743 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b1111110100110110; // vC= -714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b1111110100011010; // vC= -742 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010101; // iC=-1771 
// vC = 14'b1111110110110101; // vC= -587 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b1111110110011110; // vC= -610 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011010; // iC=-1958 
// vC = 14'b1111110010111101; // vC= -835 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000100; // iC=-1724 
// vC = 14'b1111110101101111; // vC= -657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010011; // iC=-1901 
// vC = 14'b1111110101111011; // vC= -645 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000001; // iC=-1727 
// vC = 14'b1111110001010110; // vC= -938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b1111110001011010; // vC= -934 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b1111110101010111; // vC= -681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001001; // iC=-1719 
// vC = 14'b1111110010011100; // vC= -868 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000111; // iC=-1849 
// vC = 14'b1111110011110101; // vC= -779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011010; // iC=-1702 
// vC = 14'b1111110000111000; // vC= -968 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b1111110001110011; // vC= -909 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001001; // iC=-1719 
// vC = 14'b1111110001011110; // vC= -930 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b1111110001001000; // vC= -952 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000000; // iC=-1664 
// vC = 14'b1111110010100011; // vC= -861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b1111110001110011; // vC= -909 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b1111110001011000; // vC= -936 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111001; // iC=-1799 
// vC = 14'b1111110100000000; // vC= -768 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001100; // iC=-1844 
// vC = 14'b1111110001101011; // vC= -917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010100; // iC=-1644 
// vC = 14'b1111110001100111; // vC= -921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001101; // iC=-1779 
// vC = 14'b1111110000101000; // vC= -984 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010100; // iC=-1644 
// vC = 14'b1111110100001010; // vC= -758 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011001; // iC=-1831 
// vC = 14'b1111110010001001; // vC= -887 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000100; // iC=-1660 
// vC = 14'b1111110011011010; // vC= -806 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b1111110001101100; // vC= -916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010100; // iC=-1644 
// vC = 14'b1111110000110010; // vC= -974 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111001; // iC=-1607 
// vC = 14'b1111101111110011; // vC=-1037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100001; // iC=-1759 
// vC = 14'b1111110011010100; // vC= -812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110100; // iC=-1676 
// vC = 14'b1111101111100001; // vC=-1055 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001000; // iC=-1848 
// vC = 14'b1111101111001101; // vC=-1075 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010101; // iC=-1643 
// vC = 14'b1111101111110101; // vC=-1035 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011010; // iC=-1702 
// vC = 14'b1111110010101000; // vC= -856 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110101; // iC=-1867 
// vC = 14'b1111110010111101; // vC= -835 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110000; // iC=-1680 
// vC = 14'b1111101110001000; // vC=-1144 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110101; // iC=-1611 
// vC = 14'b1111110010101011; // vC= -853 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101001; // iC=-1879 
// vC = 14'b1111110010010110; // vC= -874 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110111; // iC=-1737 
// vC = 14'b1111101101110101; // vC=-1163 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011111; // iC=-1569 
// vC = 14'b1111101110010100; // vC=-1132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110100; // iC=-1804 
// vC = 14'b1111101111101000; // vC=-1048 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011001; // iC=-1831 
// vC = 14'b1111110000010111; // vC=-1001 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011000; // iC=-1832 
// vC = 14'b1111110010000010; // vC= -894 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101011; // iC=-1557 
// vC = 14'b1111101101100111; // vC=-1177 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001011; // iC=-1717 
// vC = 14'b1111110000001000; // vC=-1016 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110001; // iC=-1807 
// vC = 14'b1111101101111111; // vC=-1153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011010; // iC=-1702 
// vC = 14'b1111110000011110; // vC= -994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001111; // iC=-1649 
// vC = 14'b1111110001010110; // vC= -938 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111100; // iC=-1796 
// vC = 14'b1111110000001001; // vC=-1015 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111110; // iC=-1602 
// vC = 14'b1111101101110001; // vC=-1167 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111001; // iC=-1671 
// vC = 14'b1111101110010100; // vC=-1132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111011; // iC=-1605 
// vC = 14'b1111101101110011; // vC=-1165 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000101; // iC=-1659 
// vC = 14'b1111101100010000; // vC=-1264 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001011; // iC=-1525 
// vC = 14'b1111101100110111; // vC=-1225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001010; // iC=-1654 
// vC = 14'b1111101101111110; // vC=-1154 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110110; // iC=-1802 
// vC = 14'b1111101111101000; // vC=-1048 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000110; // iC=-1658 
// vC = 14'b1111110000100111; // vC= -985 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011100; // iC=-1572 
// vC = 14'b1111101101100101; // vC=-1179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100110; // iC=-1690 
// vC = 14'b1111101110100000; // vC=-1120 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011101; // iC=-1699 
// vC = 14'b1111101100101010; // vC=-1238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100110; // iC=-1562 
// vC = 14'b1111101100001111; // vC=-1265 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001110; // iC=-1650 
// vC = 14'b1111101101011011; // vC=-1189 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100011; // iC=-1501 
// vC = 14'b1111101110011101; // vC=-1123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101010; // iC=-1750 
// vC = 14'b1111101101000010; // vC=-1214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b1111101101000001; // vC=-1215 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011100; // iC=-1700 
// vC = 14'b1111101111110111; // vC=-1033 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001111; // iC=-1585 
// vC = 14'b1111101101000010; // vC=-1214 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010100; // iC=-1452 
// vC = 14'b1111101111100011; // vC=-1053 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011111; // iC=-1633 
// vC = 14'b1111101110111011; // vC=-1093 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100001; // iC=-1631 
// vC = 14'b1111101101011101; // vC=-1187 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101011; // iC=-1685 
// vC = 14'b1111101111000011; // vC=-1085 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000010010; // iC=-1518 
// vC = 14'b1111101100100000; // vC=-1248 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101111; // iC=-1489 
// vC = 14'b1111101011101001; // vC=-1303 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111110011; // iC=-1549 
// vC = 14'b1111101110100011; // vC=-1117 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111011; // iC=-1413 
// vC = 14'b1111101011111000; // vC=-1288 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101101; // iC=-1491 
// vC = 14'b1111101100111000; // vC=-1224 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000110; // iC=-1402 
// vC = 14'b1111101101010101; // vC=-1195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100111; // iC=-1561 
// vC = 14'b1111101100100001; // vC=-1247 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110000; // iC=-1680 
// vC = 14'b1111101010111111; // vC=-1345 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001010; // iC=-1398 
// vC = 14'b1111101011100100; // vC=-1308 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000111; // iC=-1529 
// vC = 14'b1111101010100100; // vC=-1372 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100111; // iC=-1433 
// vC = 14'b1111101101010100; // vC=-1196 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011010; // iC=-1382 
// vC = 14'b1111101010011001; // vC=-1383 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010011; // iC=-1389 
// vC = 14'b1111101100000100; // vC=-1276 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001010; // iC=-1654 
// vC = 14'b1111101010011111; // vC=-1377 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111100; // iC=-1540 
// vC = 14'b1111101001010100; // vC=-1452 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101011; // iC=-1429 
// vC = 14'b1111101010101100; // vC=-1364 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000101; // iC=-1595 
// vC = 14'b1111101100010010; // vC=-1262 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010100; // iC=-1644 
// vC = 14'b1111101010111000; // vC=-1352 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111000; // iC=-1608 
// vC = 14'b1111101011110101; // vC=-1291 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111000000; // iC=-1600 
// vC = 14'b1111101000100101; // vC=-1499 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011011; // iC=-1445 
// vC = 14'b1111101011101110; // vC=-1298 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000000; // iC=-1472 
// vC = 14'b1111101001101011; // vC=-1429 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000001; // iC=-1343 
// vC = 14'b1111101100110111; // vC=-1225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100111; // iC=-1561 
// vC = 14'b1111101000101101; // vC=-1491 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000000000; // iC=-1536 
// vC = 14'b1111101010001011; // vC=-1397 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000001011; // iC=-1525 
// vC = 14'b1111101010110100; // vC=-1356 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011001; // iC=-1383 
// vC = 14'b1111100111100101; // vC=-1563 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011011; // iC=-1509 
// vC = 14'b1111101010010011; // vC=-1389 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001110; // iC=-1394 
// vC = 14'b1111101001001001; // vC=-1463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011001; // iC=-1511 
// vC = 14'b1111101011000010; // vC=-1342 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110111; // iC=-1417 
// vC = 14'b1111100111111000; // vC=-1544 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111011111; // iC=-1569 
// vC = 14'b1111101000100110; // vC=-1498 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101011; // iC=-1557 
// vC = 14'b1111100111100001; // vC=-1567 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111100; // iC=-1284 
// vC = 14'b1111101011000000; // vC=-1344 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101010; // iC=-1430 
// vC = 14'b1111100111111110; // vC=-1538 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011110; // iC=-1314 
// vC = 14'b1111101001001111; // vC=-1457 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101011; // iC=-1557 
// vC = 14'b1111101001100011; // vC=-1437 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100111; // iC=-1497 
// vC = 14'b1111100111001110; // vC=-1586 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011101; // iC=-1443 
// vC = 14'b1111101000011001; // vC=-1511 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011001; // iC=-1319 
// vC = 14'b1111101011010100; // vC=-1324 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000010; // iC=-1406 
// vC = 14'b1111101010111010; // vC=-1350 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000000; // iC=-1472 
// vC = 14'b1111101000101010; // vC=-1494 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101101; // iC=-1235 
// vC = 14'b1111100111110001; // vC=-1551 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011110; // iC=-1378 
// vC = 14'b1111101001000011; // vC=-1469 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111001; // iC=-1479 
// vC = 14'b1111100110000010; // vC=-1662 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010010; // iC=-1198 
// vC = 14'b1111100111101011; // vC=-1557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100101; // iC=-1435 
// vC = 14'b1111100111100110; // vC=-1562 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100001010; // iC=-1270 
// vC = 14'b1111101000100001; // vC=-1503 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011001; // iC=-1447 
// vC = 14'b1111101001011010; // vC=-1446 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111110; // iC=-1282 
// vC = 14'b1111100111100000; // vC=-1568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100100; // iC=-1436 
// vC = 14'b1111100111001011; // vC=-1589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010001; // iC=-1455 
// vC = 14'b1111100110100110; // vC=-1626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011101; // iC=-1379 
// vC = 14'b1111101001001110; // vC=-1458 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110100; // iC=-1356 
// vC = 14'b1111100110010010; // vC=-1646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111111; // iC=-1409 
// vC = 14'b1111101000011111; // vC=-1505 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010011010; // iC=-1382 
// vC = 14'b1111101001100000; // vC=-1440 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100111110; // iC=-1218 
// vC = 14'b1111100110000111; // vC=-1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110010; // iC=-1422 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110010; // iC=-1166 
// vC = 14'b1111100110100010; // vC=-1630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100001; // iC=-1311 
// vC = 14'b1111100100111010; // vC=-1734 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110101; // iC=-1291 
// vC = 14'b1111101000110010; // vC=-1486 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111101; // iC=-1283 
// vC = 14'b1111101001100101; // vC=-1435 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110110; // iC=-1098 
// vC = 14'b1111101000010011; // vC=-1517 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010010; // iC=-1262 
// vC = 14'b1111100110001101; // vC=-1651 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101000001; // iC=-1215 
// vC = 14'b1111100101101000; // vC=-1688 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110101; // iC=-1099 
// vC = 14'b1111100101100010; // vC=-1694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110100; // iC=-1228 
// vC = 14'b1111100100110000; // vC=-1744 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001010; // iC=-1206 
// vC = 14'b1111101000101100; // vC=-1492 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100101; // iC=-1307 
// vC = 14'b1111101000111101; // vC=-1475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011101001; // iC=-1303 
// vC = 14'b1111100101111111; // vC=-1665 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010110; // iC=-1130 
// vC = 14'b1111100111010010; // vC=-1582 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011010; // iC=-1318 
// vC = 14'b1111100101010001; // vC=-1711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110000; // iC=-1296 
// vC = 14'b1111101000010100; // vC=-1516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110110; // iC=-1226 
// vC = 14'b1111100100010100; // vC=-1772 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110101010; // iC=-1110 
// vC = 14'b1111100110111100; // vC=-1604 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111000; // iC=-1096 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000000111; // iC=-1017 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001100; // iC=-1076 
// vC = 14'b1111100111010111; // vC=-1577 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110000; // iC=-1232 
// vC = 14'b1111100011100111; // vC=-1817 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011110; // iC=-1314 
// vC = 14'b1111100100110100; // vC=-1740 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001011; // iC=-1077 
// vC = 14'b1111100101001111; // vC=-1713 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001100; // iC=-1076 
// vC = 14'b1111100100010111; // vC=-1769 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001110; // iC=-1074 
// vC = 14'b1111100110010110; // vC=-1642 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011100; // iC=-1188 
// vC = 14'b1111100101010111; // vC=-1705 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110001011; // iC=-1141 
// vC = 14'b1111100101001011; // vC=-1717 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011110; // iC=-1186 
// vC = 14'b1111100110000111; // vC=-1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101001; // iC= -983 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010011; // iC=-1197 
// vC = 14'b1111100101101010; // vC=-1686 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011001; // iC=-1191 
// vC = 14'b1111100110001100; // vC=-1652 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111011100; // iC=-1060 
// vC = 14'b1111100110110111; // vC=-1609 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000000; // iC=-1088 
// vC = 14'b1111100111000000; // vC=-1600 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110101; // iC=-1099 
// vC = 14'b1111100101100111; // vC=-1689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001010; // iC=-1206 
// vC = 14'b1111100101111000; // vC=-1672 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000001001; // iC=-1015 
// vC = 14'b1111100100111000; // vC=-1736 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110100; // iC=-1036 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100000; // iC= -992 
// vC = 14'b1111100011011111; // vC=-1825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000101011; // iC= -981 
// vC = 14'b1111100010011100; // vC=-1892 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111101000; // iC=-1048 
// vC = 14'b1111100101111010; // vC=-1670 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010111; // iC=-1001 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000000; // iC= -960 
// vC = 14'b1111100100001000; // vC=-1784 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000110011; // iC= -973 
// vC = 14'b1111100100001101; // vC=-1779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111000; // iC= -904 
// vC = 14'b1111100001101010; // vC=-1942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100100; // iC=-1180 
// vC = 14'b1111100010111110; // vC=-1858 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100100; // iC=-1116 
// vC = 14'b1111100011000111; // vC=-1849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010001; // iC=-1071 
// vC = 14'b1111100010010001; // vC=-1903 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000011010; // iC= -998 
// vC = 14'b1111100100101111; // vC=-1745 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111110110; // iC=-1034 
// vC = 14'b1111100110000100; // vC=-1660 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111000; // iC= -904 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100111; // iC= -985 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111111; // iC= -961 
// vC = 14'b1111100011101000; // vC=-1816 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010010; // iC=-1006 
// vC = 14'b1111100011000011; // vC=-1853 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110101; // iC= -843 
// vC = 14'b1111100001010010; // vC=-1966 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100101; // iC= -987 
// vC = 14'b1111100010101001; // vC=-1879 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111001101; // iC=-1075 
// vC = 14'b1111100101010010; // vC=-1710 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110110110; // iC=-1098 
// vC = 14'b1111100100101101; // vC=-1747 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100100; // iC= -860 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010110; // iC=-1002 
// vC = 14'b1111100010101101; // vC=-1875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001110101; // iC= -907 
// vC = 14'b1111100100111001; // vC=-1735 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111101; // iC= -963 
// vC = 14'b1111100101010100; // vC=-1708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010101; // iC= -939 
// vC = 14'b1111100101101100; // vC=-1684 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111010111; // iC=-1065 
// vC = 14'b1111100100101111; // vC=-1745 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111100; // iC= -836 
// vC = 14'b1111100001100000; // vC=-1952 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100000; // iC= -736 
// vC = 14'b1111100010011011; // vC=-1893 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011111010; // iC= -774 
// vC = 14'b1111100101011001; // vC=-1703 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010011; // iC= -749 
// vC = 14'b1111100001010101; // vC=-1963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010110; // iC= -746 
// vC = 14'b1111100100100111; // vC=-1753 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000100001; // iC= -991 
// vC = 14'b1111100001010110; // vC=-1962 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010001100; // iC= -884 
// vC = 14'b1111100001111100; // vC=-1924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111100; // iC= -964 
// vC = 14'b1111100011000001; // vC=-1855 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000111100; // iC= -964 
// vC = 14'b1111100001100001; // vC=-1951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111111; // iC= -833 
// vC = 14'b1111100001111101; // vC=-1923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001111100; // iC= -900 
// vC = 14'b1111100100011001; // vC=-1767 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001101110; // iC= -914 
// vC = 14'b1111100011010101; // vC=-1835 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101011; // iC= -661 
// vC = 14'b1111100011111111; // vC=-1793 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101000; // iC= -792 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101101110; // iC= -658 
// vC = 14'b1111100001101111; // vC=-1937 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101010100; // iC= -684 
// vC = 14'b1111100011011010; // vC=-1830 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011011; // iC= -869 
// vC = 14'b1111100001000010; // vC=-1982 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001011; // iC= -629 
// vC = 14'b1111100000110011; // vC=-1997 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011001110; // iC= -818 
// vC = 14'b1111100000000000; // vC=-2048 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011110101; // iC= -779 
// vC = 14'b1111100100000011; // vC=-1789 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011000001; // iC= -831 
// vC = 14'b1111100001001111; // vC=-1969 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101001; // iC= -855 
// vC = 14'b1111100000101001; // vC=-2007 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100101000; // iC= -728 
// vC = 14'b1111100001100110; // vC=-1946 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010000010; // iC= -894 
// vC = 14'b1111100001010110; // vC=-1962 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111001; // iC= -647 
// vC = 14'b1111100000101010; // vC=-2006 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100110000; // iC= -720 
// vC = 14'b1111011111111011; // vC=-2053 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100010; // iC= -734 
// vC = 14'b1111100000110100; // vC=-1996 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011010; // iC= -678 
// vC = 14'b1111100010111111; // vC=-1857 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100011011; // iC= -741 
// vC = 14'b1111100001100101; // vC=-1947 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011010100; // iC= -812 
// vC = 14'b1111100001100111; // vC=-1945 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111010; // iC= -838 
// vC = 14'b1111100001001001; // vC=-1975 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011100; // iC= -804 
// vC = 14'b1111011111001111; // vC=-2097 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011111; // iC= -609 
// vC = 14'b1111100010011110; // vC=-1890 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101111101; // iC= -643 
// vC = 14'b1111100011101000; // vC=-1816 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100001101; // iC= -755 
// vC = 14'b1111100001100100; // vC=-1948 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100101; // iC= -795 
// vC = 14'b1111011111100011; // vC=-2077 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101101; // iC= -595 
// vC = 14'b1111100011000011; // vC=-1853 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100010111; // iC= -745 
// vC = 14'b1111100001011101; // vC=-1955 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011111; // iC= -481 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111001; // iC= -455 
// vC = 14'b1111100000001110; // vC=-2034 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110011; // iC= -589 
// vC = 14'b1111100001100001; // vC=-1951 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101110001; // iC= -655 
// vC = 14'b1111100011101110; // vC=-1810 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001001001; // iC= -439 
// vC = 14'b1111100010001011; // vC=-1909 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111001000; // iC= -568 
// vC = 14'b1111011111011110; // vC=-2082 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110110011; // iC= -589 
// vC = 14'b1111011111111000; // vC=-2056 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101011111; // iC= -673 
// vC = 14'b1111100001110001; // vC=-1935 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111101100; // iC= -532 
// vC = 14'b1111100011100010; // vC=-1822 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010001100; // iC= -372 
// vC = 14'b1111100010110010; // vC=-1870 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000101101; // iC= -467 
// vC = 14'b1111100001101011; // vC=-1941 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000010001; // iC= -495 
// vC = 14'b1111100001110000; // vC=-1936 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000000000; // iC= -512 
// vC = 14'b1111011110011000; // vC=-2152 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110101001; // iC= -599 
// vC = 14'b1111100001111001; // vC=-1927 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000100010; // iC= -478 
// vC = 14'b1111100000101000; // vC=-2008 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000001; // iC= -383 
// vC = 14'b1111100010001010; // vC=-1910 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100000101; // iC= -251 
// vC = 14'b1111100001001111; // vC=-1969 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000011001; // iC= -487 
// vC = 14'b1111100000011100; // vC=-2020 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010110111; // iC= -329 
// vC = 14'b1111011111011110; // vC=-2082 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010001; // iC= -239 
// vC = 14'b1111011111010011; // vC=-2093 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001010000; // iC= -432 
// vC = 14'b1111100001000110; // vC=-1978 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010111111; // iC= -321 
// vC = 14'b1111100000001111; // vC=-2033 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001101; // iC= -179 
// vC = 14'b1111100010010010; // vC=-1902 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111101; // iC= -387 
// vC = 14'b1111100000100111; // vC=-2009 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101111100; // iC= -132 
// vC = 14'b1111100000101011; // vC=-2005 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010000; // iC= -304 
// vC = 14'b1111100010010101; // vC=-1899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010000101; // iC= -379 
// vC = 14'b1111100000000101; // vC=-2043 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110011110; // iC=  -98 
// vC = 14'b1111100011000110; // vC=-1850 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001000; // iC= -248 
// vC = 14'b1111100010101110; // vC=-1874 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100000; // iC= -160 
// vC = 14'b1111100001101001; // vC=-1943 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110111111; // iC=  -65 
// vC = 14'b1111100011000001; // vC=-1855 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101001110; // iC= -178 
// vC = 14'b1111100000110110; // vC=-1994 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111011101; // iC=  -35 
// vC = 14'b1111100000000000; // vC=-2048 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111100100; // iC=  -28 
// vC = 14'b1111100000111110; // vC=-1986 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100011110; // iC= -226 
// vC = 14'b1111100000110000; // vC=-2000 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111010100; // iC=  -44 
// vC = 14'b1111100000110000; // vC=-2000 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111001001; // iC=  -55 
// vC = 14'b1111011110110010; // vC=-2126 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010110; // iC=   22 
// vC = 14'b1111011110010001; // vC=-2159 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101100001; // iC= -159 
// vC = 14'b1111100011000000; // vC=-1856 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000100; // iC= -124 
// vC = 14'b1111011111100111; // vC=-2073 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101110110; // iC= -138 
// vC = 14'b1111100000101011; // vC=-2005 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001111001; // iC=  121 
// vC = 14'b1111100001001100; // vC=-1972 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110001; // iC=  177 
// vC = 14'b1111100010000101; // vC=-1915 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001110010; // iC=  114 
// vC = 14'b1111011110101100; // vC=-2132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110111; // iC=  183 
// vC = 14'b1111011110011010; // vC=-2150 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101000; // iC=  104 
// vC = 14'b1111011111010100; // vC=-2092 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010000101; // iC=  133 
// vC = 14'b1111100000101010; // vC=-2006 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010001010; // iC=  138 
// vC = 14'b1111011110110100; // vC=-2124 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111110; // iC=  190 
// vC = 14'b1111100000011001; // vC=-2023 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000110; // iC=  326 
// vC = 14'b1111100000000101; // vC=-2043 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011101; // iC=  157 
// vC = 14'b1111100010110111; // vC=-1865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010111110; // iC=  190 
// vC = 14'b1111011111011001; // vC=-2087 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100100111; // iC=  295 
// vC = 14'b1111011111000111; // vC=-2105 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111000010; // iC=  450 
// vC = 14'b1111100000000011; // vC=-2045 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100111100; // iC=  316 
// vC = 14'b1111100001010100; // vC=-1964 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101001; // iC=  425 
// vC = 14'b1111100011001000; // vC=-1848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110000100; // iC=  388 
// vC = 14'b1111011110101100; // vC=-2132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111001110; // iC=  462 
// vC = 14'b1111100000100001; // vC=-2015 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101111100; // iC=  380 
// vC = 14'b1111100001000011; // vC=-1981 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111101; // iC=  445 
// vC = 14'b1111100001110110; // vC=-1930 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110111; // iC=  631 
// vC = 14'b1111100010101101; // vC=-1875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110111; // iC=  503 
// vC = 14'b1111100011011110; // vC=-1826 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110111110; // iC=  446 
// vC = 14'b1111100011001111; // vC=-1841 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110011111; // iC=  415 
// vC = 14'b1111011111100100; // vC=-2076 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100110; // iC=  550 
// vC = 14'b1111100010100110; // vC=-1882 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111100101; // iC=  485 
// vC = 14'b1111100000111100; // vC=-1988 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100100; // iC=  740 
// vC = 14'b1111100001010011; // vC=-1965 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101111; // iC=  687 
// vC = 14'b1111100010000100; // vC=-1916 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110010; // iC=  626 
// vC = 14'b1111100000011000; // vC=-2024 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100110; // iC=  614 
// vC = 14'b1111100001001010; // vC=-1974 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100000; // iC=  608 
// vC = 14'b1111100010010100; // vC=-1900 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010001; // iC=  785 
// vC = 14'b1111100000010001; // vC=-2031 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001111; // iC=  911 
// vC = 14'b1111011111111100; // vC=-2052 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100111; // iC=  615 
// vC = 14'b1111100010101011; // vC=-1877 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011010100; // iC=  724 
// vC = 14'b1111100000111000; // vC=-1992 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010111; // iC=  855 
// vC = 14'b1111100010101010; // vC=-1878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010011; // iC=  851 
// vC = 14'b1111100011111110; // vC=-1794 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101010100; // iC=  852 
// vC = 14'b1111011111011100; // vC=-2084 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101110; // iC=  942 
// vC = 14'b1111100011010111; // vC=-1833 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101111111; // iC=  895 
// vC = 14'b1111100011000101; // vC=-1851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101000011; // iC=  835 
// vC = 14'b1111100010101111; // vC=-1873 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110010; // iC=  882 
// vC = 14'b1111100000110111; // vC=-1993 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000110001; // iC= 1073 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100101; // iC= 1125 
// vC = 14'b1111100001011111; // vC=-1953 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100111; // iC=  871 
// vC = 14'b1111100001111011; // vC=-1925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110010100; // iC=  916 
// vC = 14'b1111100011001011; // vC=-1845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001001; // iC= 1097 
// vC = 14'b1111100001000111; // vC=-1977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110100; // iC= 1012 
// vC = 14'b1111100100010010; // vC=-1774 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101101; // iC=  941 
// vC = 14'b1111100000011111; // vC=-2017 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000100111; // iC= 1063 
// vC = 14'b1111100011110111; // vC=-1801 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011111000; // iC= 1272 
// vC = 14'b1111100000111110; // vC=-1986 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001010; // iC= 1034 
// vC = 14'b1111100001100101; // vC=-1947 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100000; // iC= 1120 
// vC = 14'b1111100001000111; // vC=-1977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101010; // iC= 1194 
// vC = 14'b1111100011110100; // vC=-1804 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011011110; // iC= 1246 
// vC = 14'b1111100001011010; // vC=-1958 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010001; // iC= 1361 
// vC = 14'b1111100011000101; // vC=-1851 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110100; // iC= 1396 
// vC = 14'b1111100101100000; // vC=-1696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000110; // iC= 1286 
// vC = 14'b1111100011000111; // vC=-1849 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110001; // iC= 1393 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110010000; // iC= 1424 
// vC = 14'b1111100100100110; // vC=-1754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111101; // iC= 1469 
// vC = 14'b1111100100001010; // vC=-1782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111001; // iC= 1465 
// vC = 14'b1111100100100101; // vC=-1755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011010; // iC= 1306 
// vC = 14'b1111100110001000; // vC=-1656 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011010; // iC= 1498 
// vC = 14'b1111100100011011; // vC=-1765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010110; // iC= 1366 
// vC = 14'b1111100010001110; // vC=-1906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101100; // iC= 1260 
// vC = 14'b1111100010101010; // vC=-1878 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100010000; // iC= 1296 
// vC = 14'b1111100010001110; // vC=-1906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110000; // iC= 1328 
// vC = 14'b1111100011000010; // vC=-1854 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000111; // iC= 1607 
// vC = 14'b1111100011111100; // vC=-1796 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000100; // iC= 1476 
// vC = 14'b1111100110110111; // vC=-1609 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001000; // iC= 1352 
// vC = 14'b1111100100110001; // vC=-1743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011100; // iC= 1500 
// vC = 14'b1111100111001111; // vC=-1585 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101010; // iC= 1514 
// vC = 14'b1111100100000010; // vC=-1790 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000110101; // iC= 1589 
// vC = 14'b1111100110010111; // vC=-1641 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001101011; // iC= 1643 
// vC = 14'b1111100110111101; // vC=-1603 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101001; // iC= 1449 
// vC = 14'b1111100100010101; // vC=-1771 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010010; // iC= 1682 
// vC = 14'b1111100111011010; // vC=-1574 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011011; // iC= 1435 
// vC = 14'b1111100011001100; // vC=-1844 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111101111; // iC= 1519 
// vC = 14'b1111100101100100; // vC=-1692 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111011000; // iC= 1496 
// vC = 14'b1111100110100111; // vC=-1625 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010100; // iC= 1492 
// vC = 14'b1111100111010100; // vC=-1580 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000001; // iC= 1537 
// vC = 14'b1111101000011101; // vC=-1507 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011001; // iC= 1561 
// vC = 14'b1111100100101010; // vC=-1750 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010111; // iC= 1751 
// vC = 14'b1111100011110001; // vC=-1807 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010111110; // iC= 1726 
// vC = 14'b1111101000000001; // vC=-1535 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b1111100110011101; // vC=-1635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100001; // iC= 1761 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011110; // iC= 1694 
// vC = 14'b1111100101100101; // vC=-1691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010010011; // iC= 1683 
// vC = 14'b1111100101001110; // vC=-1714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110110; // iC= 1654 
// vC = 14'b1111101001000010; // vC=-1470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010101; // iC= 1621 
// vC = 14'b1111101000011101; // vC=-1507 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110010; // iC= 1714 
// vC = 14'b1111101001000011; // vC=-1469 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011000111; // iC= 1735 
// vC = 14'b1111100101001110; // vC=-1714 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110100; // iC= 1780 
// vC = 14'b1111101001001000; // vC=-1464 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001001; // iC= 1801 
// vC = 14'b1111101010000010; // vC=-1406 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111110; // iC= 1662 
// vC = 14'b1111100101011110; // vC=-1698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110100; // iC= 1844 
// vC = 14'b1111101000011000; // vC=-1512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b1111100101111001; // vC=-1671 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100001101; // iC= 1805 
// vC = 14'b1111100110010001; // vC=-1647 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001010; // iC= 1930 
// vC = 14'b1111100111010000; // vC=-1584 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100100; // iC= 1956 
// vC = 14'b1111101000110100; // vC=-1484 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010110; // iC= 1878 
// vC = 14'b1111101000011110; // vC=-1506 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000010; // iC= 1922 
// vC = 14'b1111100111001101; // vC=-1587 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111010; // iC= 2042 
// vC = 14'b1111101001111010; // vC=-1414 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000101; // iC= 1797 
// vC = 14'b1111101001100000; // vC=-1440 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111000; // iC= 1784 
// vC = 14'b1111101010000000; // vC=-1408 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011110; // iC= 1886 
// vC = 14'b1111101011100011; // vC=-1309 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111100; // iC= 1916 
// vC = 14'b1111100110110000; // vC=-1616 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b1111100111100110; // vC=-1562 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b1111101010001110; // vC=-1394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010010; // iC= 2066 
// vC = 14'b1111101001111101; // vC=-1411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010001; // iC= 2065 
// vC = 14'b1111101001100001; // vC=-1439 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010010; // iC= 1938 
// vC = 14'b1111101000010000; // vC=-1520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000100; // iC= 2052 
// vC = 14'b1111101100000100; // vC=-1276 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b1111101000000101; // vC=-1531 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101010; // iC= 1962 
// vC = 14'b1111101001010001; // vC=-1455 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011100; // iC= 2076 
// vC = 14'b1111101001001101; // vC=-1459 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010010; // iC= 2002 
// vC = 14'b1111101000001110; // vC=-1522 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100100; // iC= 1892 
// vC = 14'b1111101011100101; // vC=-1307 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b1111101001010011; // vC=-1453 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000000; // iC= 1984 
// vC = 14'b1111101011110001; // vC=-1295 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100000; // iC= 2080 
// vC = 14'b1111101101000001; // vC=-1215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b1111101011100100; // vC=-1308 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011111; // iC= 2079 
// vC = 14'b1111101010000001; // vC=-1407 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b1111101010010011; // vC=-1389 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011110; // iC= 2142 
// vC = 14'b1111101001010101; // vC=-1451 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101101; // iC= 2093 
// vC = 14'b1111101010010000; // vC=-1392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100011; // iC= 1891 
// vC = 14'b1111101101101000; // vC=-1176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001000; // iC= 1864 
// vC = 14'b1111101010110011; // vC=-1357 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101101; // iC= 2093 
// vC = 14'b1111101110101000; // vC=-1112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010010; // iC= 2066 
// vC = 14'b1111101011011100; // vC=-1316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010100; // iC= 2132 
// vC = 14'b1111101011111111; // vC=-1281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101011; // iC= 1963 
// vC = 14'b1111101101001100; // vC=-1204 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b1111101010101010; // vC=-1366 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b1111101100100001; // vC=-1247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b1111101011111001; // vC=-1287 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001111; // iC= 1871 
// vC = 14'b1111101010110010; // vC=-1358 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101001; // iC= 2153 
// vC = 14'b1111101100001000; // vC=-1272 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b1111101111111010; // vC=-1030 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111101011000010; // vC=-1342 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001010; // iC= 2186 
// vC = 14'b1111101110001000; // vC=-1144 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011010; // iC= 2074 
// vC = 14'b1111101100010010; // vC=-1262 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b1111101101110101; // vC=-1163 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111101101111110; // vC=-1154 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001011; // iC= 2187 
// vC = 14'b1111101100000001; // vC=-1279 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010001; // iC= 1937 
// vC = 14'b1111101111100100; // vC=-1052 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000111; // iC= 1927 
// vC = 14'b1111101111101101; // vC=-1043 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111110; // iC= 1918 
// vC = 14'b1111101110001010; // vC=-1142 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011100; // iC= 1884 
// vC = 14'b1111101110011101; // vC=-1123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100110; // iC= 1958 
// vC = 14'b1111110000100010; // vC= -990 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111101110010010; // vC=-1134 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001010; // iC= 2186 
// vC = 14'b1111101110100010; // vC=-1118 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010010; // iC= 2066 
// vC = 14'b1111101111001000; // vC=-1080 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b1111110000011101; // vC= -995 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110101; // iC= 1973 
// vC = 14'b1111101110101010; // vC=-1110 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001100; // iC= 1996 
// vC = 14'b1111101110110001; // vC=-1103 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110110; // iC= 2038 
// vC = 14'b1111101110010111; // vC=-1129 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001101; // iC= 2189 
// vC = 14'b1111110010010011; // vC= -877 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b1111110000011100; // vC= -996 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001110010; // iC= 2162 
// vC = 14'b1111110010010100; // vC= -876 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000000; // iC= 2048 
// vC = 14'b1111101110001001; // vC=-1143 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110010; // iC= 2034 
// vC = 14'b1111101111011101; // vC=-1059 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111010; // iC= 2170 
// vC = 14'b1111101111011110; // vC=-1058 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000110; // iC= 2182 
// vC = 14'b1111110011011111; // vC= -801 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010000; // iC= 2064 
// vC = 14'b1111110001101101; // vC= -915 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110011; // iC= 2227 
// vC = 14'b1111110011101001; // vC= -791 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111000; // iC= 2168 
// vC = 14'b1111110000101111; // vC= -977 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b1111110010001010; // vC= -886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111110011011110; // vC= -802 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111000; // iC= 2104 
// vC = 14'b1111110100011000; // vC= -744 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000110; // iC= 2054 
// vC = 14'b1111101111111101; // vC=-1027 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000100; // iC= 1988 
// vC = 14'b1111110100000001; // vC= -767 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001111; // iC= 2063 
// vC = 14'b1111110100010110; // vC= -746 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000011; // iC= 1987 
// vC = 14'b1111110011101100; // vC= -788 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001101; // iC= 1933 
// vC = 14'b1111110000100101; // vC= -987 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110111; // iC= 2039 
// vC = 14'b1111110001111111; // vC= -897 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111110; // iC= 2110 
// vC = 14'b1111110100100010; // vC= -734 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001000; // iC= 2056 
// vC = 14'b1111110010000111; // vC= -889 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001000; // iC= 2120 
// vC = 14'b1111110101010110; // vC= -682 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b1111110100101101; // vC= -723 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000110; // iC= 2118 
// vC = 14'b1111110010111000; // vC= -840 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000101; // iC= 2053 
// vC = 14'b1111110010010000; // vC= -880 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001111; // iC= 2127 
// vC = 14'b1111110101010001; // vC= -687 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001010; // iC= 2186 
// vC = 14'b1111110011111001; // vC= -775 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b1111110100011111; // vC= -737 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000000; // iC= 1984 
// vC = 14'b1111110011000111; // vC= -825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b1111110110010101; // vC= -619 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010110; // iC= 2070 
// vC = 14'b1111110011011010; // vC= -806 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110110; // iC= 2102 
// vC = 14'b1111110010001010; // vC= -886 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000101; // iC= 1989 
// vC = 14'b1111110010010011; // vC= -877 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000101; // iC= 2117 
// vC = 14'b1111110110011100; // vC= -612 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101110; // iC= 2158 
// vC = 14'b1111110010101011; // vC= -853 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111101; // iC= 2109 
// vC = 14'b1111110101011101; // vC= -675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111001; // iC= 2041 
// vC = 14'b1111110101101001; // vC= -663 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000000; // iC= 2112 
// vC = 14'b1111110110010010; // vC= -622 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001111; // iC= 2127 
// vC = 14'b1111110101101110; // vC= -658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001110; // iC= 2062 
// vC = 14'b1111110011101111; // vC= -785 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b1111110101110001; // vC= -655 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010101; // iC= 2005 
// vC = 14'b1111110111010010; // vC= -558 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011011; // iC= 1947 
// vC = 14'b1111110100111010; // vC= -710 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101011; // iC= 2091 
// vC = 14'b1111110111110000; // vC= -528 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101001; // iC= 2217 
// vC = 14'b1111110101011010; // vC= -678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110011; // iC= 2035 
// vC = 14'b1111110111101010; // vC= -534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010011; // iC= 2259 
// vC = 14'b1111110110001111; // vC= -625 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010111; // iC= 2071 
// vC = 14'b1111110101110010; // vC= -654 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010101; // iC= 2197 
// vC = 14'b1111110111010000; // vC= -560 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000110; // iC= 2182 
// vC = 14'b1111110110001000; // vC= -632 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111111; // iC= 2175 
// vC = 14'b1111110111010111; // vC= -553 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011010001; // iC= 2257 
// vC = 14'b1111110110011111; // vC= -609 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011110; // iC= 2142 
// vC = 14'b1111111000111111; // vC= -449 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000001; // iC= 2177 
// vC = 14'b1111110111010001; // vC= -559 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000101100; // iC= 2092 
// vC = 14'b1111110111000011; // vC= -573 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110111; // iC= 2039 
// vC = 14'b1111110111100110; // vC= -538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111001; // iC= 2169 
// vC = 14'b1111111010010110; // vC= -362 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001101; // iC= 2125 
// vC = 14'b1111111000000000; // vC= -512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010111; // iC= 2135 
// vC = 14'b1111110111101101; // vC= -531 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001011; // iC= 2059 
// vC = 14'b1111111001110000; // vC= -400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101011; // iC= 2155 
// vC = 14'b1111110110110001; // vC= -591 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010110100; // iC= 2228 
// vC = 14'b1111111011000100; // vC= -316 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100000; // iC= 2080 
// vC = 14'b1111110110100011; // vC= -605 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001111; // iC= 2191 
// vC = 14'b1111111000100101; // vC= -475 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110111; // iC= 1975 
// vC = 14'b1111111000000001; // vC= -511 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111111; // iC= 2239 
// vC = 14'b1111111001101101; // vC= -403 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b1111111000111110; // vC= -450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000001111; // iC= 2063 
// vC = 14'b1111111011100011; // vC= -285 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111111; // iC= 2047 
// vC = 14'b1111111010011110; // vC= -354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100101; // iC= 2021 
// vC = 14'b1111111011010000; // vC= -304 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100011001001; // iC= 2249 
// vC = 14'b1111111011101010; // vC= -278 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111011; // iC= 2171 
// vC = 14'b1111111010100101; // vC= -347 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010011; // iC= 1939 
// vC = 14'b1111111100101010; // vC= -214 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111010011; // iC= 2003 
// vC = 14'b1111111010001011; // vC= -373 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001000; // iC= 2184 
// vC = 14'b1111111001110010; // vC= -398 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100001; // iC= 2145 
// vC = 14'b1111111101001100; // vC= -180 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b1111111001111001; // vC= -391 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b1111111011010111; // vC= -297 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101111; // iC= 2031 
// vC = 14'b1111111000110001; // vC= -463 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011111; // iC= 2079 
// vC = 14'b1111111011011000; // vC= -296 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b1111111101111110; // vC= -130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111011; // iC= 2043 
// vC = 14'b1111111100100100; // vC= -220 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111000; // iC= 1976 
// vC = 14'b1111111001100110; // vC= -410 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b1111111110010000; // vC= -112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100101; // iC= 2085 
// vC = 14'b1111111010011110; // vC= -354 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100101; // iC= 1957 
// vC = 14'b1111111100011100; // vC= -228 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100011; // iC= 1955 
// vC = 14'b1111111101111101; // vC= -131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101000; // iC= 2152 
// vC = 14'b1111111101000011; // vC= -189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111111110001101; // vC= -115 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100000; // iC= 2016 
// vC = 14'b1111111010100010; // vC= -350 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010011000; // iC= 2200 
// vC = 14'b1111111111000011; // vC=  -61 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101001; // iC= 1961 
// vC = 14'b1111111101111110; // vC= -130 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011000; // iC= 2008 
// vC = 14'b1111111110000011; // vC= -125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b1111111011001110; // vC= -306 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010100; // iC= 2196 
// vC = 14'b1111111100010100; // vC= -236 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111100; // iC= 2236 
// vC = 14'b1111111100001010; // vC= -246 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111100011; // iC= 2019 
// vC = 14'b1111111100000101; // vC= -251 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010111100; // iC= 2236 
// vC = 14'b1111111111100100; // vC=  -28 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001001; // iC= 2121 
// vC = 14'b0000000000100010; // vC=   34 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010010011; // iC= 2195 
// vC = 14'b1111111110011011; // vC= -101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110100; // iC= 2100 
// vC = 14'b1111111111011101; // vC=  -35 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010101111; // iC= 2223 
// vC = 14'b1111111101001111; // vC= -177 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011010; // iC= 1946 
// vC = 14'b1111111101010000; // vC= -176 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111001; // iC= 1977 
// vC = 14'b0000000001010010; // vC=   82 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110010; // iC= 2034 
// vC = 14'b1111111111110111; // vC=   -9 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110101; // iC= 2037 
// vC = 14'b1111111110000011; // vC= -125 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101011; // iC= 2027 
// vC = 14'b1111111101110001; // vC= -143 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100001; // iC= 2081 
// vC = 14'b1111111101000111; // vC= -185 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001010110; // iC= 2134 
// vC = 14'b1111111111111011; // vC=   -5 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011110; // iC= 2142 
// vC = 14'b0000000001111011; // vC=  123 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001111001; // iC= 2169 
// vC = 14'b0000000000101110; // vC=   46 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001101100; // iC= 2156 
// vC = 14'b0000000001111001; // vC=  121 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b1111111111111001; // vC=   -7 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011101; // iC= 1949 
// vC = 14'b0000000001100000; // vC=   96 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110000; // iC= 1904 
// vC = 14'b0000000000110010; // vC=   50 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000110110; // iC= 2102 
// vC = 14'b1111111111010110; // vC=  -42 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001110; // iC= 1998 
// vC = 14'b1111111111110011; // vC=  -13 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000001; // iC= 2177 
// vC = 14'b0000000011001001; // vC=  201 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b1111111111101010; // vC=  -22 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101010; // iC= 2026 
// vC = 14'b0000000011001100; // vC=  204 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011010; // iC= 2074 
// vC = 14'b0000000011010111; // vC=  215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010010; // iC= 2066 
// vC = 14'b0000000010100000; // vC=  160 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000010; // iC= 1922 
// vC = 14'b1111111111001110; // vC=  -50 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000110; // iC= 1990 
// vC = 14'b0000000001110010; // vC=  114 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011011; // iC= 2139 
// vC = 14'b0000000010111100; // vC=  188 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010001000; // iC= 2184 
// vC = 14'b0000000011110011; // vC=  243 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b0000000000100011; // vC=   35 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111111000; // iC= 2040 
// vC = 14'b0000000011101110; // vC=  238 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100000; // iC= 2144 
// vC = 14'b0000000000100011; // vC=   35 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101100; // iC= 2028 
// vC = 14'b0000000001100010; // vC=   98 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000111110; // iC= 2110 
// vC = 14'b0000000011000101; // vC=  197 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000100111; // iC= 2087 
// vC = 14'b0000000011000111; // vC=  199 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010011; // iC= 1875 
// vC = 14'b0000000100100100; // vC=  292 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011010; // iC= 2010 
// vC = 14'b0000000100100110; // vC=  294 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100111; // iC= 2151 
// vC = 14'b0000000010010100; // vC=  148 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110000000; // iC= 1920 
// vC = 14'b0000000010001001; // vC=  137 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001100011; // iC= 2147 
// vC = 14'b0000000101111000; // vC=  376 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100010000111; // iC= 2183 
// vC = 14'b0000000010000011; // vC=  131 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000000; // iC= 1984 
// vC = 14'b0000000101010101; // vC=  341 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001011100; // iC= 2140 
// vC = 14'b0000000010001101; // vC=  141 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000011; // iC= 2051 
// vC = 14'b0000000101001100; // vC=  332 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001111; // iC= 1871 
// vC = 14'b0000000011101010; // vC=  234 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011111; // iC= 1951 
// vC = 14'b0000000001111000; // vC=  120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111001000; // iC= 1992 
// vC = 14'b0000000001101111; // vC=  111 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000111; // iC= 2119 
// vC = 14'b0000000101001011; // vC=  331 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011100; // iC= 1884 
// vC = 14'b0000000101110010; // vC=  370 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000000000; // iC= 2048 
// vC = 14'b0000000110000101; // vC=  389 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110110001; // iC= 1969 
// vC = 14'b0000000110001001; // vC=  393 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001011; // iC= 1867 
// vC = 14'b0000000100011001; // vC=  281 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b0000000101010111; // vC=  343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000010; // iC= 2114 
// vC = 14'b0000000111101001; // vC=  489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111010; // iC= 1914 
// vC = 14'b0000000110100000; // vC=  416 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101001111; // iC= 1871 
// vC = 14'b0000000100010010; // vC=  274 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101100; // iC= 1836 
// vC = 14'b0000001000001000; // vC=  520 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001100; // iC= 2124 
// vC = 14'b0000000101001001; // vC=  329 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001011; // iC= 2123 
// vC = 14'b0000000011110111; // vC=  247 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000010; // iC= 2114 
// vC = 14'b0000000100000101; // vC=  261 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b0000000111011001; // vC=  473 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011101; // iC= 2077 
// vC = 14'b0000000111011000; // vC=  472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111011101; // iC= 2013 
// vC = 14'b0000000100101100; // vC=  300 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000010011; // iC= 2067 
// vC = 14'b0000000111111011; // vC=  507 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110111; // iC= 1911 
// vC = 14'b0000000110100010; // vC=  418 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111010; // iC= 1850 
// vC = 14'b0000000110001010; // vC=  394 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001001011; // iC= 2123 
// vC = 14'b0000000111100110; // vC=  486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100000011011; // iC= 2075 
// vC = 14'b0000000111011010; // vC=  474 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011010; // iC= 1882 
// vC = 14'b0000001000010110; // vC=  534 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000010; // iC= 1858 
// vC = 14'b0000000111111101; // vC=  509 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101011; // iC= 1835 
// vC = 14'b0000000110011011; // vC=  411 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110111111; // iC= 1983 
// vC = 14'b0000000110010000; // vC=  400 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010100; // iC= 1812 
// vC = 14'b0000000110111001; // vC=  441 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000100001000001; // iC= 2113 
// vC = 14'b0000000111001001; // vC=  457 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b0000000111000001; // vC=  449 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110101; // iC= 1781 
// vC = 14'b0000001001011000; // vC=  600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010000; // iC= 1936 
// vC = 14'b0000000111011010; // vC=  474 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101110; // iC= 1838 
// vC = 14'b0000001000000000; // vC=  512 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110100; // iC= 1908 
// vC = 14'b0000000111000010; // vC=  450 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011000; // iC= 1880 
// vC = 14'b0000001000101000; // vC=  552 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100011; // iC= 1955 
// vC = 14'b0000001001011010; // vC=  602 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101100; // iC= 1964 
// vC = 14'b0000000111010110; // vC=  470 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011011; // iC= 1819 
// vC = 14'b0000001011010010; // vC=  722 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011011; // iC= 1883 
// vC = 14'b0000001000011010; // vC=  538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101110101; // iC= 1909 
// vC = 14'b0000001001010001; // vC=  593 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101000; // iC= 1960 
// vC = 14'b0000000111000100; // vC=  452 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b0000001010111010; // vC=  698 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110001001; // iC= 1929 
// vC = 14'b0000000111101110; // vC=  494 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101111101; // iC= 1917 
// vC = 14'b0000001011111110; // vC=  766 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010110; // iC= 1942 
// vC = 14'b0000001000100000; // vC=  544 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110001; // iC= 2033 
// vC = 14'b0000001011100001; // vC=  737 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111101101; // iC= 2029 
// vC = 14'b0000001100011001; // vC=  793 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011010100; // iC= 1748 
// vC = 14'b0000001010010010; // vC=  658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111110010; // iC= 2034 
// vC = 14'b0000001010010001; // vC=  657 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100111; // iC= 1959 
// vC = 14'b0000001000010001; // vC=  529 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101101; // iC= 1965 
// vC = 14'b0000001011100101; // vC=  741 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011010; // iC= 1882 
// vC = 14'b0000001011101010; // vC=  746 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011001; // iC= 1945 
// vC = 14'b0000001001110100; // vC=  628 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110101011; // iC= 1963 
// vC = 14'b0000001011110111; // vC=  759 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100000100; // iC= 1796 
// vC = 14'b0000001101000010; // vC=  834 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110010; // iC= 1714 
// vC = 14'b0000001001010101; // vC=  597 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100011; // iC= 1827 
// vC = 14'b0000001100111000; // vC=  824 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011111; // iC= 1759 
// vC = 14'b0000001101100001; // vC=  865 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110011011; // iC= 1947 
// vC = 14'b0000001100101000; // vC=  808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011111000001; // iC= 1985 
// vC = 14'b0000001011101101; // vC=  749 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110010100; // iC= 1940 
// vC = 14'b0000001101111111; // vC=  895 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101110; // iC= 1710 
// vC = 14'b0000001010110011; // vC=  691 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010010; // iC= 1810 
// vC = 14'b0000001010001001; // vC=  649 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101111; // iC= 1711 
// vC = 14'b0000001011110011; // vC=  755 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110000; // iC= 1840 
// vC = 14'b0000001110011010; // vC=  922 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110111; // iC= 1847 
// vC = 14'b0000001011011000; // vC=  728 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100000; // iC= 1888 
// vC = 14'b0000001010100100; // vC=  676 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100011001; // iC= 1817 
// vC = 14'b0000001101001110; // vC=  846 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000000; // iC= 1664 
// vC = 14'b0000001010010110; // vC=  662 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011110100000; // iC= 1952 
// vC = 14'b0000001110001010; // vC=  906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011110101; // iC= 1781 
// vC = 14'b0000001011001111; // vC=  719 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000111; // iC= 1671 
// vC = 14'b0000001101111101; // vC=  893 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101000111; // iC= 1863 
// vC = 14'b0000001011110000; // vC=  752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100111; // iC= 1703 
// vC = 14'b0000001110000100; // vC=  900 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001000; // iC= 1736 
// vC = 14'b0000001101010000; // vC=  848 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101010000; // iC= 1872 
// vC = 14'b0000001100111011; // vC=  827 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100000; // iC= 1696 
// vC = 14'b0000001111111010; // vC= 1018 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100101; // iC= 1701 
// vC = 14'b0000001100000001; // vC=  769 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111101; // iC= 1853 
// vC = 14'b0000001101100011; // vC=  867 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100010; // iC= 1634 
// vC = 14'b0000001110011011; // vC=  923 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001110110; // iC= 1654 
// vC = 14'b0000001111101111; // vC= 1007 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011100; // iC= 1884 
// vC = 14'b0000001110001001; // vC=  905 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100010001; // iC= 1809 
// vC = 14'b0000001110000010; // vC=  898 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111010; // iC= 1658 
// vC = 14'b0000001101100100; // vC=  868 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101100011; // iC= 1891 
// vC = 14'b0000010001001111; // vC= 1103 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011001100; // iC= 1740 
// vC = 14'b0000001101111000; // vC=  888 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000100; // iC= 1668 
// vC = 14'b0000001100110010; // vC=  818 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100110; // iC= 1830 
// vC = 14'b0000001111000111; // vC=  967 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011101011010; // iC= 1882 
// vC = 14'b0000001110001110; // vC=  910 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000110; // iC= 1606 
// vC = 14'b0000001101011010; // vC=  858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100101; // iC= 1765 
// vC = 14'b0000010000100011; // vC= 1059 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110101; // iC= 1845 
// vC = 14'b0000001101101011; // vC=  875 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100000; // iC= 1696 
// vC = 14'b0000001111010111; // vC=  983 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111000; // iC= 1656 
// vC = 14'b0000010010010110; // vC= 1174 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011100111; // iC= 1767 
// vC = 14'b0000001110101100; // vC=  940 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100101000; // iC= 1832 
// vC = 14'b0000010001011000; // vC= 1112 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001001100; // iC= 1612 
// vC = 14'b0000001101100101; // vC=  869 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001111; // iC= 1551 
// vC = 14'b0000001111011101; // vC=  989 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100111011; // iC= 1851 
// vC = 14'b0000010001001100; // vC= 1100 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111000; // iC= 1656 
// vC = 14'b0000001110110110; // vC=  950 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100110011; // iC= 1843 
// vC = 14'b0000010000111000; // vC= 1080 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111011; // iC= 1659 
// vC = 14'b0000001111010011; // vC=  979 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011100100100; // iC= 1828 
// vC = 14'b0000010011010101; // vC= 1237 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000010; // iC= 1538 
// vC = 14'b0000001111010110; // vC=  982 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000000000; // iC= 1536 
// vC = 14'b0000010001000111; // vC= 1095 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011101; // iC= 1757 
// vC = 14'b0000001110110001; // vC=  945 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011001; // iC= 1561 
// vC = 14'b0000010000001101; // vC= 1037 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111111; // iC= 1791 
// vC = 14'b0000010011000010; // vC= 1218 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011011110; // iC= 1758 
// vC = 14'b0000010011000011; // vC= 1219 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111000; // iC= 1784 
// vC = 14'b0000010000010001; // vC= 1041 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111010; // iC= 1530 
// vC = 14'b0000010011101000; // vC= 1256 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000011010; // iC= 1562 
// vC = 14'b0000010100001100; // vC= 1292 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011011111100; // iC= 1788 
// vC = 14'b0000010000000101; // vC= 1029 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111010; // iC= 1594 
// vC = 14'b0000010001101100; // vC= 1132 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110001; // iC= 1521 
// vC = 14'b0000010000001010; // vC= 1034 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111110; // iC= 1662 
// vC = 14'b0000010001001101; // vC= 1101 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001100100; // iC= 1636 
// vC = 14'b0000010000101001; // vC= 1065 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010000; // iC= 1616 
// vC = 14'b0000010010101101; // vC= 1197 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011100; // iC= 1692 
// vC = 14'b0000010011001110; // vC= 1230 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100110; // iC= 1702 
// vC = 14'b0000010001100001; // vC= 1121 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001100; // iC= 1548 
// vC = 14'b0000010010100101; // vC= 1189 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010000001; // iC= 1665 
// vC = 14'b0000010010011111; // vC= 1183 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000111011; // iC= 1595 
// vC = 14'b0000010011011010; // vC= 1242 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001010111; // iC= 1623 
// vC = 14'b0000010100100111; // vC= 1319 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010110100; // iC= 1716 
// vC = 14'b0000010000111010; // vC= 1082 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010011000; // iC= 1688 
// vC = 14'b0000010010101010; // vC= 1194 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001100; // iC= 1484 
// vC = 14'b0000010100101110; // vC= 1326 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001001; // iC= 1673 
// vC = 14'b0000010001101000; // vC= 1128 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010010; // iC= 1490 
// vC = 14'b0000010010111010; // vC= 1210 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010100000; // iC= 1696 
// vC = 14'b0000010011001100; // vC= 1228 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010001110; // iC= 1678 
// vC = 14'b0000010010111111; // vC= 1215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011010101010; // iC= 1706 
// vC = 14'b0000010001100000; // vC= 1120 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101100; // iC= 1452 
// vC = 14'b0000010101010010; // vC= 1362 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111010101; // iC= 1493 
// vC = 14'b0000010011001100; // vC= 1228 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111101; // iC= 1533 
// vC = 14'b0000010100101001; // vC= 1321 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100101; // iC= 1445 
// vC = 14'b0000010010111000; // vC= 1208 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101110101; // iC= 1397 
// vC = 14'b0000010011010010; // vC= 1234 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000100100; // iC= 1572 
// vC = 14'b0000010010100100; // vC= 1188 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001100; // iC= 1548 
// vC = 14'b0000010101010010; // vC= 1362 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001111101; // iC= 1661 
// vC = 14'b0000010010111111; // vC= 1215 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101110; // iC= 1390 
// vC = 14'b0000010011011101; // vC= 1245 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111111010; // iC= 1530 
// vC = 14'b0000010101101111; // vC= 1391 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011010; // iC= 1434 
// vC = 14'b0000010011000110; // vC= 1222 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001011011; // iC= 1627 
// vC = 14'b0000010011010011; // vC= 1235 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011001000010; // iC= 1602 
// vC = 14'b0000010101110000; // vC= 1392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001110; // iC= 1422 
// vC = 14'b0000010100111111; // vC= 1343 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101111; // iC= 1327 
// vC = 14'b0000010111001110; // vC= 1486 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110011111; // iC= 1439 
// vC = 14'b0000010100011101; // vC= 1309 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000000; // iC= 1408 
// vC = 14'b0000010011000111; // vC= 1223 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000011; // iC= 1475 
// vC = 14'b0000010011001111; // vC= 1231 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111100; // iC= 1340 
// vC = 14'b0000010110011101; // vC= 1437 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111011; // iC= 1403 
// vC = 14'b0000010101110000; // vC= 1392 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011011; // iC= 1307 
// vC = 14'b0000010100010110; // vC= 1302 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110001; // iC= 1521 
// vC = 14'b0000010011111011; // vC= 1275 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100010; // iC= 1314 
// vC = 14'b0000010111000000; // vC= 1472 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111110001; // iC= 1521 
// vC = 14'b0000010100101000; // vC= 1320 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000101001; // iC= 1577 
// vC = 14'b0000010100110010; // vC= 1330 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110101; // iC= 1269 
// vC = 14'b0000010101101011; // vC= 1387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101001; // iC= 1321 
// vC = 14'b0000010110110000; // vC= 1456 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100100; // iC= 1316 
// vC = 14'b0000010111011000; // vC= 1496 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100000100; // iC= 1284 
// vC = 14'b0000010110111001; // vC= 1465 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000011000001001; // iC= 1545 
// vC = 14'b0000010110000101; // vC= 1413 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111001010; // iC= 1482 
// vC = 14'b0000010100100111; // vC= 1319 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110001101; // iC= 1421 
// vC = 14'b0000011001001010; // vC= 1610 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010001; // iC= 1361 
// vC = 14'b0000010101011100; // vC= 1372 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000011; // iC= 1475 
// vC = 14'b0000010110011100; // vC= 1436 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100100010; // iC= 1314 
// vC = 14'b0000010101101011; // vC= 1387 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101100100; // iC= 1380 
// vC = 14'b0000010101101010; // vC= 1386 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011010101; // iC= 1237 
// vC = 14'b0000010111111000; // vC= 1528 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110101110; // iC= 1454 
// vC = 14'b0000010111111000; // vC= 1528 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100011101; // iC= 1309 
// vC = 14'b0000011001000000; // vC= 1600 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101111000; // iC= 1400 
// vC = 14'b0000011000110000; // vC= 1584 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100100; // iC= 1444 
// vC = 14'b0000011000001010; // vC= 1546 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011110111; // iC= 1271 
// vC = 14'b0000011001100011; // vC= 1635 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011101; // iC= 1181 
// vC = 14'b0000011000000010; // vC= 1538 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110111100; // iC= 1468 
// vC = 14'b0000010111100100; // vC= 1508 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000000; // iC= 1472 
// vC = 14'b0000010111011111; // vC= 1503 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100011; // iC= 1251 
// vC = 14'b0000011001101110; // vC= 1646 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010111000110; // iC= 1478 
// vC = 14'b0000010111001000; // vC= 1480 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000011; // iC= 1411 
// vC = 14'b0000010101111111; // vC= 1407 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110000000; // iC= 1408 
// vC = 14'b0000010101111101; // vC= 1405 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010000000; // iC= 1152 
// vC = 14'b0000011000011110; // vC= 1566 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010110100110; // iC= 1446 
// vC = 14'b0000010111101011; // vC= 1515 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101101010; // iC= 1386 
// vC = 14'b0000011001111010; // vC= 1658 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111011; // iC= 1339 
// vC = 14'b0000011010001000; // vC= 1672 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100001001; // iC= 1289 
// vC = 14'b0000011000111111; // vC= 1599 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110011; // iC= 1331 
// vC = 14'b0000011000110011; // vC= 1587 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010111; // iC= 1367 
// vC = 14'b0000011011000011; // vC= 1731 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101110; // iC= 1134 
// vC = 14'b0000011001001000; // vC= 1608 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100001; // iC= 1121 
// vC = 14'b0000010111111001; // vC= 1529 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101010010; // iC= 1362 
// vC = 14'b0000011000110110; // vC= 1590 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010101011; // iC= 1195 
// vC = 14'b0000010110111111; // vC= 1471 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100110001; // iC= 1329 
// vC = 14'b0000011000110010; // vC= 1586 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011101; // iC= 1117 
// vC = 14'b0000011011111111; // vC= 1791 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010010101; // iC= 1173 
// vC = 14'b0000011011111000; // vC= 1784 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100110; // iC= 1190 
// vC = 14'b0000011011001101; // vC= 1741 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000111001; // iC= 1081 
// vC = 14'b0000011011000100; // vC= 1732 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001001100; // iC= 1100 
// vC = 14'b0000010111010001; // vC= 1489 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100111001; // iC= 1337 
// vC = 14'b0000011010111010; // vC= 1722 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010101001100; // iC= 1356 
// vC = 14'b0000011001100100; // vC= 1636 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101111; // iC= 1071 
// vC = 14'b0000011000010011; // vC= 1555 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011100011; // iC= 1251 
// vC = 14'b0000011011100101; // vC= 1765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000101010; // iC= 1066 
// vC = 14'b0000011001110100; // vC= 1652 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010100101010; // iC= 1322 
// vC = 14'b0000011011011010; // vC= 1754 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001010010; // iC= 1106 
// vC = 14'b0000011000011100; // vC= 1564 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110001; // iC= 1137 
// vC = 14'b0000011011100101; // vC= 1765 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100011; // iC=  995 
// vC = 14'b0000011000000101; // vC= 1541 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011010; // iC= 1178 
// vC = 14'b0000011010010001; // vC= 1681 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110110; // iC= 1142 
// vC = 14'b0000011000001111; // vC= 1551 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110100; // iC= 1012 
// vC = 14'b0000011011101100; // vC= 1772 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010000; // iC= 1040 
// vC = 14'b0000011100111111; // vC= 1855 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010111; // iC= 1047 
// vC = 14'b0000011011001000; // vC= 1736 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101101; // iC= 1133 
// vC = 14'b0000011000011011; // vC= 1563 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011101101; // iC= 1261 
// vC = 14'b0000011000100100; // vC= 1572 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111010011; // iC=  979 
// vC = 14'b0000011101100010; // vC= 1890 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111100101; // iC=  997 
// vC = 14'b0000011010001011; // vC= 1675 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010011000010; // iC= 1218 
// vC = 14'b0000011001001011; // vC= 1611 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001101110; // iC= 1134 
// vC = 14'b0000011010000100; // vC= 1668 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100010; // iC= 1122 
// vC = 14'b0000011100001010; // vC= 1802 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001101; // iC= 1037 
// vC = 14'b0000011001010001; // vC= 1617 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010011001; // iC= 1177 
// vC = 14'b0000011010111101; // vC= 1725 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001011; // iC= 1035 
// vC = 14'b0000011010100100; // vC= 1700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011010; // iC=  986 
// vC = 14'b0000011011110110; // vC= 1782 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001110100; // iC= 1140 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000001001; // iC= 1033 
// vC = 14'b0000011011010011; // vC= 1747 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110110; // iC=  886 
// vC = 14'b0000011101110010; // vC= 1906 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010010100110; // iC= 1190 
// vC = 14'b0000011010100100; // vC= 1700 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001100001; // iC= 1121 
// vC = 14'b0000011100110101; // vC= 1845 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101000; // iC= 1000 
// vC = 14'b0000011001110011; // vC= 1651 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010111; // iC= 1047 
// vC = 14'b0000011101101101; // vC= 1901 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110100; // iC=  884 
// vC = 14'b0000011010010011; // vC= 1683 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000110; // iC= 1030 
// vC = 14'b0000011110000101; // vC= 1925 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111000; // iC= 1016 
// vC = 14'b0000011110000111; // vC= 1927 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010001011011; // iC= 1115 
// vC = 14'b0000011010111100; // vC= 1724 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111110011; // iC= 1011 
// vC = 14'b0000011010100000; // vC= 1696 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101100010; // iC=  866 
// vC = 14'b0000011110001111; // vC= 1935 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111001; // iC=  825 
// vC = 14'b0000011011011000; // vC= 1752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001011; // iC=  907 
// vC = 14'b0000011010000111; // vC= 1671 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000010111; // iC= 1047 
// vC = 14'b0000011010001110; // vC= 1678 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000011111; // iC= 1055 
// vC = 14'b0000011010001111; // vC= 1679 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111000011; // iC=  963 
// vC = 14'b0000011100111100; // vC= 1852 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111011111; // iC=  991 
// vC = 14'b0000011011011000; // vC= 1752 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111011; // iC= 1019 
// vC = 14'b0000011011100100; // vC= 1764 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110011010; // iC=  922 
// vC = 14'b0000011100010010; // vC= 1810 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101000; // iC=  936 
// vC = 14'b0000011010100101; // vC= 1701 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111111; // iC=  831 
// vC = 14'b0000011100100001; // vC= 1825 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000010000000000; // iC= 1024 
// vC = 14'b0000011011000001; // vC= 1729 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101100; // iC=  940 
// vC = 14'b0000011101101110; // vC= 1902 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000010; // iC=  898 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111111010; // iC= 1018 
// vC = 14'b0000011101001111; // vC= 1871 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011111111; // iC=  767 
// vC = 14'b0000011101000010; // vC= 1858 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110101001; // iC=  937 
// vC = 14'b0000011110111111; // vC= 1983 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011110001; // iC=  753 
// vC = 14'b0000011010110110; // vC= 1718 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101001; // iC= 1001 
// vC = 14'b0000011111010111; // vC= 2007 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001111101111; // iC= 1007 
// vC = 14'b0000011101011111; // vC= 1887 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110100001; // iC=  929 
// vC = 14'b0000011100010000; // vC= 1808 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011011; // iC=  731 
// vC = 14'b0000011101101110; // vC= 1902 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110000011; // iC=  899 
// vC = 14'b0000011100111010; // vC= 1850 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100010111; // iC=  791 
// vC = 14'b0000011011001111; // vC= 1743 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011011; // iC=  795 
// vC = 14'b0000011110110111; // vC= 1975 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011000001; // iC=  705 
// vC = 14'b0000011111010011; // vC= 2003 
// sigma = 2'b01; // sigma=01 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110101; // iC=  885 
// vC = 14'b0000011100100010; // vC= 1826 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100110; // iC=  678 
// vC = 14'b0000011101011110; // vC= 1886 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011100111; // iC=  743 
// vC = 14'b0000011111111111; // vC= 2047 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001111; // iC=  911 
// vC = 14'b0000011100011101; // vC= 1821 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010000101; // iC=  645 
// vC = 14'b0000011111011100; // vC= 2012 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111010; // iC=  634 
// vC = 14'b0000011110101010; // vC= 1962 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100111011; // iC=  827 
// vC = 14'b0000011111110101; // vC= 2037 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101001111; // iC=  847 
// vC = 14'b0000011110100100; // vC= 1956 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111001; // iC=  633 
// vC = 14'b0000011011101111; // vC= 1775 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001110001011; // iC=  907 
// vC = 14'b0000011101001010; // vC= 1866 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001100110; // iC=  614 
// vC = 14'b0000011100001101; // vC= 1805 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001100; // iC=  780 
// vC = 14'b0000011111100001; // vC= 2017 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011001011; // iC=  715 
// vC = 14'b0000011110110111; // vC= 1975 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001101110110; // iC=  886 
// vC = 14'b0000011110011011; // vC= 1947 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101001; // iC=  681 
// vC = 14'b0000011101101000; // vC= 1896 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001111111; // iC=  639 
// vC = 14'b0000100000110101; // vC= 2101 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100101; // iC=  549 
// vC = 14'b0000011100000101; // vC= 1797 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100011101; // iC=  797 
// vC = 14'b0000011110101110; // vC= 1966 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001110010; // iC=  626 
// vC = 14'b0000011111100001; // vC= 2017 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011101101; // iC=  749 
// vC = 14'b0000100001000101; // vC= 2117 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001001100; // iC=  588 
// vC = 14'b0000100000000000; // vC= 2048 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100001011; // iC=  779 
// vC = 14'b0000011110110001; // vC= 1969 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011010; // iC=  666 
// vC = 14'b0000011111001010; // vC= 1994 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001101100; // iC=  620 
// vC = 14'b0000011100011111; // vC= 1823 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001100000101; // iC=  773 
// vC = 14'b0000100000110101; // vC= 2101 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101100; // iC=  684 
// vC = 14'b0000011110101000; // vC= 1960 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010011111; // iC=  671 
// vC = 14'b0000100001000111; // vC= 2119 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010101000; // iC=  680 
// vC = 14'b0000011101101001; // vC= 1897 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001011011101; // iC=  733 
// vC = 14'b0000011100011110; // vC= 1822 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010100000; // iC=  672 
// vC = 14'b0000011101110101; // vC= 1909 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001010001000; // iC=  648 
// vC = 14'b0000100000001001; // vC= 2057 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001000010; // iC=  578 
// vC = 14'b0000100001100100; // vC= 2148 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000100001; // iC=  545 
// vC = 14'b0000011100111110; // vC= 1854 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110010101; // iC=  405 
// vC = 14'b0000011100101110; // vC= 1838 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101110111; // iC=  375 
// vC = 14'b0000100001011111; // vC= 2143 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000010100; // iC=  532 
// vC = 14'b0000011111001011; // vC= 1995 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001001011001; // iC=  601 
// vC = 14'b0000011101001110; // vC= 1870 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111011011; // iC=  475 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111110100; // iC=  500 
// vC = 14'b0000011111011110; // vC= 2014 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000001000110010; // iC=  562 
// vC = 14'b0000100001011110; // vC= 2142 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000111101100; // iC=  492 
// vC = 14'b0000100001000000; // vC= 2112 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000110101001; // iC=  425 
// vC = 14'b0000011101100001; // vC= 1889 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100001; // iC=  225 
// vC = 14'b0000011101101101; // vC= 1901 
// sigma = 2'b00; // sigma=00 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101100101; // iC=  357 
// vC = 14'b0000011100111001; // vC= 1849 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100010101; // iC=  277 
// vC = 14'b0000011110101000; // vC= 1960 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100011111; // iC=  287 
// vC = 14'b0000011101010000; // vC= 1872 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101001; // iC=  361 
// vC = 14'b0000011110110110; // vC= 1974 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100110010; // iC=  306 
// vC = 14'b0000100000110100; // vC= 2100 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011001111; // iC=  207 
// vC = 14'b0000011110011111; // vC= 1951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101001011; // iC=  331 
// vC = 14'b0000100001101101; // vC= 2157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101101101; // iC=  365 
// vC = 14'b0000011110101101; // vC= 1965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111101; // iC=  253 
// vC = 14'b0000100000011111; // vC= 2079 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000101000001; // iC=  321 
// vC = 14'b0000011110000000; // vC= 1920 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000100101011; // iC=  299 
// vC = 14'b0000011111110001; // vC= 2033 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001100001; // iC=   97 
// vC = 14'b0000100001010100; // vC= 2132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100001; // iC=   33 
// vC = 14'b0000011101011000; // vC= 1880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010011010; // iC=  154 
// vC = 14'b0000011101111100; // vC= 1916 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011111001; // iC=  249 
// vC = 14'b0000100001110100; // vC= 2164 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000011100000; // iC=  224 
// vC = 14'b0000011111000110; // vC= 1990 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010010011; // iC=  147 
// vC = 14'b0000100001110110; // vC= 2166 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001101000; // iC=  104 
// vC = 14'b0000011110110011; // vC= 1971 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111000110; // iC=  -58 
// vC = 14'b0000011111111011; // vC= 2043 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000001; // iC= -127 
// vC = 14'b0000011101001101; // vC= 1869 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000010110000; // iC=  176 
// vC = 14'b0000011101010011; // vC= 1875 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000111011; // iC=   59 
// vC = 14'b0000011111100011; // vC= 2019 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010110; // iC=   22 
// vC = 14'b0000011101101110; // vC= 1902 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000001011011; // iC=   91 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000100000; // iC=   32 
// vC = 14'b0000100010000010; // vC= 2178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b0000000000010101; // iC=   21 
// vC = 14'b0000100000000111; // vC= 2055 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111110000101; // iC= -123 
// vC = 14'b0000100000101111; // vC= 2095 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111111011111; // iC=  -33 
// vC = 14'b0000011110000100; // vC= 1924 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010101; // iC= -235 
// vC = 14'b0000011101010110; // vC= 1878 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100010110; // iC= -234 
// vC = 14'b0000100001111010; // vC= 2170 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100110101; // iC= -203 
// vC = 14'b0000100001000101; // vC= 2117 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111010010100; // iC= -364 
// vC = 14'b0000100000100111; // vC= 2087 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111100001100; // iC= -244 
// vC = 14'b0000100000101010; // vC= 2090 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111000; // iC= -392 
// vC = 14'b0000011111000101; // vC= 1989 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111101110100; // iC= -140 
// vC = 14'b0000100000110110; // vC= 2102 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011010110; // iC= -298 
// vC = 14'b0000100001010101; // vC= 2133 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011011111; // iC= -289 
// vC = 14'b0000011110011111; // vC= 1951 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000111010; // iC= -454 
// vC = 14'b0000011110111101; // vC= 1981 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100101; // iC= -539 
// vC = 14'b0000011101101000; // vC= 1896 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111100100; // iC= -540 
// vC = 14'b0000011110110100; // vC= 1972 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110000; // iC= -400 
// vC = 14'b0000011110011110; // vC= 1950 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111011000111; // iC= -313 
// vC = 14'b0000011110100000; // vC= 1952 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110011100; // iC= -612 
// vC = 14'b0000011111000100; // vC= 1988 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001111110; // iC= -386 
// vC = 14'b0000011111111001; // vC= 2041 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110111110001; // iC= -527 
// vC = 14'b0000011100111000; // vC= 1848 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111001110101; // iC= -395 
// vC = 14'b0000100000001101; // vC= 2061 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111111000000100; // iC= -508 
// vC = 14'b0000011110011011; // vC= 1947 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110111111; // iC= -577 
// vC = 14'b0000100000101000; // vC= 2088 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100110; // iC= -730 
// vC = 14'b0000100000111000; // vC= 2104 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101100111; // iC= -665 
// vC = 14'b0000100000001111; // vC= 2063 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110110001010; // iC= -630 
// vC = 14'b0000011110010100; // vC= 1940 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001111; // iC= -689 
// vC = 14'b0000011110101111; // vC= 1967 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010011111; // iC= -865 
// vC = 14'b0000100000100011; // vC= 2083 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011100001; // iC= -799 
// vC = 14'b0000011101110001; // vC= 1905 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010101010; // iC= -854 
// vC = 14'b0000011110101011; // vC= 1963 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101001011; // iC= -693 
// vC = 14'b0000011110100000; // vC= 1952 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010100001; // iC= -863 
// vC = 14'b0000100000000000; // vC= 2048 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110101000111; // iC= -697 
// vC = 14'b0000011101000101; // vC= 1861 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011101001; // iC= -791 
// vC = 14'b0000011101111001; // vC= 1913 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110011011100; // iC= -804 
// vC = 14'b0000011111101010; // vC= 2026 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110100100001; // iC= -735 
// vC = 14'b0000011100110001; // vC= 1841 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010110110; // iC= -842 
// vC = 14'b0000011100010100; // vC= 1812 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111000011; // iC=-1085 
// vC = 14'b0000011101110111; // vC= 1911 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101111100100; // iC=-1052 
// vC = 14'b0000011111011101; // vC= 2013 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110010111110; // iC= -834 
// vC = 14'b0000011100000011; // vC= 1795 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110000010000; // iC=-1008 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110100000; // iC=-1120 
// vC = 14'b0000011100101101; // vC= 1837 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001000100; // iC= -956 
// vC = 14'b0000011011011110; // vC= 1758 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111110001010000; // iC= -944 
// vC = 14'b0000011111110101; // vC= 2037 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100101100; // iC=-1236 
// vC = 14'b0000011111011101; // vC= 2013 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100001; // iC=-1183 
// vC = 14'b0000011110101101; // vC= 1965 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110111010; // iC=-1094 
// vC = 14'b0000011110111000; // vC= 1976 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110010100; // iC=-1132 
// vC = 14'b0000011110111011; // vC= 1979 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110110; // iC=-1290 
// vC = 14'b0000011101000011; // vC= 1859 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101010111; // iC=-1193 
// vC = 14'b0000011100001011; // vC= 1803 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010111; // iC=-1321 
// vC = 14'b0000011110011101; // vC= 1949 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101110000010; // iC=-1150 
// vC = 14'b0000011111001010; // vC= 1994 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100100111; // iC=-1241 
// vC = 14'b0000011101100101; // vC= 1893 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011010; // iC=-1190 
// vC = 14'b0000011110111011; // vC= 1979 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100000; // iC=-1376 
// vC = 14'b0000011110111110; // vC= 1982 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101100111; // iC=-1177 
// vC = 14'b0000011011010010; // vC= 1746 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011111010; // iC=-1286 
// vC = 14'b0000011010001101; // vC= 1677 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010010; // iC=-1262 
// vC = 14'b0000011010101100; // vC= 1708 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100011011; // iC=-1253 
// vC = 14'b0000011001111111; // vC= 1663 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100010011; // iC=-1261 
// vC = 14'b0000011010000100; // vC= 1668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011000111; // iC=-1337 
// vC = 14'b0000011010110010; // vC= 1714 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010110000; // iC=-1360 
// vC = 14'b0000011101101011; // vC= 1899 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110110; // iC=-1418 
// vC = 14'b0000011101101000; // vC= 1896 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000011000; // iC=-1512 
// vC = 14'b0000011100101100; // vC= 1836 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101001; // iC=-1559 
// vC = 14'b0000011010000000; // vC= 1664 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110110; // iC=-1418 
// vC = 14'b0000011001110010; // vC= 1650 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101111; // iC=-1553 
// vC = 14'b0000011100100010; // vC= 1826 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011101; // iC=-1635 
// vC = 14'b0000011100001001; // vC= 1801 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000010; // iC=-1470 
// vC = 14'b0000011101001000; // vC= 1864 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111111; // iC=-1537 
// vC = 14'b0000011000111100; // vC= 1596 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111111010; // iC=-1542 
// vC = 14'b0000011001111001; // vC= 1657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010011; // iC=-1645 
// vC = 14'b0000011100010111; // vC= 1815 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101001; // iC=-1623 
// vC = 14'b0000011000110010; // vC= 1586 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100111; // iC=-1433 
// vC = 14'b0000011000111111; // vC= 1599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110011001; // iC=-1639 
// vC = 14'b0000011010101011; // vC= 1707 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111000; // iC=-1736 
// vC = 14'b0000011010000011; // vC= 1667 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101011; // iC=-1685 
// vC = 14'b0000011011110011; // vC= 1779 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110011; // iC=-1741 
// vC = 14'b0000011100011110; // vC= 1822 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110110; // iC=-1802 
// vC = 14'b0000011000110101; // vC= 1589 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100001; // iC=-1567 
// vC = 14'b0000011001101110; // vC= 1646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010111; // iC=-1577 
// vC = 14'b0000011100011111; // vC= 1823 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101001; // iC=-1687 
// vC = 14'b0000011001100001; // vC= 1633 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101001; // iC=-1751 
// vC = 14'b0000011010011110; // vC= 1694 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001011; // iC=-1589 
// vC = 14'b0000011011001111; // vC= 1743 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100000; // iC=-1760 
// vC = 14'b0000011000110001; // vC= 1585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100010; // iC=-1822 
// vC = 14'b0000010111011111; // vC= 1503 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000011; // iC=-1853 
// vC = 14'b0000010111000101; // vC= 1477 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101101; // iC=-1811 
// vC = 14'b0000011010011101; // vC= 1693 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110001; // iC=-1615 
// vC = 14'b0000010111111110; // vC= 1534 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101110; // iC=-1874 
// vC = 14'b0000010111101101; // vC= 1517 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101101; // iC=-1747 
// vC = 14'b0000011010110000; // vC= 1712 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001110; // iC=-1650 
// vC = 14'b0000011000101010; // vC= 1578 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000111; // iC=-1657 
// vC = 14'b0000011000101111; // vC= 1583 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011101; // iC=-1763 
// vC = 14'b0000010110001011; // vC= 1419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010001; // iC=-1903 
// vC = 14'b0000011001011110; // vC= 1630 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101011; // iC=-1685 
// vC = 14'b0000010111110001; // vC= 1521 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101011; // iC=-1749 
// vC = 14'b0000010110111010; // vC= 1466 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010110; // iC=-1706 
// vC = 14'b0000010111100111; // vC= 1511 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000110; // iC=-1914 
// vC = 14'b0000010101101001; // vC= 1385 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101101; // iC=-1811 
// vC = 14'b0000011001111010; // vC= 1658 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101010; // iC=-1942 
// vC = 14'b0000010110000110; // vC= 1414 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011111; // iC=-1953 
// vC = 14'b0000011000100000; // vC= 1568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b0000010101111000; // vC= 1400 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101010; // iC=-1814 
// vC = 14'b0000010100110110; // vC= 1334 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b0000010101001101; // vC= 1357 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110110; // iC=-2058 
// vC = 14'b0000010101011111; // vC= 1375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010011; // iC=-2093 
// vC = 14'b0000011000111100; // vC= 1596 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011000; // iC=-1832 
// vC = 14'b0000010110101110; // vC= 1454 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011101; // iC=-1891 
// vC = 14'b0000010101100111; // vC= 1383 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010110; // iC=-1962 
// vC = 14'b0000011000100011; // vC= 1571 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000010101100101; // vC= 1381 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101111; // iC=-1937 
// vC = 14'b0000010011100110; // vC= 1254 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111011; // iC=-1797 
// vC = 14'b0000010101001111; // vC= 1359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100011; // iC=-1949 
// vC = 14'b0000010111011111; // vC= 1503 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100000; // iC=-2016 
// vC = 14'b0000010100110010; // vC= 1330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000011; // iC=-1853 
// vC = 14'b0000010100100001; // vC= 1313 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000010011111100; // vC= 1276 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000010101101101; // vC= 1389 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111110; // iC=-1922 
// vC = 14'b0000010111011110; // vC= 1502 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110000; // iC=-2064 
// vC = 14'b0000010011111100; // vC= 1276 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111110; // iC=-1986 
// vC = 14'b0000010010100010; // vC= 1186 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011110; // iC=-2082 
// vC = 14'b0000010010101011; // vC= 1195 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011110; // iC=-1890 
// vC = 14'b0000010111000001; // vC= 1473 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011000; // iC=-2152 
// vC = 14'b0000010100110110; // vC= 1334 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011000; // iC=-2152 
// vC = 14'b0000010110010110; // vC= 1430 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001001; // iC=-2039 
// vC = 14'b0000010011100010; // vC= 1250 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b0000010001101100; // vC= 1132 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000101; // iC=-2171 
// vC = 14'b0000010100010011; // vC= 1299 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110101; // iC=-2123 
// vC = 14'b0000010010011011; // vC= 1179 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101011; // iC=-2069 
// vC = 14'b0000010100000010; // vC= 1282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111001; // iC=-2055 
// vC = 14'b0000010100101110; // vC= 1326 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110010; // iC=-2062 
// vC = 14'b0000010001110110; // vC= 1142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b0000010010010001; // vC= 1169 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b0000010011111110; // vC= 1278 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001001; // iC=-2167 
// vC = 14'b0000010000110100; // vC= 1076 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111000; // iC=-1928 
// vC = 14'b0000010011010010; // vC= 1234 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010101101; // iC=-1875 
// vC = 14'b0000010011001001; // vC= 1225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101100; // iC=-2132 
// vC = 14'b0000010000100010; // vC= 1058 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100010; // iC=-2142 
// vC = 14'b0000010000110010; // vC= 1074 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010111; // iC=-2089 
// vC = 14'b0000010010111011; // vC= 1211 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111001; // iC=-1927 
// vC = 14'b0000010000100101; // vC= 1061 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001110; // iC=-2162 
// vC = 14'b0000010011111001; // vC= 1273 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111111; // iC=-2177 
// vC = 14'b0000010011000000; // vC= 1216 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b0000010001101111; // vC= 1135 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010111; // iC=-2025 
// vC = 14'b0000010011100001; // vC= 1249 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010101; // iC=-2091 
// vC = 14'b0000010010000110; // vC= 1158 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011100; // iC=-2084 
// vC = 14'b0000010001011010; // vC= 1114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000010010000000; // vC= 1152 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000011; // iC=-2109 
// vC = 14'b0000010011010000; // vC= 1232 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011011; // iC=-2213 
// vC = 14'b0000001110011001; // vC=  921 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000101; // iC=-2107 
// vC = 14'b0000010000101100; // vC= 1068 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010000; // iC=-2160 
// vC = 14'b0000010000000101; // vC= 1029 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011000; // iC=-1960 
// vC = 14'b0000010010100101; // vC= 1189 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111010; // iC=-1990 
// vC = 14'b0000001111100110; // vC=  998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011000; // iC=-2024 
// vC = 14'b0000001111010100; // vC=  980 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b0000001111011000; // vC=  984 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011010; // iC=-2022 
// vC = 14'b0000010000101110; // vC= 1070 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101010; // iC=-2134 
// vC = 14'b0000010001010001; // vC= 1105 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000010000110110; // vC= 1078 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b0000001110000101; // vC=  901 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100111; // iC=-1945 
// vC = 14'b0000001111010110; // vC=  982 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b0000001111100001; // vC=  993 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b0000001101110001; // vC=  881 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b0000001100100110; // vC=  806 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111001; // iC=-2183 
// vC = 14'b0000001110110010; // vC=  946 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111100; // iC=-2052 
// vC = 14'b0000001100011001; // vC=  793 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011100; // iC=-2148 
// vC = 14'b0000010000100101; // vC= 1061 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100011; // iC=-1949 
// vC = 14'b0000001101100110; // vC=  870 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110110; // iC=-2122 
// vC = 14'b0000001111100001; // vC=  993 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011000; // iC=-2216 
// vC = 14'b0000001110111100; // vC=  956 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111010; // iC=-1926 
// vC = 14'b0000001011011100; // vC=  732 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100110; // iC=-2138 
// vC = 14'b0000001101110110; // vC=  886 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101011; // iC=-1941 
// vC = 14'b0000001101000000; // vC=  832 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010111; // iC=-2089 
// vC = 14'b0000001101001110; // vC=  846 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100111011; // iC=-2245 
// vC = 14'b0000001011111100; // vC=  764 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b0000001011101010; // vC=  746 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000001; // iC=-2111 
// vC = 14'b0000001110010101; // vC=  917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b0000001100001101; // vC=  781 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001010; // iC=-2166 
// vC = 14'b0000001011110110; // vC=  758 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001010; // iC=-2102 
// vC = 14'b0000001101110010; // vC=  882 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b0000001101001010; // vC=  842 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011011; // iC=-2149 
// vC = 14'b0000001101010000; // vC=  848 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001010; // iC=-2166 
// vC = 14'b0000001101000000; // vC=  832 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000001110010111; // vC=  919 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101101; // iC=-2259 
// vC = 14'b0000001100110100; // vC=  820 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101001; // iC=-1943 
// vC = 14'b0000001010001110; // vC=  654 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110100; // iC=-2188 
// vC = 14'b0000001101101100; // vC=  876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000100; // iC=-2236 
// vC = 14'b0000001011110101; // vC=  757 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101111; // iC=-2193 
// vC = 14'b0000001100100011; // vC=  803 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b0000001000101001; // vC=  553 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000001101001100; // vC=  844 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b0000001100111000; // vC=  824 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011110; // iC=-2018 
// vC = 14'b0000001011111000; // vC=  760 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111000; // iC=-2184 
// vC = 14'b0000001011011001; // vC=  729 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001011; // iC=-2037 
// vC = 14'b0000001010000110; // vC=  646 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110010; // iC=-2254 
// vC = 14'b0000001010101001; // vC=  681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000111; // iC=-2105 
// vC = 14'b0000001100000001; // vC=  769 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000001111; // iC=-2033 
// vC = 14'b0000001100000010; // vC=  770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101111101; // iC=-2179 
// vC = 14'b0000001011110111; // vC=  759 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110100; // iC=-2252 
// vC = 14'b0000001000000100; // vC=  516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011000; // iC=-2216 
// vC = 14'b0000001010001010; // vC=  650 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001001; // iC=-1975 
// vC = 14'b0000001001011101; // vC=  605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b0000001000000100; // vC=  516 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110101; // iC=-2187 
// vC = 14'b0000000110111001; // vC=  441 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100110011; // iC=-2253 
// vC = 14'b0000000111110011; // vC=  499 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110101; // iC=-2123 
// vC = 14'b0000000111101111; // vC=  495 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010011; // iC=-1965 
// vC = 14'b0000001000000111; // vC=  519 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b0000000110001000; // vC=  392 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001001; // iC=-2167 
// vC = 14'b0000001001100101; // vC=  613 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110101; // iC=-2059 
// vC = 14'b0000001010011111; // vC=  671 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000000; // iC=-2176 
// vC = 14'b0000001000110110; // vC=  566 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101000; // iC=-2072 
// vC = 14'b0000000110100011; // vC=  419 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000000; // iC=-2112 
// vC = 14'b0000000110100010; // vC=  418 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100100; // iC=-2076 
// vC = 14'b0000000110101011; // vC=  427 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000000111111101; // vC=  509 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000101; // iC=-2043 
// vC = 14'b0000000110001011; // vC=  395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100001; // iC=-2015 
// vC = 14'b0000000101111110; // vC=  382 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010010; // iC=-2094 
// vC = 14'b0000000110001011; // vC=  395 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b0000001001010000; // vC=  592 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100100; // iC=-1948 
// vC = 14'b0000001000001011; // vC=  523 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000100; // iC=-2172 
// vC = 14'b0000000111101101; // vC=  493 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110001; // iC=-2063 
// vC = 14'b0000000110100010; // vC=  418 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011100101010; // iC=-2262 
// vC = 14'b0000000011111011; // vC=  251 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000111; // iC=-2233 
// vC = 14'b0000001000001110; // vC=  526 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100110; // iC=-1946 
// vC = 14'b0000000110100100; // vC=  420 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b0000000110101000; // vC=  424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101011; // iC=-2197 
// vC = 14'b0000000110011010; // vC=  410 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000000; // iC=-2048 
// vC = 14'b0000000100111101; // vC=  317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b0000000101100111; // vC=  359 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100010; // iC=-2206 
// vC = 14'b0000000110101001; // vC=  425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001110; // iC=-1970 
// vC = 14'b0000000101011111; // vC=  351 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000000; // iC=-2240 
// vC = 14'b0000000011110001; // vC=  241 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100000; // iC=-1952 
// vC = 14'b0000000111001111; // vC=  463 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010001; // iC=-1967 
// vC = 14'b0000000010010010; // vC=  146 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100001; // iC=-2079 
// vC = 14'b0000000101011100; // vC=  348 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100101; // iC=-2139 
// vC = 14'b0000000100011110; // vC=  286 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100110; // iC=-2202 
// vC = 14'b0000000011011000; // vC=  216 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b0000000011001010; // vC=  202 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101101000; // iC=-2200 
// vC = 14'b0000000101101110; // vC=  366 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100100; // iC=-2140 
// vC = 14'b0000000010101100; // vC=  172 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010100; // iC=-2156 
// vC = 14'b0000000101001000; // vC=  328 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100010; // iC=-1950 
// vC = 14'b0000000001011011; // vC=   91 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110000; // iC=-2192 
// vC = 14'b0000000010100011; // vC=  163 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b0000000011001101; // vC=  205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010101; // iC=-2219 
// vC = 14'b0000000011111000; // vC=  248 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111101; // iC=-1987 
// vC = 14'b0000000010101010; // vC=  170 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000100; // iC=-2108 
// vC = 14'b0000000001011101; // vC=   93 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111000111; // iC=-2105 
// vC = 14'b0000000001000110; // vC=   70 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b0000000011001011; // vC=  203 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011101; // iC=-1955 
// vC = 14'b0000000000010010; // vC=   18 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111100000; // iC=-2080 
// vC = 14'b0000000001101101; // vC=  109 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101001; // iC=-2135 
// vC = 14'b0000000011111111; // vC=  255 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101011001; // iC=-2215 
// vC = 14'b0000000010000011; // vC=  131 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000000100000111; // vC=  263 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101000100; // iC=-2236 
// vC = 14'b0000000010011011; // vC=  155 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111111; // iC=-2113 
// vC = 14'b0000000001011110; // vC=   94 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b0000000011110110; // vC=  246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100100; // iC=-2204 
// vC = 14'b0000000011101100; // vC=  236 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101001101; // iC=-2227 
// vC = 14'b1111111110111110; // vC=  -66 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111100; // iC=-1988 
// vC = 14'b0000000001000101; // vC=   69 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001010101; // iC=-1963 
// vC = 14'b0000000010001110; // vC=  142 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001100; // iC=-2100 
// vC = 14'b1111111110111101; // vC=  -67 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010001; // iC=-2159 
// vC = 14'b0000000001000101; // vC=   69 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110101; // iC=-1995 
// vC = 14'b1111111110100110; // vC=  -90 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000010; // iC=-1982 
// vC = 14'b0000000000001111; // vC=   15 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101010000; // iC=-2224 
// vC = 14'b1111111111111100; // vC=   -4 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001011; // iC=-1909 
// vC = 14'b1111111101100100; // vC= -156 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110011; // iC=-1997 
// vC = 14'b0000000000110110; // vC=   54 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011101; // iC=-2083 
// vC = 14'b0000000001110010; // vC=  114 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001000; // iC=-1912 
// vC = 14'b1111111101100011; // vC= -157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100000; // iC=-2144 
// vC = 14'b1111111110101000; // vC=  -88 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011011; // iC=-2085 
// vC = 14'b1111111110100101; // vC=  -91 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001000; // iC=-2168 
// vC = 14'b1111111110100010; // vC=  -94 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000100; // iC=-2044 
// vC = 14'b0000000001000110; // vC=   70 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101110011; // iC=-2189 
// vC = 14'b1111111100100001; // vC= -223 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110101101; // iC=-2131 
// vC = 14'b1111111101010101; // vC= -171 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001011; // iC=-2101 
// vC = 14'b1111111110101010; // vC=  -86 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001000; // iC=-2104 
// vC = 14'b1111111111011100; // vC=  -36 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110011; // iC=-2061 
// vC = 14'b1111111100111010; // vC= -198 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101110; // iC=-2002 
// vC = 14'b1111111100110101; // vC= -203 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011101100011; // iC=-2205 
// vC = 14'b1111111100001010; // vC= -246 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000110100; // iC=-1996 
// vC = 14'b1111111110111000; // vC=  -72 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001101; // iC=-1971 
// vC = 14'b0000000000010001; // vC=   17 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110111; // iC=-1929 
// vC = 14'b1111111101001110; // vC= -178 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b1111111110001101; // vC= -115 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111111; // iC=-2113 
// vC = 14'b1111111101101101; // vC= -147 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b1111111100111000; // vC= -200 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010010010; // iC=-1902 
// vC = 14'b1111111110010110; // vC= -106 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110010; // iC=-2126 
// vC = 14'b1111111110101101; // vC=  -83 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101000; // iC=-1944 
// vC = 14'b1111111011001101; // vC= -307 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110111110; // iC=-2114 
// vC = 14'b1111111101011111; // vC= -161 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100111; // iC=-1881 
// vC = 14'b1111111101000111; // vC= -185 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000100; // iC=-2172 
// vC = 14'b1111111101011101; // vC= -163 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100100; // iC=-1948 
// vC = 14'b1111111100000000; // vC= -256 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b1111111101100011; // vC= -157 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110011000; // iC=-2152 
// vC = 14'b1111111001101011; // vC= -405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110000011; // iC=-2173 
// vC = 14'b1111111101010000; // vC= -176 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001001; // iC=-2167 
// vC = 14'b1111111010011000; // vC= -360 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110001110; // iC=-2162 
// vC = 14'b1111111001011100; // vC= -420 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111101111; // iC=-2065 
// vC = 14'b1111111010111110; // vC= -322 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110100101; // iC=-2139 
// vC = 14'b1111111100101111; // vC= -209 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111001111; // iC=-2097 
// vC = 14'b1111111011101110; // vC= -274 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110010100; // iC=-2156 
// vC = 14'b1111111100011111; // vC= -225 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111011; // iC=-1925 
// vC = 14'b1111111000101000; // vC= -472 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010000; // iC=-1840 
// vC = 14'b1111111001010010; // vC= -430 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b1111111011101000; // vC= -280 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100011; // iC=-2013 
// vC = 14'b1111111001100010; // vC= -414 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b1111110111111010; // vC= -518 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011001101; // iC=-1843 
// vC = 14'b1111111001110001; // vC= -399 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000011100; // iC=-2020 
// vC = 14'b1111111000011101; // vC= -483 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111001; // iC=-1863 
// vC = 14'b1111111100100101; // vC= -219 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111010; // iC=-2054 
// vC = 14'b1111111000101100; // vC= -468 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001010; // iC=-1974 
// vC = 14'b1111110111101001; // vC= -535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110111; // iC=-2057 
// vC = 14'b1111111100000100; // vC= -252 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011110110000; // iC=-2128 
// vC = 14'b1111110111101011; // vC= -533 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111101; // iC=-2051 
// vC = 14'b1111111000100100; // vC= -476 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100011; // iC=-1885 
// vC = 14'b1111111010110110; // vC= -330 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b1111110110101110; // vC= -594 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001000; // iC=-1976 
// vC = 14'b1111111010010101; // vC= -363 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111010001; // iC=-2095 
// vC = 14'b1111110111001000; // vC= -568 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111111011; // iC=-2053 
// vC = 14'b1111111000110011; // vC= -461 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111110000; // iC=-2064 
// vC = 14'b1111111011000110; // vC= -314 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000010; // iC=-2046 
// vC = 14'b1111111001001000; // vC= -440 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b1111111001011100; // vC= -420 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110000; // iC=-1936 
// vC = 14'b1111111000110111; // vC= -457 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111100; // iC=-1860 
// vC = 14'b1111111001110110; // vC= -394 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001011011; // iC=-1957 
// vC = 14'b1111110101011101; // vC= -675 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011110000; // iC=-1808 
// vC = 14'b1111111000000010; // vC= -510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000000; // iC=-1792 
// vC = 14'b1111111010001001; // vC= -375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011011100; // iC=-1828 
// vC = 14'b1111111001101010; // vC= -406 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010100000; // iC=-1888 
// vC = 14'b1111110111000001; // vC= -575 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110101; // iC=-1867 
// vC = 14'b1111111001101011; // vC= -405 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111011111011010; // iC=-2086 
// vC = 14'b1111111000101001; // vC= -471 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101011; // iC=-1813 
// vC = 14'b1111110110101001; // vC= -599 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010110; // iC=-1834 
// vC = 14'b1111110101001101; // vC= -691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101111; // iC=-1937 
// vC = 14'b1111111000010010; // vC= -494 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b1111110100011100; // vC= -740 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000111; // iC=-1977 
// vC = 14'b1111111000000010; // vC= -510 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b1111110101101101; // vC= -659 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100110; // iC=-2010 
// vC = 14'b1111110110101101; // vC= -595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010001001; // iC=-1911 
// vC = 14'b1111110101010111; // vC= -681 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b1111110100111011; // vC= -709 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010111000; // iC=-1864 
// vC = 14'b1111110100100000; // vC= -736 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010011; // iC=-2029 
// vC = 14'b1111110011100110; // vC= -794 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000110; // iC=-1914 
// vC = 14'b1111110011101000; // vC= -792 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000010010; // iC=-2030 
// vC = 14'b1111110011111101; // vC= -771 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000000111; // iC=-2041 
// vC = 14'b1111110101000010; // vC= -702 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101110; // iC=-1810 
// vC = 14'b1111110011111110; // vC= -770 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001111100; // iC=-1924 
// vC = 14'b1111110111000010; // vC= -574 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000100100; // iC=-2012 
// vC = 14'b1111110101101111; // vC= -657 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100000; // iC=-1824 
// vC = 14'b1111110100000101; // vC= -763 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011100101; // iC=-1819 
// vC = 14'b1111110110101011; // vC= -597 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110110; // iC=-1866 
// vC = 14'b1111110010010000; // vC= -880 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010011011; // iC=-1893 
// vC = 14'b1111110110110111; // vC= -585 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011111; // iC=-1761 
// vC = 14'b1111110010011111; // vC= -865 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001001111; // iC=-1969 
// vC = 14'b1111110100001011; // vC= -757 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001000000; // iC=-1984 
// vC = 14'b1111110011111111; // vC= -769 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000111000; // iC=-1992 
// vC = 14'b1111110101010100; // vC= -684 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011010010; // iC=-1838 
// vC = 14'b1111110100101011; // vC= -725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100000101011; // iC=-2005 
// vC = 14'b1111110001101010; // vC= -918 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100011011; // iC=-1765 
// vC = 14'b1111110010011001; // vC= -871 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101100; // iC=-1940 
// vC = 14'b1111110010111111; // vC= -833 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100101100; // iC=-1748 
// vC = 14'b1111110010010100; // vC= -876 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100001000; // iC=-1784 
// vC = 14'b1111110001101011; // vC= -917 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010000011; // iC=-1917 
// vC = 14'b1111110101100100; // vC= -668 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100010110100; // iC=-1868 
// vC = 14'b1111110011000111; // vC= -825 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010001; // iC=-1711 
// vC = 14'b1111110101001100; // vC= -692 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100100; // iC=-1692 
// vC = 14'b1111110100111001; // vC= -711 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110011; // iC=-1933 
// vC = 14'b1111110100101011; // vC= -725 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001101110; // iC=-1938 
// vC = 14'b1111110011110111; // vC= -777 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110000; // iC=-1680 
// vC = 14'b1111110001011011; // vC= -933 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001100001; // iC=-1951 
// vC = 14'b1111110010100000; // vC= -864 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110110; // iC=-1738 
// vC = 14'b1111110000011010; // vC= -998 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110001110; // iC=-1650 
// vC = 14'b1111110010101011; // vC= -853 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101010100; // iC=-1708 
// vC = 14'b1111110011111101; // vC= -771 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100100; // iC=-1692 
// vC = 14'b1111110011100001; // vC= -799 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100100; // iC=-1756 
// vC = 14'b1111110010111010; // vC= -838 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100001110101; // iC=-1931 
// vC = 14'b1111110010101101; // vC= -851 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111110; // iC=-1730 
// vC = 14'b1111110001011000; // vC= -936 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011000011; // iC=-1853 
// vC = 14'b1111110001101111; // vC= -913 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101100; // iC=-1620 
// vC = 14'b1111110001000011; // vC= -957 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101111; // iC=-1681 
// vC = 14'b1111101111111101; // vC=-1027 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001111; // iC=-1713 
// vC = 14'b1111110011100011; // vC= -797 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100110000; // iC=-1744 
// vC = 14'b1111110000001001; // vC=-1015 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111101; // iC=-1795 
// vC = 14'b1111110000101011; // vC= -981 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100000; // iC=-1696 
// vC = 14'b1111101111110001; // vC=-1039 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100111; // iC=-1625 
// vC = 14'b1111110001010010; // vC= -942 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000001; // iC=-1727 
// vC = 14'b1111110000000110; // vC=-1018 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101001; // iC=-1687 
// vC = 14'b1111110001100011; // vC= -925 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101001; // iC=-1623 
// vC = 14'b1111110001000101; // vC= -955 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111110; // iC=-1602 
// vC = 14'b1111110000101010; // vC= -982 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101100111; // iC=-1689 
// vC = 14'b1111101101100100; // vC=-1180 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101001; // iC=-1687 
// vC = 14'b1111110001001101; // vC= -947 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011001; // iC=-1703 
// vC = 14'b1111101110011011; // vC=-1125 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010010; // iC=-1774 
// vC = 14'b1111110001001000; // vC= -952 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111100; // iC=-1668 
// vC = 14'b1111110000011111; // vC= -993 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110110; // iC=-1674 
// vC = 14'b1111110001100101; // vC= -923 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011101110; // iC=-1810 
// vC = 14'b1111101111001101; // vC=-1075 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111111; // iC=-1793 
// vC = 14'b1111101110011010; // vC=-1126 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100010101; // iC=-1771 
// vC = 14'b1111101111001110; // vC=-1074 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100100101; // iC=-1755 
// vC = 14'b1111110000000001; // vC=-1023 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101111; // iC=-1617 
// vC = 14'b1111101110100111; // vC=-1113 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101110110; // iC=-1674 
// vC = 14'b1111101101100010; // vC=-1182 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010100; // iC=-1580 
// vC = 14'b1111101101110111; // vC=-1161 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100000011; // iC=-1789 
// vC = 14'b1111101101011010; // vC=-1190 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111010001; // iC=-1583 
// vC = 14'b1111101101100010; // vC=-1182 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010001; // iC=-1647 
// vC = 14'b1111101100001101; // vC=-1267 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100011111101; // iC=-1795 
// vC = 14'b1111101111100000; // vC=-1056 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101101010; // iC=-1686 
// vC = 14'b1111101110010111; // vC=-1129 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101000001; // iC=-1727 
// vC = 14'b1111101100100100; // vC=-1244 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111101; // iC=-1667 
// vC = 14'b1111101111100110; // vC=-1050 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101001010; // iC=-1718 
// vC = 14'b1111101110010001; // vC=-1135 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111000; // iC=-1608 
// vC = 14'b1111101011111001; // vC=-1287 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010011; // iC=-1645 
// vC = 14'b1111101011111110; // vC=-1282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110000100; // iC=-1660 
// vC = 14'b1111101111101001; // vC=-1047 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100100111101; // iC=-1731 
// vC = 14'b1111101110011000; // vC=-1128 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001001; // iC=-1463 
// vC = 14'b1111101011000101; // vC=-1339 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001111; // iC=-1457 
// vC = 14'b1111101011000101; // vC=-1339 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110100111; // iC=-1625 
// vC = 14'b1111101101011100; // vC=-1188 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010101; // iC=-1451 
// vC = 14'b1111101011101010; // vC=-1302 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011110; // iC=-1698 
// vC = 14'b1111101011111110; // vC=-1282 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111100001; // iC=-1567 
// vC = 14'b1111101100010101; // vC=-1259 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110110011; // iC=-1613 
// vC = 14'b1111101100001111; // vC=-1265 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000000; // iC=-1472 
// vC = 14'b1111101101111111; // vC=-1153 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101101; // iC=-1427 
// vC = 14'b1111101011010111; // vC=-1321 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101011011; // iC=-1701 
// vC = 14'b1111101011011011; // vC=-1317 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110010001; // iC=-1647 
// vC = 14'b1111101011100001; // vC=-1311 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100111; // iC=-1497 
// vC = 14'b1111101010011011; // vC=-1381 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010011; // iC=-1453 
// vC = 14'b1111101100101101; // vC=-1235 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010010010; // iC=-1390 
// vC = 14'b1111101110100010; // vC=-1118 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111011; // iC=-1477 
// vC = 14'b1111101110011101; // vC=-1123 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111011; // iC=-1669 
// vC = 14'b1111101100110001; // vC=-1231 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001110010; // iC=-1422 
// vC = 14'b1111101001111011; // vC=-1413 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001001; // iC=-1591 
// vC = 14'b1111101101010111; // vC=-1193 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110111111; // iC=-1601 
// vC = 14'b1111101101001011; // vC=-1205 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100110101001; // iC=-1623 
// vC = 14'b1111101010100111; // vC=-1369 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111001; // iC=-1671 
// vC = 14'b1111101100111010; // vC=-1222 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100101111000; // iC=-1672 
// vC = 14'b1111101101100001; // vC=-1183 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100100; // iC=-1500 
// vC = 14'b1111101010001000; // vC=-1400 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010111011; // iC=-1349 
// vC = 14'b1111101001100101; // vC=-1435 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001100; // iC=-1588 
// vC = 14'b1111101100101100; // vC=-1236 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100011; // iC=-1437 
// vC = 14'b1111101000100111; // vC=-1497 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100101; // iC=-1371 
// vC = 14'b1111101011011101; // vC=-1315 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000101010; // iC=-1494 
// vC = 14'b1111101011111000; // vC=-1288 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001001; // iC=-1591 
// vC = 14'b1111101010111101; // vC=-1347 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111001001; // iC=-1591 
// vC = 14'b1111101000000010; // vC=-1534 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111000; // iC=-1480 
// vC = 14'b1111101100101010; // vC=-1238 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000111; // iC=-1465 
// vC = 14'b1111101001101010; // vC=-1430 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000100000; // iC=-1504 
// vC = 14'b1111101011000010; // vC=-1342 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101010; // iC=-1366 
// vC = 14'b1111101011010000; // vC=-1328 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100011; // iC=-1373 
// vC = 14'b1111101011111100; // vC=-1284 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111100111101110; // iC=-1554 
// vC = 14'b1111101100000001; // vC=-1279 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100001; // iC=-1311 
// vC = 14'b1111101011000100; // vC=-1340 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100000010; // iC=-1278 
// vC = 14'b1111101000100110; // vC=-1498 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010010; // iC=-1454 
// vC = 14'b1111100111000101; // vC=-1595 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001010; // iC=-1462 
// vC = 14'b1111101010100001; // vC=-1375 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100010; // iC=-1310 
// vC = 14'b1111101000100011; // vC=-1501 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001001011; // iC=-1461 
// vC = 14'b1111100111110010; // vC=-1550 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101000111101; // iC=-1475 
// vC = 14'b1111101000011111; // vC=-1505 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010100; // iC=-1452 
// vC = 14'b1111100111111010; // vC=-1542 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011000; // iC=-1448 
// vC = 14'b1111101000111101; // vC=-1475 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001000110; // iC=-1466 
// vC = 14'b1111101011001111; // vC=-1329 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011010101; // iC=-1323 
// vC = 14'b1111101011001101; // vC=-1331 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001111011; // iC=-1413 
// vC = 14'b1111100110110100; // vC=-1612 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101100; // iC=-1428 
// vC = 14'b1111100110100110; // vC=-1626 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010000011; // iC=-1405 
// vC = 14'b1111101001010001; // vC=-1455 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001100010; // iC=-1438 
// vC = 14'b1111100110111011; // vC=-1605 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001011000; // iC=-1448 
// vC = 14'b1111101001110000; // vC=-1424 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101111; // iC=-1425 
// vC = 14'b1111101000010110; // vC=-1514 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011100010; // iC=-1310 
// vC = 14'b1111101010100000; // vC=-1376 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101011000; // iC=-1192 
// vC = 14'b1111100111101101; // vC=-1555 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101001100; // iC=-1204 
// vC = 14'b1111101001101110; // vC=-1426 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010001101; // iC=-1395 
// vC = 14'b1111100101100111; // vC=-1689 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001101001; // iC=-1431 
// vC = 14'b1111101000000001; // vC=-1535 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101101110111; // iC=-1161 
// vC = 14'b1111100110010001; // vC=-1647 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101001010100; // iC=-1452 
// vC = 14'b1111101001101010; // vC=-1430 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010100000; // iC=-1376 
// vC = 14'b1111101001101111; // vC=-1425 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011001101; // iC=-1331 
// vC = 14'b1111100101100101; // vC=-1691 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101010101001; // iC=-1367 
// vC = 14'b1111100111110100; // vC=-1548 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011011111; // iC=-1313 
// vC = 14'b1111100111101011; // vC=-1557 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101011110101; // iC=-1291 
// vC = 14'b1111101000101111; // vC=-1489 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;
// clk_100M = 1'b1;
// iC = 14'b1111101100110000; // iC=-1232 
// vC = 14'b1111100111101101; // vC=-1555 
// sigma = 2'b11; // sigma=11 
// #5;
// clk_100M = 1'b0;
// #5;




// end





endmodule