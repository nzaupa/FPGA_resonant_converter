��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C���TWNĆ9�_��4[���~��E����B
2�\���.�}��]`�3.H|/�����H�1�@Jg]�2��U�;��X:�4A.�z�F5]�ox��1�^��Pi��I�~�V�I��}a�m���v�4��⒀M
rzx�Of]�Ц~QEX�N�d����f�*қ�J�)U�G��/��:6���"qc3YԨ�S7]�L��k�� ��Sf�'}󲶥x���5Y�ߗ�Xtx���i��q��j���2�B�1�=ѹ�������-p�^~�m&�X
"U!��Q:��'�����oDp�����R R�L������o}������Z�Y\�F
�芍�gE�K4J8�Ѓ�\��}�ʮ�e�g;������R��*�VL�/^��^it?�Ʊ��!���؊�fȰ%�?��ʐ��}��T������3�n�)
1�����}_��MG|�@X��.��t�H�~^�
�T|�H��qݳap�?G��L�qØ"��?���5�53[����.֬C�uxW���Uh���=��b�0�+p�"�x5B��iiW4�O�]x��H��p��Lp�7���^��/�om�%�ȟ��͚����)��s�LyM��D~�l�f�� F"���٦���o�7�<=r/"?�a���n��#z�-��8�Xo jiY5	��- �rx�(�ұ�gо]�c@����Ll��h�NbxG�b�Ɔ��>O�H���s�ޚ[5��fx�z{�OT��EL1�j�X<#�P�T0��N�	:��H	c2o`����_��"<;C��Y�y� (E�_csL俉��j�:
V�P�wT���0�W �ve
�X:d[�s�@��k�Rnk��M>+`1.��O���:
`�����)YN��[c� ��_�Q0�����_~��-ɗxp������h�!v������<��F��~B�g��;{��_�~�5p�&��NPy��4i:1Z�S�Pi�����`�d��R�i�<]���5N�ߤ`�)�=�^����@] �p$L;©�_�?ڤ]�K]-���/���v2��ʽ󄇂qC3�{� �m2*��.֕Zց쯨�>���75A��Y�Q�գ�@zDߥx�O��P7�l/uu�^�$���u��Y蜎SY;�+��Ü<����e��D
k�q'Ѓ&Ҽx�(�u�4nrL:�V��J�g�-?�~	J��[)/��.:�Z�ԲX��/�Ȇ�KI(�뒐���b+o1�j�^�Ү1d�xA�u�HI@=�g^���"*O����-):��f�l{�b_�Rgd�٤z��3�*X[�WY���?�21t筡�ZoxΗ���N�A_�) �(!�U��!MpF�y���º���Gƥ�]�>��kb3�:�sV�a�_��d��&�vf��{�����y���pB��N�sF|����х6���B2F��7l���x�3��u%"�T�C+:���-t,^�� �c��a�̯�b�~��+�O`?2���73�X/=�،��Dt�ڥ�����OC�����ﻘ<��_�9e�m=lj�IM��ҷ<Si��~�м��ɬi�f�D;'C��7Φ�/����og9c,}���,=`� ��lN96��9�ЂwE�(�)Kb%/,U��9!9r݅잎�x�\���n���߃��S��-ڽ~��C	y!���_-� �/ዂ��B7x���Vdx���K��k��h���:M8���G�0��.�A4��T�2y�o��� ���rn���G'���I ���/����΅��%Pk��C��p9��O[� *\t��iF�6wIi� ��B��:�`�� ��'�:��n�:aCe�"��p1]c��IxW�}�����&���T�`+G�o���03��a�%(�#��.�>l3��B4C=�$f��~q�<=���N5�!/��Z��֟��)�~�xP/J܍o2usT��}�,;�0ߡ8�����ρ�@AC*6.��ĉ�4Mhָ7%��i��A��q�F����ݎ���;��9Fq_7ш�Q^pU	�f1�����ؓV����t��6A����CA�vi2�[���{v�p�f���;�F�YK8H�;�A4P�� �����b��ܽ�7�S@�"�|�u���,�!���=���3(�e�`�C^��&��)���FO[P��y��B6��>�}Q�dK��(j���L�n��	A�/�L�՝L�a�W�j��5�m>�?��xh��6P���-mT�4�HxZ�P,���듯Ì�/m�(�J����ԆG��(��Bmd�K����F�mLU�}<���N�g��Gܡ'yDVk@Ӑ��%�,�f�+��1��QH���(���^3�z��W�9���I�h�@��j{Qc����p5Kȇ�w�X�n������q�ؾ��'����1�@y	��u�7n��e��\,)�j�VN�Xӯ��A���եy�W7U�Ǿ��|c<ۇl��}�@LG �0Ej忞�X;u9�L����`�y�b��:��`v�.�H;op�nc0�<���X�)���B�58 �5O���~�Ljq����|osc{���;���<U\�����L�`���#32'w�(�ѱ������H�����J��BC�zI����
H�����puq	Uh4/Li�C3����⅘�����=�,��DiS�'RcD�ܶի"�����gVJ��
RӍ��R�$�g���a_��؏���^�\m��yc��>�b*A�-���*._u��6�8�x�q�/ꢁuF6��ɭ� ʨhm����yX���	����Y�
X g��J��')������T8ϝ���8��3|�3�S_�^�,���)�����e��L�Ez���z�^�i¹R�b����ܴ=�n2è���R��˒����K�<�G��0�������р�T�p�в&���^9��K�*���p}H1m߯��z�v����'����Hp�(X7�ԅ�n�&�a|H�i�1��u��p��h&F�S�ʏ74��s�h[8E>�ZI
N�|��*P2�������M��Փ���ߕ�B�����P7�� Rp1�gES6��R]�;&�`��r�b����C�-�������:��t�f��Ol�\����Ѝk��J֚Ȇ�&�B_p��r�7#�;:ܮM�8-4 �/���r�[vʗ��L��m�o5$],VI�o/�v�����@\Dd��M�eI�B���Z���޺��9)i[ǰ�FOW��=�Ю��T�a�~�t�����\�!��[����3���s~T���ZjA(.7U-��V��[*F�"s�K�ϲ,��/�A�� �8�%O����0g����I�����	B���[�!�?wL�fT]D�\�(C�](s�h����vt�>cV��0����Π�,Cm�s��D��#��T�N>�
�T�M�.��?h���2w��1��hE���!��ˉ����8��ya��1�ؒ9^�8�^k��TTB\�pÎ�l�k|9�u[�B#����RU!��0N��H@�l[�M��d="SE
�$�� a$x9���W���z  "��]�D�U3H����d��7~~��F���sV/��U�-%��ӕi������$�Bz>�b�}�_F���1/j4y6ㆰ�T��I&Q; %-Y��1�{1���/#ġ�\���Ќ��5G� ̗T��>Lj�h��`�������!ſ]k����a���5�;l��75��� �cr�o��
A�fޔ���{�Lx���J�q������<u�
�!��c�mU�Z��b��2��Q訟��p)gNx��n��F3Bp��R<����kx�>�Q�V���-p�h�ij�]�z@a�����C�R��� �<6�G\4�L��<�X�W�9���ol3��[/��+%r��ߝJ냡�f'�Ώn=2`�I�B��r�eke�'l�d���7��u��js��3�#�;��@O� ���=E�Pi�ϨMid�߽�Kw+�������I]wo�x��'i,��"0`t�Z������T!��D�9� ���D��T�+�٬&e./u��
s)�� �Hc`X�e��+��X��߈����%�]�L}DS
��Ƅ��|�5���P7I�a̹�y�5y}���$ܷ��U��!UO_��*��:����du�6ͣ��ѱq`�2B1!��[J7�)��wVr8$�p7�رp�3i%�K��%��P0��l�