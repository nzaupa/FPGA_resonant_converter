-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UnjORBdNah/1md4jgyELI6ubHmZIxmkWlxF7QzVFaM3qCc+PKjMY1Z0qK/dWQ9rmY6/vsdaXW95O
GrmtgjuWFir3Sz75Rvvwvg0pKkKqFQDMyzJ7ZI2AoELkeZ/uHL6WhgSJOaBRu+FkgGoscy53JRmh
Jaj0z5/oD7CIwUL7HAcDAYLuW3uHraz5qPipHvrsOHDSktWNQgATxE8acw0U2HhSr0eD45sj/24N
hYO8heh6CEa9srXyWhIDNhLqm1PpckSLraHqcJhgbhFiR6LGG6XwThR7i5kHG9GJLfGxzxhpjEvb
ZtQRUijWOauadkAYAMySq9opyePuk9XlN/vR0A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7296)
`protect data_block
yH9EqMyLITzYkPmNooH2ftR/9Vo/+mpmvPymU6ndvdFdJIFSTOfRNzL6Wf11So5/E2GkDsvZ4cXQ
Ng/Y1hZDdCmW6c/erRfrakgVnvtOCCK/pmuant2rOUK+7YxmD04w9FLWIzgAdDevh+xM9Kxs36Gt
MQSbgUQ7KhVbYAoZGa1zyKpignd7QIAvTpN5WvwONrYq4PkTPYcZViktZ/m2sEFf1dOvBqZPn9gB
qOoWOQn2u6xUiA8Boo7VSUcoasiX1nhfMsPS9xLb1J1bekdtPyMVAkzqc/4Gl72CBAar8gccNAjm
5h18mPwU+QeFTni/inU0qj7g0EjQp5aTx4UMY+qdPx9d0YzfQT7deWPDpjfmtXkGljLdTV48pTTk
Ma9qAJjDmReEydfr1dupqjsL/5aPLKHgON7/JPuIb6/21nKSrBxvT5UptfEPvZkzB//UlRqQ3Rn9
PXZ2jcjJsEYyriKZLGGKUqIBboEk8QULpPheKtLlG7/YAVWDI9qSn2CrTZQApIECZI85WNkQK2MN
rbOqZuLzDg4xLeVxfRryDDj0LA70nJl3FJzyi001bQ5SDlIbkNHwVgiVHBN1Vcq2sUokxwT9CAC6
FnsCNrG1ofdEGA4kuhXYV9AhvFt43PCWS6gLyhm/S46vbH2FxmIUF5KEmVL7KBeKDWjvMxLjnbdt
sxJlRpJSUoCV13CFgudIxzR+lmQ2rDAq0pkpVwswSrSkJq2Ovekaono6HvniKkgkbrug6eOrJoAN
kKNmpQLiepJJ2Qg+CIyBR67lGhuRRdZh9hh0XZTp2KJZgP5juhG6Xdb+9wPBsy36K1YMDAJPySoE
mjOHwE86A5vaH2IJynC44njjpfF7TvNA0LJg7cgUfPQdfNSkG6M+VvibHLQHHe041Zp8pf3gU+I3
ZZ64gekcvNPv94SqecxOW5b8tpXl1AqcPVgzN1nCWRYd7PovUwCpr/9B/tzzJ//PlBPvvUS/v5nZ
YpieqsoPrpVFRlgY1kGwwFp8dFCACj2F07553s0LbGnOcZ66srBmzTdLtYL2G7RsAnUckeA7xSNE
Kj2YwO/hAu5xCjpHlHO/zuD6A0MgOu/5tMXY8lGjf7klDRO6mMhz2sqhx/JVCxWwtmFMF+EX+11s
URMdCEkVFWeazjC2G2fZr9E4Zk2tgsxqCq97i7Dln8qhWbnrWkEEOeyqW13hKLr0WsBXZJkFw3Ve
4C19VW9u4C4kWECVj/hVI/9ppBCqLVWK7M8QJzaD/ZNQthmwrSxhSoNyM80NpdMlXkVdV0ne4cq2
CIvSKj85Vnn3lCOiyRaQNKMDOs5C/XETUvMPU0mRZCGrJYFBjTO1KFtWSHJlCY/39xL3cQ6qC4X0
yhZCw3KfASmDyBZBq0M0XUyDjeiF3rX6hQV2tjglprUJXLbeaBHU/9Qby+4S0c1saryc1ixcW8QS
gByP+TWHXN/CTb9TTfvnn328kDonHxZNT/Lo+1rHd1dGbSTEY8R0xVzeudSwK0pCcQ4m9WN7sAs3
ssXVfKdwUq0v4ZjbfMkrAq0E+agLMI/EjHRq+qvRwL5f1KnBSFMHzd+CNEtznuBNu2mz8a44oHYA
Zo9J8uFq63Mb7h6Z0vY/ZR7XjjBPosP2AjG/MtecM/dBbOzUSsWNtZR3oXgDQ49CneBlQhPKRYmp
ZBYjxwYLjl2cKo83Ut4tDnu//ABpXnutnlRLzXID758WRiPRnWM23LkRnBQKgn4giwezwlMEsIqM
zMys6oIqPBciUTH3wVdGlPKVjfYEAc534Fe1RNmSRxG+jWV+fXDB6jbGQ80ctx+5KOmslHvuE2xM
r9QvlSYnibUG9s5kJlOeArWWfbAIBkJdzh19o1bkm+8sQfOgs5oPf1xUqYgeXfNG4SgJHNHg+Tgy
nE1f5Y6POkEpU/iJLkTe1JqNnT5WyCxNyDVTwpe0KJYtwSRyDbb+yaoj/MPMZ8+8w9BTm9XavA+w
5fVKCFwqwGphJ3OZG7uocWcmoFEj/f/GR55c+bv8mbw7HgT9NxV1joYmaB3kiENCkS2fdpPqbYK+
gIs8zzIhX4QDl70SutP36mIBqR8JeRKB6sLiF9ccEmKvtBXc4mu7llPeepTulNaJw+Nh+sVn19R5
zgXtEtdmOaFTL+yKRNwZ+UscxnvjXcZKZF9JpQIi2VhwDHteVdco/cDouZjhoNOQ7w5pOBVxFPlp
jb9+1swrCH0kFZ06Bv2C8lhypMngoe+oJRPM7xQ4+E3OZP4ICaingHP4qorUXap44h5O+SlWTPXH
yYs6+yG2t0IpdDjMT0w2y/YTiOqNTwFmdzdp2J3cEa5e2JfmDZM+g4dpJBqBCLV3eHTao7YIU9vE
8aOUE8KzaMHRP0p2zvXLTAi6cNxmvxQX8r3YNKsZFauBKT/EXImHWOajiVi9o6zIzAROn56hZOBW
r3R+Uz9pxkblbj3eW4SOicpZmTJ6FBhci8XzDTU8Gt0K6vkMWeRhoL56NG6cin+U2YJBJQ3HaftG
qjUJeCOPIy/r6yqwzbARqy3ntKYZsZdCV1SG1ydD6c3p/kEqdAXwKf/4ArqmWuP7oIKbVHaDeYQh
FsPrlT0eC6Uq1Pi2QVKBxEmxX/j/Ecuwyr6F6BRVcIXm8oxHKZNlocjPkOjX2YrQyjciSMlfVC+V
+M57UdimHW0S8c63U+nrPwheJ997wmhM05O1xNjst2fpXxdV3gm82mGnpmLeB+RuRDQUAk3sMlv9
77tFGtDmwcVa2BJ1NNK71aCJ7pZm9C7Ks+yOMwfxNVEA+KEn0H7bT3gDQyMOAn8csyF6x1LkmKI0
vEb4ycm2wg1Ad7usDaDCRdceknOLBPTliVgpQ8HIwKCWHxVSLs/tgCTTXt8oZJlJskNJLD+ZFv+t
V6iScTT+dOx3Qvlx9hQRsWAv1iO1ni2eYhH6XZAQiuA/jRKcAzFZx1cMcyZPBJRS0yYz0XzjEM2Q
70NzYmuYCZawJwnaohrD4agRwq09XMP0J+dBpGqc56AuMz7a9mL8QeP5NWk5I4amz40bW4UR8zm1
05aOU2tKEPAMRm5G0QA5P+7KZh+Xr7qERI7TJZwGc7WrkgHvkv/OPSfrNEB9se6DrZxuYS0PHpF9
ncnXXe4e3uWMAP7cewJC9nN6XW8UNLApMG4rh+ugdBnClMhCgoh766N8UAuJMCQzLaaZxH7m6rS3
vVTeN/F2pHKLADUf8I/7/XgpkH/vu+0ZaK+GUZxd0JgtIllI+1Vu/lpOhMcSmMDLSrQw8P2b9BjD
VJOUApzgeI1Y7aHntA8XQ1DD+JHbEzS7mGuOJegef+gp7bDec9jnsTIKsFNdjg+nN7rN6sopcA63
0fYA9TmBMDMt0Dm889dQs9XuQnA4xw/3JSJ+8q8C7DhUi0kOKjJyT42kqq9wZoN/vtw9bJxcyc2q
aME3YQL2K4X9YUCTT68RD1kLJ67ysRCAfQmBpP+dTvIxFSiMXFL6Vod2XDh+mCgTzJmPRWWKpHUy
zI7ma/+o/8sjvP76RD+gRHOrbjEIg81dehb7zHMQsx52ueX4Jg5qolHlOIdKnaKNuMgVy87n9k6Q
TT/h4nVNx0/4ilmmUL8hv0qpWxJlfjCa+9kUFpKRYfzpBex4ISoOZcuXs9pvBVi0sfPdvM4grbEy
T3ZkQGcPMflejoV9pcdpjWcGn2b9Ne7Tp7jcxKTgEpGeTby3IpN6aRTgE7sb98qsrq7eRUgI1nfD
dkx+t3PO36LZOVcN19VC0UPwOMudS4s6YWPtG8TTji74o4T9DMMpDAXJcpAzIr175gULOs4AFfri
6jUWFK7Tf/lI8RP1OHbHgGhxI+ZwEr8ld4mppjlaPNoiWJDz8wqScdmdwrmQVI94ii3SexIhowWV
K+fiIh1XFKu/GUj1VO9ZOZl19rTXJEk8R2dzesUoEUX58JmO31HPozCIGAhTt21WOi/BFjUvswyM
OpsnzUjC8ATUwcY7KH7hS1TDpvapze4vv1ApUnpvZazjjh9T6qip5OZJUlK3Ayt9DAZDtFq0NEdy
Makxg4U7jLdWtnrL3cQfujr6NDDVJLWeiDoX0jESqYJQWqiVsMvxEuNp2apTx1Qvkwsji8yYazIx
CXkiGkc0GKH+2HsDUWPrR61nxF9jdq+kdYLhylO2P+2bgia79C41GAYf5tU/ZFWaJPh3uCXxrB0P
6XuYyfL7EvJ//DVJABJ6mveBHLQMtt5GiXfwyczbcviqKDKX577VnhNVgHBpWzdHnRQbPAvVX35e
lz93AxlairRRhz2HVA26RkegSrXKmapXyzFImB2xe1AQP+FTij9eiTsMMBFPP0LBgHJIf6wFYn8x
jOLzQg3a5j8OgNedEFiiwR9ViwdvKAxcTxY2QdaGAGiaPrR/VZzHEp2itABN5fkzWCyz5NHKUldA
vvQe7d8LSmK1TcqR7H0xgaAPwcX0y9bGMlggzyP1EeK3w6EH4F1KJtRH00ZXtB2RUxlg2JjDDMPm
IkmR4iXQdr2IkVCXgj/QbQHmxbyU3lG4C/dmkXns+8MrHdMTpHDJU3h/YBJSDQx0RZ3rZ8ZVlVFh
CS2apnQwbOj9mNrLs3p2hDcNvXyxFUksaYkUQkceNbwdDmU1QP2C3UzJ1ql4g7O7rr6H472CclTb
NqZ4DSVEfGgxGj8IMTzlHYw5OsKEjRM3qMWDsXDn8EQVt1pTaXSE1eNmwOe01v9Ad885oEziVHTL
uPvvsR1SVQ0x9Oc0T1t0Bue28Z7GVBHFKxplwQxnaTm1lTCIfOUpUve1KmbZFMSGUqu4mJQsrXFf
J0nt6+DRKG+Ly0/P7PheKq6ObuHe7cgw4PXXkTPNOki9gFnpO5GKBtMu3t5pNzhgXcw+EjosPd9h
i2b8u54B1ZjLMD9v5qNrWq/6cBd98k9xuo+cj3+Q633WkRszd1Lz/uw4ofBIqVIQd26iHlkhQfkt
/7XJx+K/rk/kYsdgC2KtNkU3rFRR9puWOxSypU6SzEo6MdVSf2KG/FM5qhjM2fuN7EltsnwkbPLQ
hIlgaLNU7zsuzZoeDkUbCLCALItkT6ArKu0NdpC69fIvL8mGuwAhSc/p40XtjnFDvStk5yKNONJh
RAsk7pz/bWSGVkTpiy5sgKvCldhoGhJFBR2zwlVQgaY0wdiNAosLIWNplIC67EFNrvHTxiNcX4Tq
KVgE+IlMPzcb8xnBDP9GRGUxbIGjyAnnHtNjCSPa1CnUiDoMfF9hOgAe8ax2HdOtOuc5klDvRo+t
EqgQU5351sp7QkigDFT+4tNscS59o7Fn5TcobtGSrHDxzHDs3GUCLptvddI82rfaKQS2Qpl/acGv
FgQ/pnaxCHQ0J2+9wVcHELWG/1+gnhnGCuhi37Wl4/je8dLjKZ5VMcCbqD5tdO0AS7zvkTA2ss5d
tb10l0H1XUbL6ljltoqSDsrJO5XuMfvnD21743flys+/NRtcTvFvH6GP/Uw+xFWop6NSxm50qDdT
+rRSiwLM0t6/erBNMOxxo/J5ZOEapHDZbFYR3VR3y3h1oAB1Sc6L119+R+OyM7C/Kus1W7f1XoLU
ohBHhKKh8fUJMa5A8pSwv4CgbxxoCtAEqml1h8WzrnaZksEgVrgaFgVQ1nf4/xXK4ushj6i0w+A1
tUE3/rneA4c5PISB99gwbgV+/MpdiYHmiqNscD7XX2QeBIV+6sOVZDv+D5J7D4oPA8EScojD9wnJ
MH9SdXsm8iPqMKqiM7wXM5GwsV3/vF9YWiBRtMpyEt5V2jtAzw6OB52+Op1AWhkmNYhqvPx+7uhl
925EGSOoBoUxtlj8rDtZBdLuXVvZ7K87vO+9Ubv2YwUtGZzZcqbKtoTJ/tX+0Hs3eHewTVK9YojS
bf37r/b1u6pTFHy7shFkyTk+DpmN2qAZU4pMpo+2WtecsPyc75vRSqPmmIoL+5WiUR1Ss0m5gg9B
W8zyFbFmkaiXCnlmRCmOEBaWXRRZLQ8U74QwhGattyxrucSYOlEq/mVWloM6SJDl3JJUoWthWSum
one3X6nqGfJlfZkdLhcc7vTnfaSt4U2UN74/sgI5JFfhyRKjGXbqfZB1N8ic1pF96re/70cKhu6Q
LGA0+GRa58PTw9RpW3BmJtVsNYpIq6KSaeaAKxptpOj3Hdeh40/BQGXEMPVie7mrS7GR+I1SmN2y
t/lSRULur9asE/4/fvD6zJY6YUPC9x0nRigyvvSIha+XbdR+86D9djqkWcPzTdX2+zqjCKOvFnqU
G3b3ggiJzYNYml40YjgaS0P3Kz3r3NKtTUsY6hOrgeO9q9CaDY8sluCxgKvHxJUcjfqI4Zx0qypq
+OMcx2IfastVEW2ndoEx8VMVDeqUbNmhpqlPsbQLfZ8srtnBhDXa5ZsdJDTgOoiGxDgiyIdhGIMz
94t3CnFYwoqKW9nDxYYSToHjb6VKUrofqtcKZuZ2F4sW1S7jE9KGFOQMfql7Ek6hVsGKTMp2x+/n
NIV8pJ6fucbRd0Y2AbkgLqTWPk/ufL8kCsT8ZAga12IizBRh3R/LIPqHRkdV4hXg2jZnUhx6a+12
yhIi7arGRaGM9oAkYdz6sbf83AMydUdOcDROb0Q5t+UW1k5wGCEtzMZikmZdA456rWjaFNT0/BI0
AVq4xdIHiieyUNn5nfdusaR/q5LLOe+AVjLgN1d3tzTomSaJsi/GlCm97F2HWeULc6Ky7Vx1/tEi
wseMyfOglsRiEJyfxECy6KMg3vR3beDKsHHy6fx399VrG2o0A0lg/thJTN9dkWb5cu6TCis7V12z
hgIOLPg+OxqVD929oh0wqCvuLPivbVki1Tcd8UVHKja0X8gfQq5psiWqWbEZXEIU+MGvdoJTq6R6
GBBm2lyg3cPJwz9umWuc0sl+8bsBAiCAp7rDQLBpB9PcQdL2NrRrPshujktrl1O7WE7EtPf3YOem
Q4GqlMANJ0cQ5PIK3oW//t8rtB0UNn1XAhwcS8c65tRKucnrIVvEBJJdlDWZ/8zLA6i9sWxqZdbE
mPawmZnHu0nWBjZch/B2uMnmOpl3nCfQPpUpOjdRC2WMg+F5cTyU0Tows8du2ik/HAVyQtBkRrcI
Oj1gV3RT0GrMx5kexKbt6KXJ1MKCLOcppcuuS5onnXOSmFZkLskrQRzbSTIwJDLRVXPd4llbPjTe
NzIpd9GzhgScgxnp/0UceVpMKL7eaCp8hWX1FmnyoiH7srA31PxOYTmuQe1SpEKKm0V4WnvR/lSS
8HtA1Vi8pVPKelI5KK2bVgcqC7Jl6agygAym0XHX+FxAC7HWtsFUlEtXFMvPJ8V2GowWhzF8fWpU
flLFL9Dy0hKP3576HGPNeZlrcivy7dqxhkm7/jOhej7fpyYhG/2Yfr6WLgUXOIkmycMka3j1jjpV
c5EHOhfamb4P8gKQtHqr0UdH9xwednO5NlnlwLtkz2m3ZneRZmWySyF/m+V51JCNKgZNcluMAKnw
CaUPqv8J/dLFd3xyficYtsEgftC/AhWAmnDeFQ4uF1STo2cJf4uRoySiWpVS76CAjBQL/9X8xZs/
G0IwUn7bLRn4xCR/zxVtfRdfSa2DpEd/7OqjFHNNE4XDb6Y9OqXOv5KQm+FxjWT/aS5meJNSdOei
/kPxjuE2PT5TrGxKPsJZPRoV3Xv5+ohFu4gyG6eyLGuV4pfrRF85LK8ythRQeD1LydGWl19laYgV
N5dNKLja5NGEJsICxOQRzRQfAnO8L8FRxAscXDNWludQrx214WAfOIY7lQ0ON4qpzsPoheq0/inr
M63veHnG0069GZXkRhEP9n0/GOc8Nh/UZBefB2slcKJqw4Si5uYSZYViFSbt4CnBCqqKaelZWcOU
yUdXzXXMWBXe6H2GAdO95GmEpsYu26cMab5CEzQu8q0EYfpYgxLUyu1tUsBoMIN04ZTncizYrNDx
ypKwtVyHPBC78Uvrbrgb+yXsnr0nX87xFXCU+/EYqBLWaIF5amksu3mc9YCUmU5kgAG7Vp4karFj
YTvomDR5S70cLcAVdTLfz8+q7Zl94ID2sc4CXpHyI4u0ZpiT7Zh0/SlYg+f0E9IMGNwROjvzBSoe
FcEvjUvqWMg2Rca8MybFESDD6ZT0w+Pd0PCBRZbB0U2stZrq/xrcx+ow5/6PA+s6n2Tl2seXddsY
m9zBli+CGpDLlRX2DuIG7AIowPeXn5Opt32gp0mcUOWt09EKr1A3pRiXYSravUnsmmIQIDWBInHz
M3VnX9DkLHkPkGSdOItH/IsV3qMMdjdpQ70CSgNiLlIhgyAtbuYWHTqKmK889TfdMyxPZkwbZdrt
wuiXX94EjRxdfLm6loU7ioXmRuuHGiqsOBDosmz2ZL3zO7FXk9Tf0YH8Uk20OuW/5qaDLbM2/RWQ
ipcHsoMNhilk1V/DfS0mSFiEDm3ArpS6UVUQ/nAXEblv2QiX0VpOFmsEXHfWn96JefPURl/ze7gR
SPZjnVy0GSj/76+Y43U6w81aCzdwEtcFfrPCwEvnZLmtUmPdX+2pPov5i0EyoVjNELQCHuqXzbfh
Ii2UD9OAkQNEgro1rb3CcNlVbbKE3YoOpav0TWNPGT00pAG7/t15M3LM/BGDZyo5OsPqckrHkDsc
SLu4sEBrqu73EDwxtgoeySR7TOYRZW9APN6uq4QPaAXfgnkS+34Oq0x130sgzXVs/SnFzBY33v72
S6AiOyM3B3e1jgtyOfBEJnAXr94P4ZHXaDeE2c30efTGwPm2ltgYcFteC7e7Ps0MD3xxs8ScBWbE
qUi0k+2Q7ePsyqzHHIREAQMNu2j93PF/nOHol6nQXS4DKNjKmndroWUtJCwVDhCyhaSVTStyJ73k
zhd3e7JPfdMKmxQerUdq2rT24WwDaKGDUoOhUo7IYlUMlJBiWWqd023LN4PEJVAG1K+iO5lXcblF
IUQDh7Ax9n3TbPAAo4jZBHAv8rXNfeoGaTdCUOkxZcWVaI4Yarp0+KuwcB51xcNdYPCXEkEZ6BSL
oVo1K+d+xxPio/LrsmtUxjZ2IfFfcXTt7/FLQBA9zikbFM/ixRH/iGIle26eP05oFeQ9YgXnkwg1
Xawg8utaT5xTrFdsyfUgIOPhker+MaXq+RIwbqbREhFNWiuQ+jSncrZ2IscS47rHiJMe4oeirBLm
t8ICpJhxThPfFmQVOg5TsbOv2TmpWGt7jVUMg5dEA7WZozY+Zmm1ZtDKjg68Is3yoJBKWIwFG0Dm
LjzzsCzOckCERsQMbK1n95BXcKbkYfYehkelsiPxP7zfXAme15cG99qBSe2PU6ELNL8kefgZfZZB
SFSqSAVul1c+ZVkCxLC6FQYoTfXqujtgAqjCksO495GxRqwdSBgmKtYenaLdMxXq2n8lSheP0UMl
NLcdOfLZFYrrAtQ+COMFUwiURj1D/8uEMRHj/XWqEyQWEMOFR8bOsc1oJlUrdlMRQci1RxvMzT77
qDWq/tWhYUnQgarwv2I2FIPoQVzivLwbb6GAeoyW6mOjbIia+VfCTkg0KsAFY1CmQdWNK3TXIVog
CZAvwoK0HfY87zLUM79N9qE28osRVpw7X4NdGqEffzyWOrdI+qBh3ryS78IYkXaawD9YAZqNVl6n
bPpkSvy2Z1vM2BuNXEQR71oviwDtd2vKaUoQvOZ5pvtxbAf+nf9iOUk1iCXzbHhLuScuVUvTs65B
E9DKZY7MLsXkeOESIQs18Rxof36vUDOfiefIXpck8mwrq9Oyh42XplkkbGhWIDqdda1LsG29J5qB
`protect end_protected
