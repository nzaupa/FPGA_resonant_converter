��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m��k?��V��6��"�"?&��s7.�\�ߺr�=�!�ѕzr�
`�-C�k~�����<bЉ�.�#��k��3in��퇢S���l��א��ET(/�f���&���ثC��KX1)Z3�H��x��w�!u�^L�#X�C������BԤ�ÝѶM@cb�y��J��έ��U8��+���df\�$�U����O���)�m~z\�JV�q�&)�x2�`9JCu��K��z�u�����B���(�ya�h�ѵ#pfI�͑��i^������T]����ƥ��A�ʛ8�>�w�7����IĀx�^�˾]�����9-"p)�AAxi�q{T[r3~�%����u�5S��܍5������#�(ܹ�D�e�Ve���+YE��a�'�%�V��eå��M�K��P*`dir�n>ag�5`�V���6D�n���T�K��~�q^�Q��3N�1�����%������f{��ZV���{�)�����Z�1��{��&�7��/u
�ſ�p'�� `u���5�E�9|�xvoS��̢�E����fB������-��ȥJ;<�DL%���2��e".㷏w����BP� �5�XxOQ�
;����Q�Ac��1�hy�[7������)�xxX�����k7G(���Jҟ�g��Pf����8)%�I�d���Q�&�4)�ɟȭ*��<)�v�D, >��P���&�������=z���m�b�M��f�dY:#��2�LcO[<� ZV��i|�V��28������9��|�`��V����h/`�E/0��br]�c�#��B��Ĳ;4�rщ�zM�1������ej�x�%4��5ZU�M���nq�?�)j� ��������e��G�Ģ��|��f�@�4��;_�&�1��{*-
����w��;�&X}�.7u�i��UUR*�L�{e�lȌo���6���B[9CE���~�`ʔW��"�ZG+���"��|�0L;�E*D��	Y�?���g4����]��.�¿��(۸U�:nW���$��zTPCzQj��z������x��H�S��?\v��N�Kl癕j��;Z��
��؋D��Rx��ɣ�s0�3��@���@�ﳨ�,