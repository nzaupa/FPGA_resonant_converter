-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0q2RaozJQloughhLXFj+tGpfjWxqfHFZfOcZyrUj4alyuSRQAg6BHio9UlJhMqBYnPKCo8cbxOX0
b/57gg6XMiP5mkCiiwLHqZGgGQDnBfkdCEWzTqd7wkOeJ7XCiNiYLAzgZEQHugFE4KgJiCWTfua2
wzoQVhjXkeE61WcbMRyKiOa48XirOkRKrgvYvhnkX83gqsRRp3htAKI6a3BPMgjbCnU8FNl35SiP
WSC7JInXPm3SJrObwTMxy91HRREhsmFX5ltvBPcLHdkVWUJLzMKaVBzinodcqf0EyXrzQFpHSSQG
Szc5a1WgZ0grgNnG3hmlnQw59b8L80KxygPAnQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7696)
`protect data_block
MFYEfG/xt0+7BjZS4kAdIOMUHx0yd4HOH8cXijsCRvlEgrYSxSx+x6eiEpfnnfbTQPpxXzU104j4
n/draK92h2CnRH1I9O6ZZuas65ZoOXjsQP8Ymmy6/FsfJ2dLsdms/kiXBEtWcAqgeeV5WEY7xdq0
WXqzAbzUYKe2fwI4AjtKTet+Z5cAWVjL/9CUXCrbueA0Ps4LiohvX8vfO8Eel+eixveJzc4rDzzX
/OwWmQmtP4hS07uSiBwT4i4+snqKWamoyIFEc4qHls9sCNREEL9SwOIqNxjL7943efZat86Wgl9C
9/uU+tDdxCmhVkTZ5OY6R//ZBhuG2F4QeTnGHW45fDXbPJwrqfPNJ1yo15d/ZjvWF0MhEzSxkx7G
bdK+K8MhGJc81lAolNmG+LfftppU10EXOE63g/lqp0nhy/W/7BLpjswQuhCfQgPaarqdBsTT9+B3
WEW16PBAaFhPgBXUUj+l8IkTWAhqnLRgwojNSdR49PknvOfYkJiLlr10okDAS/SLtcjwRsdoykYr
ssa4Df/2X0c5DtfM8LokRJrwXNBA+glK/gL+Qj26pexG+rzm4W57wcgmme6WPJ8MLQV1h2oekBMT
AxlKaW4mBxQLlIMLyl5ekcpkMVcm9GpgTNzHW6+LF0dO3TbHk0NV+A8llXQJ/umWYq9fxRS22LEs
DpBqizSQzUzyZn/UJp8kuMqmmSOVv0I0X5+zOGjQtEDvuYgGUSqSJRZ1REhN4WMBE4hUBPSMmdim
VXc8HsZEG2FpfwWWBsT401Lcky2lCWu1v5glPCDnk7qH+OfK1nWt/nY9cBw+L/9qT4PHWivsW910
6Jmc73NRpaXHJjCfby/EXgdA5CaEspg1s6a2UXQWXpv26wVIk3La2F8JeYjfjAjKfjV/y3vY28cN
9HwTCdkCJ3JY3ghqiMncCZsIwoqg906UPdHdnZPPqDOMllO8aaStm2kRtTFtlRRdo2a137mDSeKl
ygtxlcNZdp5j2kpdgylxDaRBMSvuXfPZiJDNLBiXU6j23GaUfZJvDOqvSAFDRnofi5uVaeTQQTf9
63wOZys4SpHJT1ahep7Ob/3j6ovvGtnZW5FaJkZAjKg3+Hqbfb8apTCyHgpDaTLj33Gs1lOLXUuw
85OInA4GpAuSjckWiALbDD2ICkGjn3AZDjXpZiDhIGRc/ilS/TQ39GR+1xzT2xie2yhBcsRrIEv+
w5jf9NRRnufe/ndEXlcdIXf0s4Rvzowg9fbR9r5a1DoH+fosNcNu281+0uVLLYB0BUGtGuEbmDFQ
JhXaGCRY8WD//ZpCo9TM4eIrcbExNu+93KGL7D9bdD8KBtVNATFtZCs+dBN2LSgRmy5tOHpKVL7W
Z3d3oYvRUamlEuHeUun1vj9v+qYP1XKXeRAGlDei73FjFDfEdUTqLOLHsi/VUOLZgIzRoEwk0q3Z
ta9/kbu55/BWlI17u7hlUmObxjFhqXitfmCgGq6oh30LiMOBBg8kSAmdrW/TEImA5+gAH7jnMTt0
kT7fewtO0qmK3PmZCfuviGeITfwsxi1IXsRKBI1J+4w5jry/MNpEdHqqvomMJUsmhWGLH8Cmraz6
K+2lwdoEZ1YZ3of73/4/d/z/n7VFmTBHw0RHvS16RnCEjfNnqhGl8npeQsxnuc5WWDcKtdyPFmb2
TAMc6D+nqbWdD0RuoktmZwhiawi+8eU0PkcfX3o7IvfeApR35IZ8Q9FoW9qWXcyfnBd+zBnkcV+s
aHLztpy2BmPI03SFTjOr5AFbVK7KiBV467h2rhuzYNYLihhLlqvDvZEdZa6tSwY+AmGlzOfXQNLm
Cmnd39gTDLpOzyEUDo4+nd1GO/G1tXCWZ3yYp5R2xVJo9bX5ZFcRyvMpl9lqf3oOKNpgLq8QgDWk
ttT0LwQTeMVze3x/CWl11VYYBvFAF6pAYEHJ0QvpmWk5b5fu9AvFzLOqHds+oafpBGWk+McuyFav
Prtc5j7VrZod+PAC2HxnDinrpZYeLFB8wNv8h+Sr0STggH71FkuE9yf/vyt1tdcYx6amGpEpbCsO
GRvKEFyO4sgn/F6/dSjoNxgrFRVYI6rvRozw+XLaYKoh0l0tlxxz6CMMrS/hPzjgO1zaWdOPzOKF
Dix1VYGFybinoSo2NxcEIEtiNOygikiyuftLoy5v6Qf5NJ/mnA1G36RdT9DApVDyb/Dn8ltaygok
IVT1q+oEWLXD6AZYHUh9IMZQvQ5C7Ce448Rxu3CT8qC4g6QI7HBbrHGu4IbwzPMUDpWahrHDbp8G
MvQcQSUWPobPuzY2Q/sxtTx7OnJ71xNwx3NH7LYTQaWAYKPa1GeJPQ48FjfHF91yU8gr126UAc9t
RSh7o6nSFFuK0j1/NMxoyms1rox6kx22l/c78KNq1pURjWN8kDBZxcmBGQAo7ujiAfyah/5ACNyJ
EInF4DTN6u92dpPzgRot1J/HwyZoKv1I3yh0Z6tmYdcogPm1KkmjRZZGluvovD6Enf3nF5hvQgJY
ulnU+qnHkxDK7+AZC5jJAyYKxNl1NJnRU7xf+L+2n19eL3d/1vZOYAM3nkYzYOCCrMo/Gmw3Ppjd
ENrotL3zJpHPrNMVlVSO065Mg6LwZ5sJzGEXY1NkqIZCdQ/LafuIiCuPKvaQkdYiWOawpvXts+Ek
LQBJ3Xmaa8I0ObpSud59P3Sdmdx8l4oBiVWQ2WIwsHrkVD3tl2kWy3JXGJqG51wmZ09fqsK57+7Q
fzLyHwLgo/KsDqMlMqLRxV1Pruo6o5661Yqc/NCKMYwyvbVArvFNRU17FgKyA4e1jGBYeAz9VdW+
gxoRQkkkJgTqukAf3h1ZGR2g8yXfeq9bs04rjofBFrIbbzi/sJmTHCJ+5lN2wT5VOQZ/3UTjDj2Q
aTTObNFgJrhQm+2EXwM0HT/Pu0WOiRH7H/wmEqSZEljoOODwrindjxNhUvN7t3LNmq+CRw+lucjX
rQv8rbbKGaNwJJsJiJTxBli91CvjhWxhhjFm9OcQ/fPD0HUx0xiRgTwo86qsaL6k23e8OSSA82cO
DClMagZlySt6sr3fp+C9t7uyhDA7FEspfi3MxpKFc0GYytzZymQdd7fJH2iiyK6HqxSQbDmIbI2m
7xpE0OhSfyk0hTaWyGykTa3XmsSe2xn0CB8+VL2FerA8pciJOQcaty7k1mDBn5Ajw0O4NzWzWKZR
wNiZvRAtBhX8n+02kmVuNbBFPr8yVVWYEGUjGDEnZ3yK0BIQ2SU7si4eeju8X/c+mRENim7K2ZQ3
wCAwTKc9Og8Hoc2ETuVE8vJsDk4m/ehvZ7vHvSsVtkMvxH52VAdh3oEo1/LAoR3OJIex4We4tfeg
6NoU1Q5ZeiHy8xQ/q5U/UUTgBpmd2s0nS31XszIbsc7u8vwv0xCK0uoWNlm8JUlaI8BoytyBA6r8
Nl0VmulAG/Glwre+YVRpHV2Cp8fsMkaHR6ed5FqOX61aw7pNPpJ0cc+DWd/DFKFOpflsY4Hb+4WZ
rU0rKEfX3yEm+v0nSW4ThPlRLcnzMREOcMFbxBL2q293JrD35XABxwHrRcTNfVT4HPiMX29Ngf+6
76FHYLjwu7YOJg/EtykV1BZA+oRDsSCQeXy/Vk6ypcenwcJ8NzV7O1NfPdSEU77FQ2zkZZlw3PxH
SX7Ce/IMmRYiw8Ee3QSEa9eWMPOlwCnr2kArOLQQTpVvs52NkpFD2oUb4QHUJSgP5nkrdZYVk0Cy
ZlTd9W9UWSMi5UUDHuPHbrHSRpYALwjkoE86L9tKV3rLvW4YhWxG5ptC/JSGOiiGIHs4POf9yqNQ
eimqznClZgjw4DvILsEEVMMHE9oy98PxPx48swZ5QUZzRaSIOe0nNtFQke2hFZkMk3kEpwbNW68u
O4/LJwGSGCPNByQHJxAn8YyNlE2PplpYYzTYL5Lp4o0I3ahGp2l6JoLxw7SkUmOKvHRYcGWHeHdH
f0T+AKP7pvHleUJtnMmDuNUArvlSbe3ONL2E2zy60AGzNS1fGzvZy7jBS1SGJr3nvwabHJ/2TyzL
AxdOUocFiw2m+EbT1b3uzxN9Y8Ki1hivgZqztQTg7suX2ROw+P4e0qAbrf+yc5kdM0QedZIqGKjo
N68c/TxcIGgyeAxhMr8xkcIR68vFc4qZhbwFtrLdoa5XUPVTHdCadL/IaWwyTdzN/dlkC1Him6AR
9O93BePGRnlny+SQ+5wNx5sUlr5xFQUBNg9Jn1M42l3I5ndEBKbGjpnlbdsCgSNLzB0N9AI5p7AQ
LzO2OHPQIG7yOjSL2XjieLbbNlDXmHxbc3Kbjw9k83116aPbH06VjKYyXqdpYZSfz9G/+M8aZxtA
csU5xhccbhXuH8zxYfRv/qGTAgLe5abr+v3t2Mcl/iyUSPLGrNSAZT/umC2zzHO0goo6zlTt1LyN
eQavTzi5dkkPhjOynYyOouL6DAByhm9d0TypfLoel2VppAM3OKS7m2FtswzXev1YL2TcAc53pC3e
tcMPRCcwoqgtpDOcBKCfKauhS3+MBk+KCZL1znArFXQwFY6zFmCQJ54cmSQoWbQ69rvGQg6Q98tV
oGoWaSvbBMIvoneCBvM7PLEYMJbanlpKsEnLjd7Jm1XifxS41ApgPr7GbqCekU4bhDpdgZ97hSRP
EJNDG3qGtSKv/vGvZ2zzLfWtNXuqUSE10U24clphZpjTF8acpYEgz3BPl383FNIEz8D+sYtT25xD
4XxIYBqIs+aewvakfixAOGzRiIk4Y8qTvOwfs0/jK6jsq6jtWQuW5hZT2Z/no22t9AaXYQurtcPF
mDIdLL6W7OyQFASIXAfcbj1Z16A0eyHzftUb++UhctH0A0bGqxZyFuLxfwD6AqktnCV+XvBR2vtd
fmj8fIDYPCzNZ+rJ1A68clXppgTY5pSUPQk8cKn9la8BW/67mUtw4oW0tWxMTQyZIgvMJPPa9UcR
mPSTuPm8Rf6+T3v81KCJknd7wPtZz87A++JAn9ZLgfRWLXlHVdB+TygqqM7Tm9fXE3/BqSO3hXnU
P3bua2m0oSlkHe7ZM8V15Ekxfhj3EXZbgXHZklbTlec0gFQVIvGCY4CjP5BpRilKduy66UbDR8xL
tO99d3H/wtEvGQPaxFixPlvMBr27oqoEDGeHvVB+PeYLkEaJf8TxDnS4jqPrkHDeVXkAMvvVoY71
FrobqYiq4aCs1EL9ZQOxeG3WHHDbEglLGDbkGby2H6kXCQFLJ9mYVGuUwOi5u8U++BQvHK9V5teM
1vv8DsWuBs81GcM53AW4J24AYgN1+HLNhLEOtVWhiW95BNlXdFeKjGRaZA0WOBQpwEQwZlJj7IVi
lbjGamBy5cP5DKdCBaaFxTVs1tCaqKvxy7fuysglXBLWrCVlWPSwIUfTnuTDbSfJeKlMGwr0w30e
w73bb/JiaX1QAjJOOyHPANkKyr61vFxQjZxKkZayEMZQeN6EBgP+cyF+L29VTyd6TW58SUa//qBF
07jfY0GoPJg1lzChXs5aKvA5y7pGp5Lpdm1RdcErsF9u9QicLOztPuFflJWOpmob5rpRrHIs5jRm
WfpCI8TAirYvzN21OBqoyDmP1hleNIOn428xV/m5BSKhwBeyEdsZPCOdGW0kgXBfyMyF+5ho9a8h
qljC5qSiHyMViK1NejBWD05psYlneukf3BEaJTlAda6A4/9mf2I1RkPRqPW9eI6G2A6zLz/sFPzr
uiUxvXD5c2892dCPbB6hAxQ2lORRqH8VfDno9Zpgc0lm9pxXo6nh64MqNcrFAkOLdqq1H+FDPJlW
rNFvMJWKfvmIgzEfyDmIBJyICBx4k+XOXu2bFuGuGpWiyeaBcAQjfo3W7vPDqyAXPtJgiDiLVIH1
F2et6jQrLorddET52qZeqSr/xIsW3FbnD8v4hee/PmVxfvFyEu6ftLXcRiOxi+jJUhW/ue2DRx+P
8MXwSLWYXFG9Z7+XsHU+fKeXUYaXvjPnJGLU7VDXTLQnWa0R3nk1I/aWpRYOXHTXVR9lgfZKmF6Y
aN4axk28K4IuGitFsOnSoqQKIzrWxWhSvYkIP0VBkArbARhjouaPCMjCAJpg5nC8gwxuf8Clg79t
HphYaj+5u+47k0ZILQS1y92mD5ySHbK7bbHlAMrypP9xoympMVpuE4jLMQtBpkpwjAbG6VVFtfZd
bcwnBOWtC7mUTZQNqw2p6f9fDylpt2nYnuFHX5g1RdBTRvmDQ53pVNblaAvJPv8j5DPV8B2jvsI3
VATMlTfCVcYGaTjpD1f9w2Sjn7MdLpw7oMjSS9ccy4gGd1Vq1E+99Z+HBe5RSNnO4sGL1IO9nMNM
cJlgmWKP48nWEvV+nUPAChH2IOqBqBwnfH9RkkHo6tgm2VDlGbx91aLiWuis0Ihu91YVL3EBvKYH
E7VS+fuqiRtzKJWkiEXEj33nDerCaAzLy5+cO2lP5Vuxb5dQblJohLK7m5Jt/ohbVAjoqmbRY0WX
G0deN7z+K0Xoj1SyOrqOmCrijqBdLI02oqYe0w5NBwTZcAr3DU6h9JdUkXF6POpXgoaSfMTYSaC2
Ntc3leM4MZMiAKFvyA00gxQLguJRsFzHp0DouPfkJFhE47zwZJJV2qe2RcJkCrhEpVcNZ2zAPACv
XgLgpJ7F4lOsEfwNhA2MuEutuy/zDB5I08YkM0lUpgX4c8OpfoGVIqDRAY/8PK3fjw3MHPZT/6Cs
/4dE7YVQOjoi3q6qNZTg97MdQMD8LLL6jIKZoEiBvXXc19QtgWjfsdpVX0VXGaaWmkXxPqrRV6dB
koS1ZI+ixU7E9skTECSoI6P96iNuhrO/Yae/PPckHlp5VQy5l+lZQTCcEmnXa2XCa9Ykusu9xphL
pDgyV/u6fkBwg4Ou9UeCOoUZ3nvNfTxLRLIQlTK8dKFhyMO01rvqDAelxavhIaQPij+xNJE8bN//
FiWb89OmvXw0Ad/T/iIHr7ZHT5IwcxoQSUxw91XH2Ftu1pWLQ70aT97WBYqZArL5Du2O/u1hjpY9
7+EIUfKjCJ9kuvsEySB653ya0NAOZi9+OdLkbv9w0IJGvUk92pF/T5wzQztwHu7ZsAMfpANZ2RR7
21TTofHjgfgXsNLd2bp4Fv/ztwPq9CpdTBbeMRSTKq3CAcvRlSTnXtTTpiJND1tNIZQyoBlPzL+G
yz+Ri2OWMMylZGKMSd2yiXK+bS3nKcozHuulDwxC8LTbpIXMrXIDZk5I7ziJN5pWdP1btp19Uy7G
atpKMNqcqWdnKX2nPBe3IQC/uZC71WZgwOBDzoaEStpctmKximRd26Lj5Px0t1kU1e1ZtjBU/gHj
Zxc7v9eLE90gXelF40kg9W7NnLHsjoUlxTHkHgr1MT2vTTA8LgJU33ohx8xrs25bFmNmKOrgjIvj
WXqDrSnV4wTlKvbrW+6NJ73w9w686JhYo8u6bImjOs4cwtkuMDlCacN+qJ7VoHSVXCnT2iitCo/R
+nRTyZkr7nZlERj6K9liGhMDcQgLMoxVrsPWNxSTdPRnfJYHVt2wyUcIJW7yg8FuQs47Gdf4gXOn
bs1QKTUkrvZ2pNxWVMn8h5delkx3y2Euqs/i90/HVWZxBz69eXvyTEymq+cvZxiC+9UrusHS2haK
VZC3yqLcZNrrejSqgUzVyhUSALAStXzllKRNNDyi310MKR+JRcIDsT42hBK67n4b3eoXIsU+I/Op
E6A4hY2EY9yyYpCdffdR3VTjPa68yUhBX2vPrL3NK3JPm2IU+v7T5R5Bm42x37/MiH6rmhtO3DLv
BuxF3Ckl030rOBqKPA2xrZpeaoJ8sLsaOHnj/+PtITakU7Hxl6+zb6wuXxmDck7xZQY2aAIWnjsx
nuqOvRaizL0zmHuPUC5vN6Bq6fLyxjtw22ExdZlAtg5RnhJf8juAzsVO8zpirJl9iGwG9PlherGT
nOfT7VQSzxCt6jvBIp5XH14RMUYu+ZzyGAv6qyfPFMLnhhaB+UJ4MojCG3YtyxjHpPwPIRJtV7dC
6qIhRt0ffW0unmGh6LYpcuaB1Izjt2mVolruZQ49hdfXZ8pNwxr6dAWEVJQpbGtp7zwSVSmzfevV
ri0pMUfeCFT3rRkRpUegB96/6r+NPnvGV0r4v/nSvXTZFugqRlovcDtONIJ+5NFtAzwQXldZR8/9
rv4gqfePuPCWd04gXVz8ALbUKUEuGOnd2KW31y+ibpvJqCIvo4NjaNaD9vIUpLX2+LN5kj+huB6e
QWdCENjBT1AYlS/4mkfstUZ7hHovIQtopOq7TcEF6Vx+xLVK55B6K0kdFcTaubslb4aSvPjkHWOK
Oa5hoHOK1M7ny8q5e+x/NKvbMOZhVtT4GNMS23umavwX3PgOcvslTyjoFlZgIQza7IvYhMOoxWWU
fP3J/9G9h8/0bBO5meFLwWNOcBR204cp7Yl+OWlqB3zkGprEPkokJKo9keHnCmGnzViCq6f+d2zB
TIhdDAYUCu67bfhkQsHCfrs58smwbu45iFpvH6qjvMmhvKkj8RloZ4JACLYsBLlv4AWug1mJ2sGq
ZsbN86Xu0OwKYKaEJXbtlPOF6vO20wXR2V/cQ7g+3vcQ/pk/k2cgWIswuBn4oCd4CjJjTZv1zI4v
qhSKz8NSBgN/mpGn3B2qsoqjykShCQhV9N+ZgFbZLM/EwiYHuJgJWXX7MXljhlg1OftJkpPWpsTG
br1zp1LLMzltBOttX3dJyJOvetT37yYy4KAMbHDqE5D7oTegTmb5WHKoLHaK/BErk70TiSf5Hpkf
kh8tD3Ee2XybKD1Az6+nqkbI3ToOW1yAbSQUPtXB+K7wwWNrs9kQRIs/NQNSIdk5P/OBv7hc60nm
QeW+JQFKbxcdQkm39flmzak5KGRjAbW3ee2CoO9nFufstZFEp/dN8sUzD2V11o1D1vc67IWJrkYn
J+Xy6beo39GGHxAHdg0blhDEb5cIjoZgWy2I/IrEROr9kStBwiUtB8kiZj7ZfsZA+4KjF/8Cb5MH
vIHVeRgguJ8P4smGpxHPN+hGm1qRa7QpXBsd3NvuNTx+KaQo2x5u3YgFDQVy/n0FdG0lbgNnZMzT
yI6VDOo9//HfDpSYSf2bYr0chiUaHwBs/dNnXeg0+zZ70QHbYBF9D9xnFLtHNu1AZYZ4oJtzFpc0
HQJb8TTgUIpDV4xGm0yDF+KAR15k1W6V0NeLkX44eOSfUeHVGgxBmXsQu2RezPIBzn4y0G6hKYVd
sVT0p8tFeK2fphqnzZjsppPSszHKGU82MKlNWI1CW/zh74HtAvY1T4pzMlAx9VTnpEe87gxRyf6a
37TqndHtUMuAlE865VmAfO40elTAgZaxW66ECaBLcmKbAVDpNJphbC+Zk1JLEyA1z24ROdBdUkU4
kcF4AWVbhnxmWA9LyqyXLlXsZQf1KHjhaFQ3WoLWhswR5a6zDK+bT/FUMx2aZedIi+fzEkVXLwnl
PtsFrPmRHeUqk4k0YYqNTnDoedhJ0tW+OijTP6kMzgu6fbGaaY2waJT1twJMCo+aBnFEIzs+FQxc
JloB0CIawQ5TPWYtF5DcxcdZlHFawjEHZluQXBNaeLTr4uvleBLUNZJW9Hj8TuELDzqRNUbaCqeX
Txmzxtxj5kZtcJILMxYMF/abm0B3LN0XcEyRcTwCf8W/EXCql8wukYwaklr8LnWs38im8gr7GgW4
SvZ5mvwq3Wm5UecNj+bnMouLE+qXRWP/3IxE5jtnwPJrs7gUH0s8+KeNYp5NeQ3vaqHjlQZXYPKr
1XzY0j2kOepuO2/9acvwgGxQZnUkP6WOcT1ezCyb4fIFo4W5UfQbftRfO09QCRBqLTeBF2AaWSlJ
2B9cWxY/7FyVAxX8hiGPBUP8FBcBjOXyoQsJeVtCMuGKxwQnD/CHTZG0Srui5zeqa+L5KMhfV+ZI
MimSnlLCDztrnUDAtAmBBmxkD7eXr5jFebItVOdvAAhelUeCO3LEcSvHrCXhqOnJvLg8V+Na/sOs
qtuGYZWQJNHQaqnZlzlZjPEeUnwU5m6vYR+Q9sBhl6T1ooLGEi5rCEXRYFVIllLT4N2hclIIsBbg
gS3UCGEqw1LNzcEdVf/8VwF93okzmVYuEujt0vuJmy8hZZPvhVdVXFy+LYacBut2Z2hT41r9+ig0
YaV15EI6wZK/qixwbg0FExZ9QFP7+ASZghPrY6jWCcczXUq5geI91zEGjEDwv4jwnzybDopPRWE8
8iAd4QNsAor4FY50cj8GKmkiyb7+t/EQfBtBSC1RajMFQiuKnhvgw2VI/hrF+XpFQkFpavAZLTUt
vw==
`protect end_protected
