// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
DV5wzWXAOPv4sY1A3UPVxhXkzooxZs0KT2BbvKLjR0BTOTfGpHuWmPRpsC1AE7j2ua50ZMmCbg6G
gDXoOBpg/PgBG0yxhQGScEf9Zm29SE1Vg7wfCoI5O0LrHpQ/dfySWpAh0/mlsutC2JxJMx8OnoFR
Q132cSjyBuWCASlwa0+O+Ja1YTZACIQYO7AS0yONQV+CaLPPfwERVqsHw1pXQy3/DoC0nvdW2uIV
fJ1koSpWD3Rj0x8zWE3sNx+/C+A/t+UlH7IxoEnEEaxb0E+nlTUeyujGYwU7D8pqQ7Xu2BnnfOh6
SzoBFyK5H7KZRBVGWKjNogcarLYimWNQ/3qmeg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14000)
N6FBx77jP1ctpDkyZPSO2FtOLPAj7guk4Mesylfzh5req+pYuxadAhJXJmPKwex1ltTKD8FPnczh
92GkvwSm9sIHnufRAKxeIavxXZpZPYgrUOkanEOOHAEQrmz/DYemFGNhp2id1qOpvB5y2/SVQW7e
4enmM6rk7LC8rzSDWqSBQ8p1zTwADLACf+jge4pgLh0v1L1UceEmaiXuXq7DwRRaIFp6CHs/NNHL
lI8Ep/i5dX+And0Y+FD6hVsw3IqxvHtphupe4lzpbC2JtfHVoh8SnDUtZVOAHv5TXciPngOZDkdi
/+8RSfcLYFrvhRLeh4EAPB1KhNju7U4yrXqcCW6PziyH4SXJ/wJdc2FEZZvUvwOPs9gHMACmsao0
YwvE1UvppkTsRXFwcXuPsg+tQuK0muqDprnpMUlY4Nd8ZpVRwY6P71ehapPPapsmsvbUiERIph9b
Jfn0nlya1ZSf8ZmT6vaSE+8oFT40RQC6E679Is9khucJ2bYe95pXx0RWgkr5DQFdMxjDvuaZrRk7
293Ke2tppXz8qmj5TPkM+QGsiWUDkdWKIZN8Wki0CCYwerDvFj0bDi3AZ67RukZ6zoILIi8KLQvs
TvA+IIz1vQutU/ZOcb5/npOdMyT8IkFq4iSZZzs+SSYwe9AD6P8UeDeDJASsVbTNvMxgOgsFbfPY
E9JkEtvkqAM0x121Ej9lcQnuWzOOSjEUPg/l/p5jWSZcwloFQbjTuOA9JB+zakqp1Bpof0lpeq2L
EOzC//a9RuyCXOBMCAAgPgG34KA1fE1K8K5sVYuz+ADEzeREx/DiMez0mTygre/IL05xOiMhymyG
xwFrraZI6jBAPPrZ8o3awfa7StdcKzh53b2Dv4Gx9lomxGH+PG27tVDNYe++VyeFOpAUuDa21zmT
OQwWfM8UIzTXGZ2med/bU9rZnvyebWbyNQO0WieJaA6puubqV3gKrM8kScilEzi+yyVsqC2EOkID
f7DMUdGaqgYxZTP1KnBToHegOjwR0cUgraxGnnNAlcFC+OYV1qGovbu4P18jHVTAe0ZNAZp81aA3
86qzleH+ShgTgYw7toN+MW8LT08aawASLpzGnSGzDGn6qikJQuP0XLRDGbqPBt1iJ56qavrxZphW
L7mtvCruXx9s64UZQytOf93BYM7oXe/qcJA4rkY7K+3cS9PmWoG/EURTvOues/78fhpsCBAbBL/w
6F6+sA5mgBU5Fudqg6VyrqfZX3vNaY9Xg4glJBPV8kfrPkd2OzIxjyv5b03JU1nbI1k6bLkQBrx9
P/st1v7bKOdOsoTe7t8HSnxcjMXTmQvOyXYWiadhfsAWnOje0/XntvcAeNI9lu6pmo7lpPWFyC2v
GOAJ1qyyUwNn6cqmzqKaMn1G0Zv1ELxznXkN2r19MDQf2iKQnqYAdivvCxlLz+C4cfAuafmHsAlW
fmQOczT/Jp2EvNYrzsXREOeaUFeN1gx6XukPsrVNmGCfL/r3FXDCnAmJ8FzwljSjW4mTBp9aymOB
12v23jxQbCb9MLF3sE48qiA75YhuFEGQNTev2G6WZMG4j4g92Lhp0+J+ZtSq3WJlpVTDkazzGQzs
wgKwHLrhQP/JR9XSBvz1M+uRx1yLEGDdjpL76YZHH/o27srR/VQ23ibOl2z1r3AC9eK6+qArm7a+
ryy9R68zmCWMmlJ90CXl77wzscaZ9VwLX+id/AKaI4Cn+FSkyhVCWl0tBd8oS+dRMM3sSc3GMot0
yLPp2dCM+qZBDF/6tiRWn48pu9ELW8oUrHgeeRbv9OXQ52WQ+F/1DGbH6rR4qAzYgjHHoQONdUNA
VZuta639CAzdnuTHhboGaA9sqa4L9d/8w7iGd5dsn4i/g1knBxo/me/Pl8dPPoGFCdCJHDwPOl5b
xBS4Oe8fwRdIxuvsrVAXPOotvvqEEq3HqlhWnZVbpwNLKZyzJKLJZhrhC2Ms842FGgYtoEP5Qy3g
Lb+ifEh1hIlAttRwGnBmNyGzqbUdJnowVvWgdckw4ShxHJ6FnaCx1KL6s6cohAFYkU97cS/+dzH5
nj0Qz3TCEUltAqAdEwD2Wx0SQ2RxdQ720Rkd6MjVuMWScgr/v1Yq7fxmsIYw5HJh6F4bOewzu39l
DUP8ht1sUS11mJceBdCNQlN5TQsPBkuMCVVQsic3RtBATPIG8oCNW9nDICvQ1Ga62D5S0Zj5aB9O
ssw2cO5DzM8hJ+nQllQCmb1wF7g2Iq3coBbx7RrzjRQwy0JQgwDZwYXTujUoSiSJLTiAlvvbxuW7
rBkl/T2lJpTIEqGcK/yuHV+gey3/gkjclQMDIYhf7zn0Lo9ow7Cahlvt1Tz5f1jDRHyjnfkKiUIR
l7+TEu98hGUMjx0Q6wXnmU5GW9DSKc7mv2Sk9VW38yp1oP2gNZUL3/IEBdXTxlhC2k87VGzB6JkH
zHbItxmeEcsGfIXN7AO2ZwTzUh+IXYQzH6bVtBNmLFQrh1HatIw877XVYmx7VfhVMACB7xe9QyS2
mCflmryBfDzck0HNJ0k/dkFaVss7sHDyPfP9UiG/QXq7/6vSuTNNE3JE2fyzZvmMNK5H4H/uhfSl
lNEf4Tge4lR/U5eeEKl+IgELlaiqEh7T5aGxkJ1zDHy6aVcXzPIr9mH8DDxlW+HRX2jai8nzKDRS
vKqEHZi3+z08zECRqlSrKsK/4Dcl948t7sarISgCbcOikNzoI4uXknAQ92/nfdAK4XmgFGvss317
vrQ0VC7Rp7Fw8jWDhpr7//Z1KRMPgxGXC4p/zLv243WfLwqBXc3tOCz50dLzTCS7I+YzCPvcQLLU
OR4oeSY7bJQhB9tKDK0gki1k+zf1E5zDK/JvHkjcB7HIrxV68MDHT10LFC+BzzWya1ryKmmsf2R6
T89iIhakctWt0ovuUzJ8YUKrOqErOSj6D9qu5oCiMIw6JHdEl+0ZRGZhYbThXzxlQNOB9C0eF3Ci
kL0gsDx59x11RyEEVSJi2wdJrG27+PqYLURzTjzezmwiHIG55qk8bhlDXTvfonyX4bv6fTfVVptl
W8KOuMvshnnzIuEdT3oizfrlC7U7beEH+BGTuBhj3PVsVK3bNlkmSIzFIrRm1tJoOVCPxqjGxz7B
WoKS3g2UveuGQRlKWQv/7012Q1mfw8DzWz+k7jGO/RtqIUqd1An4JErLGDNsXA/h+QjyquB9gnN9
iwAF5xaLY8aXyJp2yXwwHVtX1p8BEOMUNyStIqsljmZ7QCafByzefYevc6Z4wCGDJdLUgHtMMt/P
/o4bnhTj8hP76+XP8mjPoaAcU20FUDV/xKKnGGrokxOTnFyvma1qRwHxNRIfiDM3+gM+sqxzeYPN
57U1so8vio8lM3DhbVicTomRqzh9eK9gxwsgxBPBG0DVhIq2E6SFPSFj9ldA2Emhh+dYUxanQVDw
QQ7f4hagKcd8cYJY3ygqvGrl9T7DHXVvm/R8kIk8MdFqFluIIjiBxGP+Y9uyqIcMbKDuUPyUeGWg
D4/hQFRRzVErIRbW1dvqKTPGpaEH5qo9QgJ+RWTD2SBdTN18E+eOTkoN3PgV/xPuDVeG9wnhE2q+
HSfbTvMmrG3wwJZYk/8FqVqGR3nZqP5XeNHP7UN5nVQNP0tzpSCza50C5YAkkpQhF38fDHEG5vGy
HB7SYkib1/tF9VuY3n8Xu6kyuNJ7CoMkwjZFQqMLUBLJjxA0nKIogbem845Vdcoyi5sGQ1bP9Sgo
cLRkBXgtMuMdWUbKDeWFBaI30W6XMGNm42bacbRdrxDq0NBlK2SjaBONfy2ZvwTd7fihgMao0Qjz
eYIpzjxWQvYbl1qvkrm7FyGtxn+EFy3eEcGYOc+tqem1b3s5LrkJG7Ex62lrhQ1Dg91aCzWm5AT2
tqSVr3s5/WZ1NklsXHtcAtqM/XoHoi3q+TpaoPDZfZ+eMYownqmFmCvEOlf3U4MGAWPcoj1XIY73
62IUNR9/S2IXc+G7y8y4ClhyxdRvwIpzEU8gbzLFOQcNMp+7O5G5LDJqrQzDVevOlyqmAr+DO5XJ
P+rp3ni3OU8mz4MRYyG60G1a6fFJl313v9kmQsbS3CyNiDDwYRQfAVxli//pEF84egGIdk5G0aCd
QyTN5MxbVPN+Mu3ixw74ytkBc37pPFmzl/Dh0J4nSQhroChnQUdGdcDSs5AGq1KEln57PnPx7a/c
y4v+TCIV0DqUT6HTy/YIeTZi93WOL1S0Bc3lEHtSqXnFJ8qQAuQ7A171XJUwEaBafMskxK1LSHUY
aeQEFvLw4NJMqlUigMhwVmaE3DjIjFNCQHk/oNoGlekLzKivbk/ZdVHLehgFjL2OhlSazuHMUYyf
OH3oq3N3MFBJ5tVasfuRQUMMv02TtKFgstDvd60/P9JWBH2msX914g+UywLInJ7V3m1Ez0Zlopg9
5Gq3CuXYmYniIYnWR6XL0kHM2H5ydhemXHlIVA1aJR17v+eNduX2badzO0EKEFfyw4YB6YeR3i5G
Fo3w4Etf/LenVtkEmVTMyLkyYH9b+zn5N86kDTpog9nRcfDk1jR/fL5rg4tunu17Tonj89y402MY
o0n+QUg1T4V5pRjNqA21O1uyep1iSZ9jssbgY09vOHwHrC9Q5pCb5aSSuAgJ22LG+iqEwiauVVCv
kmtn30oz9veLikddxvnwOJwMIYa5YmuYW3YpKImPmKIqE39B0fV3jVKFv3VcsAEW1uTlidNTWbdV
zO3OGtdOAw+rxmJ5/A5rOLjpAHJACA4LRtzFSm9CxGWfn5IaXYNi9dnGF6tZ0PvyIN5jD2Hrtbxs
u5DJvBi6C7gxmxZs/14/W/rVWMvJce6+Qa4IRicNAVZTBqVt18y6G6ZCC28/XOWnN/HTae1J7nhE
zwRBQEGplrOV9rcZVGy4OjiVYhfdLcZz5s//oagI9XfHpTaEj+tNpET8Bg8d6PjiCXNsm7BSNMxk
+JuPsELUjripfU8YltzMtACfQ729sj4DFZGCunvxQh3PklMBmr+MEtzdWXKwqam9xAH2RBZzwniQ
mV5S7ApLLLZFZYyXUIRmUGqzVZ0JHjaGWqbceMZL6X25Efr/V8k50SX3gHKP1I9JIAFMBhSbUymv
J2dy3V8LYaoLTTUIZK4mzAhBEMKOBgl6qvAcTz2Ey/Fx3KoSZvaU483Zo3Jp4JEZaXcmgNXLP+r+
CpdpFWwUEZVz5mDeODp93bGgMBCbmG/bA6YOe45czR/dmtCTDHYu1IonFndRfR85SNOOW15sNlIi
w5srJ1Hx1zdK92LDnd+hL/vyQd6DU4qbaimPBdqAsmTN4jQMlFUNDI5bE/MtuSoIoUe869QERe+R
170LhNDlWb2ZqWdBP+Kbe4mmZasCithIB7Q2/KkM5fyB29I+y3hbJbsOT0fFgpw+HFdR1iTedSGh
EM8l9W56QcXe8au5IvctLY5gQ2XE0KeiTPPu8uQ4Ep0wWbicU2cY/m7aUWk+wGbzjGT7kVDMvQGo
Rh5tJh6+d9Mmfi6pVMnVJwNnTqzICB7q7qidXNR0EsBVod70ZRGqtnM7AfoGuxtYFjgg4aNOcrRc
5cHmSxan2/Hov1lHeY5J9TyvRimP/UkMRHFCCzwX4t5m423H7x7iCI4fFEYTAINgENwRiyXLBvKk
8KFl2W3VtLaupWoB0Jg+/O6G8mozgFPAM/S0wCpQmZcX0aHaeXIu8Vzux3E9KrIAgx/+HEZqwPZP
gIePV2vHpXJFXkNWERNjELPmOowHbTuohhufXVLIGV+XoAyVTnIM3brG82poJIeJ+kQcVpILDwRB
AOvnXawLeUrIEtb6PoPOKVgVk/J38nkK1zm5NEcisAfl9JVivc3Vby0UO0olyaip6mdvwcRddWbr
BUtnA4/j8LJFVkzmdS9GDMUMojRQH/kEthKJh0B3DPPrReNSmMMps5wYlk35p+R17r8N8UpUjtaV
FgZP9cFlTYEKG3Yvdy4gTc9saTIyrZ84sSPhzX2BXNMBOIs2mMFog+72KgfRxhXuADHdXRhrZrKr
KPMZe+EqxYdCzst8Djba2FkURQM0zFKRV0yuEFndx1s2fzEMZlylFkZIWsB5ORrqQX8S6NOeLQqM
3YgqoLf2820m7BkkK7oSnPcbTpTreQFi5Y1rFKF1VqDzGmXoTkOJ4poybxD4pfOYNjdCFTiHyvlV
ns5dE93NWMAHeGyvCXKlqqtR0AkksTuBG8yywk6mt/MpJhrm8RZTiK+qVZxRmpa4/Qx7jFURfrmR
I446zkJ8m8oOH/oC8r4ptKygp3cmJM9vfUvGW2yZYay4ZBesPCfi6fX2hqUNYwqIiA1f/l0u8amb
z0QoqNx3/547zkMb/ZADj6DMxunqUHTuJcD5kDlyVL6uCTZZrSa6HqRpzBLTUgonP2PMARGDa2H3
AyILh6T+ahQTWUB7avljYmcCHjK/gTk99Dc1cFV8Jt3vA7ZTeqoX6fmMqFtNjCEOh0kjPWxNW6NB
rT9E8L5C87iUU9WoPYarnUZey5BuuZRduN6PqtXQlBSbfnGmXVK40mhF1tIuSMjK/oeSVFeyLkZR
ODcNxLKUR3i+ZiiFLvWyrQOYUuljVoX3xk1g/GcpfjCYmvpLPiLZtsMjbqSvXxjq2m7gFQwBeqeN
Cpj5l9XMJbl+YHIrSal5V4/9I/7pD1Zo2OVknnxkZnzzqPhZHP7sA1hyJNOV/pOmjKYz57G28yf7
VWtG0Gguy5uTw65RPE+gjV2MAbKXL8Gue6sxjqFQ0Ll+wTZhNHpdvIEMoaGqOE/gU8VsCamG1agF
fsWc/fKbucgXOcEtBBS1f6a12M0EpooB0MNUR+Om7LdeO05Io7WJcb4WB8M95tngJXyllUIal8Fb
7rJ1UpYl3XmOvQN/+vpqfPDJcGnhsvA1Y5CTYKSSHzfikCjLf9HD2uzqykD1P/DJQ7qVUuqzzUTM
eP6H+kyudlW6cZUF+see+osBsSeNxySFjGVQ9G5fl1R/dDZ/0GwgusKVS3+Xu5SZHBwXyoO1iGLK
A8k13e/P0a6zCqYkIvydEDwCDbAdLoFen5M07YbitNph6OysCaoeUKOPhAOFKB4pLU1DI1UnDZ8u
XinMaEbFp8vXTYMHr7SOjNtJu74u6KZk3G9ta6JwNi3lVyla/sKUwY8jYaVaOdb4+eme28C67zso
bGCLwLB41NphjpC9ZCSehNdjCIkJdhVmedYD33+abuEvmFdq2dKnWBPWjo5AmNo6Sz+jbjZTRvzx
Py2jsbJLtOA+gTOBmdYxyGuqoO1afcFpMelvgewIYbQA1LIqtPa59cWoDvGGils9CmTTNxF9M08T
YwAuAn1GVHzwSXk3DO/cQUzrPo+tLroDzht+NXYttmHXWXlJJka2qvfiew5yq8qWdjfl5a6dmnU1
iEhDbM8oUvKOF0E3iq29A1slOySaPZqMpb0imIsMro6YLlHw7dHOWd4TxjLLeIxMJcWA0lytey2r
4P1afM0hEkimIQEZwHFeyiETV6SVAqt5ca+1L/KxHn8RVWhH/lgL4zeuyMJ8xN3WryPG0Rk08uoi
/sC/5PYRStEHV4EbOiD3Hs5mwtNGpNi2UfbXt4Dy0miJAe2y9MIlS6jGDGDKDJdYZOCi1QVMiy80
k6Jg0hmm8onwkaxfLVbUB9BIM8aczKX+bjw/ThADl3rS0DRQ5GtjfrgUdDQkYDcCNLm9+525AkoO
KQmj5iDxoGti7fYzSoXRM+lDx0dOikQwiLyPFF2CJESLCoyxMHmr4xkP3djdlgTIw2ph6ZAER8Yk
BnwKU1gIdbFsTEEUirOoN+GNVj027HS9yuUyQEwOKmQmIV0sR27U8LHPd6RUQCucyBKPWODwL+NJ
UC64wZFi0QybWUHbiOXLGXbhPTatcIHO9d3x58nAzgW6z7suJG71buPKGuosufeqW+CKN7Na1cre
EdfC+G21LTvq/pWykeKEeEGM+m7vwpq0rJfQomNXX1ajnnCUobJORvqixJwMu9upokMdNupNHIXB
Js6Ocm2W1okAzEVKGdZkcasW9jjV+rARjlNGAhw6U0rIIAu14+8r+LDJtskSodvK7OfcbHXHrh4W
CbyHFHdLM2RffcPGZdJXLMn9RDQtAtevkPTW8WLQ1YPMsCfdScjORQPYTV3xOvn3R6dCQbk+ZoMF
APgy5FrTwCCzmfQWj65x7Wa7q/Xn+RoGjOoLHktSCKAo5Inw1Tu9EJufRYpVJthhFMxJ2bzzDvzV
Zs7KzQ7KPMX6MB4a1fPs07HKTid3rCdO+sOvhP9Fask7omgxYXZB2RTZHYhfnSNaLC7fVqkxdvfC
4gQsDZZ8BRIZQckaZZzoQv0OBD10mMHJlxR34rMndyZj+n2rAKrTsXqiysYT1+K1qr/kmxF3O2na
gzO+XgWXGz+4yyk7Z25cUJ1rQsvvF7amRgN61E8IunNMAdBqwdtWO6whR3RdBpsj14lG+J7QIJ9j
0TG1bwX21foh+V9aEJM8lb//+qbqyfKugKYPpjrk3JJoRi5YQQ/Wwj6JYrUugLzirLPp/Unmuh+z
vJ2BEbyNmFeCkrvUHfzl2jyMcmzn3cdHsw41/IboigGMwDIC6lDcjjnQYRMh3xE86uLpfwzVoqzS
BqgL3uGYZvtQoIujH1HxO+4a6fWvS7BuiOGrSY3yCStrY/0aiJimTIbFgb0AnG1FJ67iz/AV4seY
1vNqNEe6JOtK/Jmgh8rwYlJes+RKL3dP3I3MFXHZ+prBg1Ax/HuLlOCAiVyq2lS71fRU6G/m80ph
U59IgP5MV2uFFKTB6eQHRR8l8vwX8DQatSkYQZBqRmwmIyfBmcm/cjUiiTWwd6vuTNK0GVGM+LPs
cNBaynmNI2m7PbB2mKGBuSYIttOPa9/J5LMc4mBN/O34B6li5VxuG+EhToK1/oGf5gjTKnLzmM6F
Yk38xPqpWe14WrD22OMptAfLoW5U6/vuATMS7cfqx5PD/tkxcPQVOf0j2rPPXBp5pUUoPvoqv/XL
Wr52WvqEUvGtJB66DmONaZfx5Cn8xH7mIMBl+LKphJWEk1UXu5O3Luj+lz4wjq+7Q+lLV6DFTkub
k9z5LQdLGqhBdq3Q6DoXA6xcEJ/fetQa2CITVOOdyVNQq6radyQutzTmFQ/oRhxAateg6bkfrMRf
JB2o9ArlvK522ZTjXMCfIhBc4955tSfgI2MbyxpcT8q9BYtGRrsS51t7WYEMcRiPpxnr+30JyiIP
HCnbsDhda/nJ8OxADB6NN4qmY3Gm8kSqRx9KkBQC4WfPhxZ82KznKy0ftfhaMoRu3ppVh/pJ/x1k
BwY+m0zzZvNi3qRdpX1jFU1+3w4pROK67aU8nho9UVuXZN8UiA9L9R3T5wo2rkJ7upqIR3wjW8IL
7b6E1FZyEh9JXi0330o8q0QThOlTmjXQQ3UYXgX2a0fCO607vFYjQymGp/mUH6MxmWPtxyvyOaZH
c/lqq1BPUz57Toh/EAWws4rhahWX/4BQgwLe/+UlL9bk+Uz327uohbo/D353Uy2a2JRjjopDBKna
V0auE7EdaP91liS2610YxNrhfn52INLprXvkDvuZpv1nzcO3uzyJg7LoQKArzrpiRo3gMYT8AwqH
XNHhwSVH3lbPRPVgn4gBVYjRY8kchmunCU9uy9dlWbaorFNFSWSmGAD9XGK1ZGc3g3RXZYw9J/Dh
8EBbwxtWlXDG990nA9u56I88SQasK+b1GgZqYeY6kh2jA4djmiyMl7qpf+gPDAv9PyR0sF1GbuqV
z8CRMjCtn+LBW7wnxu7pfjKbHlBAwMDgyrePg0bZf2R19djRoHa9MC9tyBwroolGQATdCo9WEsNv
aDNVK6suHW8bFMHfDT9bBEqyFpH/rxDDxzwaIRz86LvA4WPVcOyEU0DgzW4FuTUeZzKAhd/E1tQC
4wuMLrVBJ3WIdkCPL/fV6LnjGnjVAqRchRtx53W0kSohta9J9JypdblXnZoUDlYGwuUmuscgaaLG
uN+7UoC0dM/zQ/vT3lfa9qHdwDHed0IGcCOYJTen65t5OYSvJuCDQvfBquhKsZlCj0H9FoEDjH17
mV1TgjpUXM3ADqVwq8T8jR8AbZcJzoON6doCMMBhWewjNBkclkD5jMJKqkS63BnNuRO7q8ssWCVY
xUAgwS+pj32vRo1cMqS2Ya/X3buMewwseIH8EpKtlwI1g/B+Ljiz7kr3c/38T1i0Bt3X2enjtC9x
wzrHktv2bptI0NyG4OBHyTvLvTaGOiGf6cdc38ZLSWBIFyri1DFlyvL2SvYUUwf2lbZ609QM+MPP
s6kIsMq1QIwPZnwNso8b764Kj2A7WNvFM0Omp5FIlHew581TP1q2PBF5/4vb/HCl963DD4F70WTK
GfAno26fmuAARweXrMRafjpwFJmilhmc0V+MXLRa1eFZxH6S5k60fS50LbPJpHX7O57vu/aXgq8O
cFJ2L6zy6wU3LPxCDABabeUxuQTCKhhrhuXJDfW1HNzaTjtyygm/XO/c1OK8+KoDMc6Q/EqyFVag
Nh4tdEyhc9edTD8Fd2rppxKG27pEITiOXli/sskU8iaSmtk1wzrhtkFVyKE41/3SsBsgZNA3Wrth
9PQjdSnHflJRhEDm+0OqxqdYpu4zxFL/ID3azVsOigJPUSRk3cJp0Thba+voKjRs2NBZNP+q2u5r
iB8ZqvdnD0I2DYASv7hNXGYkeYx9e4P1bLrHxufUGe3ITstbYxFcotRjIBGjC7bCJMMolkk5vwV3
SZFg9mmNvM0H1hW1pnlxWhxooqWpGZ+2u6bs/uuPe0krnsvvKnM6qEwsheVfLlOYRvLNjuMyYnRM
QhxYFndwTRaTEdmeVwOWHEgv92/P5Q3kra5e3Q1ZfByNwO5s/nsbZQsTiyisuwzJzePccLSpEAIE
MjTj5vHFz1664jow/48raFwTYHze4W+7AxUwNHi2tn9oQvXA1Gl/sV383M2kpdLJhoo0xuYDuJtm
ig/042BRVbyOojYqVe2o93THVnd90VJq+w+mHR6bMUcHrp3yfqLHZJiWDw1RC+Wv5X1RbUDgRwXd
Q+eCVV3K17bcC7kIOnTfdLCVLk8bd46V9CNUh97Ro4Y+UYGzlWzANH7ha2FO3l8oaLWPfZHScksu
n3Uuo7SOfPuumojH+N1KduWdayFL/tdYTCYy80+yOnNCVoTWiosuoKD/8FE2yyoNIGMTRX/h4BN8
XtjGcG3slSPZb3CIARPRa0o7Dtp0LvM0XKmVp0cpSCdjnBHJJU3rJ20Llf72vxNWy2tnbe8uAdqh
DEAO1NlFppFwueJwhHGjOgQljvvmJ8nrPIQ2TneCjyx/dYzwUTlTfPfzQEI4He+BT8lfSwJpwrgm
qlW6QTilUVxSG6JsTnDGBznsUpbJrJB4MdXI8+WZTKet9LVWuwE9YpniTrxoaTEnGJQ2rcFga3KB
g3ApU3sMHMRgqo0VHwHsf5cOFfP/TklH06uEKDnopdCBluKyeZx5iyJq1LK+e5AWirjoR2gPuW0j
e5CLO8xjgxJk5oDxcKr68sV0yvcADDxD3WpJXA+BDJCgSluRI6wpe4HeIqNq9SzS2KziwZhyRoFL
YeN1sQXoZIGUAWpkEqIiTpt0eGvtCvvm5kJCxQXk/nqG3pP/W2GAK0IHNBZxdFA09SqYWqC3C/LO
1woEFcGW8Xq7ig4RdmGPsBnwCC/CFFtf+i8GlT2pPhaKWsB5fxi3ODDdqP0ReRstBrmR0VLeqCDL
1yHn24KUpA49dNtx1WTpOveypwBpA1ATNW2jkSa0KmJCyV7TIsf1aVYtzOqygOjx7TaBEj5IP/tV
nwZW1pE3y2Ccb0Y7XupMHDHH0uvpwL/VQkx1mo5xJcWVTZp6M6KDGqU6jN5+yc3Qhn8O1HAogN1B
hEr0A8eyXvXXF3a9Doau6SoRotlspEOB6/afHo49XGAvAxYPOQsBQbSfyemLZ+h10GwYNqfoDjz0
lKhbEPCaYclkocS+GOabjIoIxruCrkRtLucgqz15/fYnDXr2tfFvIcCcUMkwWadDGfWUzZympelL
9wg4J4wHAOpXh/0WrNI4YZt+vWmOA6oLigtW5ykZNXfElkWpAWxsu1+jUosHWoNIU6M9BsenLdzT
P2tR/Ut3Re35n/VEb2HbPQxwdpXUjFuMG1aQyj23/K7D+Yx45q+n4bxdp6KGzq+vT33GjHq0/SYy
QyINfEndq9FGVJbUr+J0X9pQgBe85Om5Sas8OstcAhlV2PobF1BeNNjRKkpCHmqZ07/K0lAHUHUR
QNYCeS+WjLWHBVZknBTSK08T1qo4vYfQ+iypIcBH082rdxhr0Alaqkl1VCt9JmxLmLEIn+JqsxTf
mG5KicTAnBMxsr3yPaKfOkWLbi0WEW8/tAL+s1QTnXalMcbAWXB0lETCWvvyoYT6JIGf05+NuAkL
HhPS2x/LGUDrAtjsCfR6uJJOhWdOKVdNDycXXZGcX0yY923UjpLntk347yRMq2Ed54rBWSt3GFhI
wLOAKftukUliFiq9jR5ZdY+N69JRxPdss1Tj+qsgLyUHRlGC7PUs3P3+A5R7tfv67JUbuXbzKnHf
8yKIQJ/GolgXgrOG1KAU5Ok//p6bXYnJG1EJmDPQB6z8J46dARLm5T+JjUHB1/+ZlecHn3o03YMU
SZJ/A8d4NkEEHS8+Uzd0j/lR+jZn1A6BqUWgoPi0ZFMXhpmfY6h0nqy4978kHmOyIigxdc42Bcly
YUGoTH1ckdQO+HdvzaCQif4y16VYYOLrdbn9H9PoaH/y51wMrHz4uoyfAgli4cQnI99NfzzUaKJQ
0OSjsZ6q3USAvrT6zZXj1FSWwrvH8VqGbvATlelk0vw16QCwi1+QFFX1Tvh+FWRvbnjSFN0gxKFr
yrjMgBZ6iMCeUb/khDVQAe1kBxH499lqqjCokS+pncVcLo/MWGIiEtSDU7bv1cM0Q1ZWH+QAA6RQ
psaQfWQtlZ3rwPBEVADKa3A+I6oqXaNrUu7c/fdSsoPndkHixhHhYaNt6TnxiVXWl+vS9dIe3keq
uquHi8iUKdJ131yv6hg6KvP7DD42bQZSRWNo8iRsWDZyY8LyC/2aV/V1qTxPOgDu4Y+ujbugKdbw
M/TXfjjxEOhhLvIkvDQv+/aQH517vWq7h/m4Pb2qkKyRWNIZ02QWh0OtnbpH70VI7bOGgUpEiKYu
Cwy8HDkQHDkA2pi2ZZ5ERLa3UKkFpWwEceZ8hgJUZUSsFJ9VojZTetXSgG/ILYFGPIcpk0j85Mrx
mYdhXiYc1dRl5v4xT17+SK0PU5p+UnBOunmSGKs19oVwzJKeAwTMi3XEqmtgOlxpS9D2LCLb3coF
UWsj+pUMJkLen9ayTprMv0zcTyD3yjfFk9mDxVAKJgrztSW/K0dJaszipXR28A21xE0JSyB8syEC
89RNYHyuoYsBKHCJD0qPEA8KragfIOzGrkSfz3BHaoCXjpcwxhUhpNHJszOqy8CNrqH378/MIiIZ
u/a3EBNHndPkPkjMLT9I5TUn/odjeAFv7p6Ekz8B5cKxztzeHraxw2Kcn9DEgAga56Z9H3aCiKBD
rF/Sco8nKyi1nqgdKqgdb3mvhSPpruVOccd8NMtvr3Cwr0RmzLYUvAR60O5gneTishoff9LNoMvt
pUzSXepfn+xGT5wSF1cEHMzQf9Vcl7VCeOfakQW+6yN8YieY9Mw5ymrsLTx1pG5hbZK+Hqowx1b0
cYlZovoc2yNb3Udo2erzM0jV9v6jjCVRIRuIKwwyvNdmdOfERkEEya+mm+UhC9YL3NBjaGFjhkMB
nglEjE15bGdEdVRxGCkBTNlZCUgnjFpLll/9QQsE7DIt2qYFpmECmNw2hMH/kxbXvAvG4ggk77sT
P54MpKIzqTO4iWV/KQmaQIoQMwgB8c6nPXn6QyZXx8KEl90Cvj1RoSgkI9Q+EgT/jVsSS5fnspv3
STu873sI1mIOOFF/FSfWp7XvoHK/fsf5j2st0KEQ7dalh/++oNql0xDjcAD8vi5fAEmOyNODr018
K+pLuMviPGlAVrxXm7/urOI0bpmllizNsZXtDd2PBmpZBAmgepJw9helbv6LfDv9dpitjSB/16Cm
fPbcpRvkG3zH1KEs5nknWzSt9l4QxzCIaJdpS61oWMXoRdxd5iVpyXrHP5Fz1XiRRTko6GcLJVau
BzioI/vki1rQiovpYgl3JKR2HqiJmRNlv9ai4LGQ7aEvM6YVgOl6laC9DlCHrvlRt/4q2wS8hZgL
qTi6MCbVGAEJGNuFokn5HYjXpIrDTZ9eI//j2dVeUkc8DtMEdMK30cUTTpWD6L7vYsMLoo8czhnF
7RdAmS+6beMX+zaReNgCiHa2+42FGpjO58GrM1m61Gv8d8CxN65YcXA3cPfpKPP+bYii+MMQzYG7
RVQqTI0fscLEc9+ni2X9x6ZZwsFYLvrz7uPYR1TolxWDSKeU3nA32aC3rs0yuAQ0VasakSD8JN7M
Z40H3ICz71CjDvDD8nk78g5zR7sn3oK5WJGHgDuZo4LFMUvGYS1h8K5DdvRIfxPuomKlMbCAKWQm
frZSitHklgCjgsB1zV/HgZWQOv+kCw52skA+7oNNEZMUTjY+6zLWMOQD9s+7qHUtEGzzmaV8Ews/
Qcw08zS9XCltxvzLnFySBW30zuu4xHbOPOu6nOBEk5jQdG1nSgmtaNWmB89Yre69X2yiiCXp03Q2
Ct/ii/72FMd+eMMdliDIBwpSwm8aovldw67WYcD99xa8a8InlCqq5ehTauNnndLiMSMchP2by6RG
Szgrp698YxYCqDKn7wItUwI0Y6D/3ohxZHIPolvVh3ibMyOJwIguV5l1lvyjBqPvxJCTFG5E8noE
ZftnddfwVKC2BdFFsinPPgj2KrXkq1yS6R1I2fGvZoPkgG308A9ArbGL4exWeugXzXiGk8lMM0BW
6XcidxDfq/X30efqeU5EGWHOhZyChR/Tyld+7xP1s7gNRadkrLNlwYeJWpti94e/SgCKRqsgk81F
vc3CIqnZrLPYx/8E3qZFg1/t9QlRLubL/c9x4T1rcpMrPtqrNoGrFTNi2fdxMXV153R280E1Nn0t
a+7spPOAOexzx3IzR4c2fXZ7M+yuFVpM7GkpA8AszyiDXTYEeDY/kUzkDPENtfsNC5LArPG44iE5
jcvn4IQ9RFIeZHVkS8UADZBqj5RC2AxJpTP48yfYtmbl4I0hE1ewBe77WhtV6L9eWHlfjWwT6mwo
KM5ri5qGwYbU2ADmjf8tzFg7WHDgU5ituZdGYspVsG+oC9niyVKzevPISvA6rcrL4FovPsF0TwC3
ZlTv4vSN1ZjwGF0q66P3WAc/VOb0Jqr8H9v5fNR6WaHNAIzV41bhx7OSGa6ciHJ9EzK9/v+pnbYS
hAQMYWGcx+k3ez6MRETzZ2pf0tRxDxHF861aXZjo3yUZUBI1WZHoLip34z6FeVypoIIrTXVt8uXp
4zHxQgEUAAyXhJe/6HzYBojD2hvekwamIjRnyGEgYKaOImNlIGPgEfxiaooSj48odq8RadQB5baa
qqoMIE1qPROAdJhFumDX0eUTz7sjGK07kIb6wEYVuENkzEsBU98W1lPVNriTnwRmmY/dbCcPVIj2
tjq1oJ9yH/XLhDXNUGvCTS6b1fBEeBYsZFYt+xbOjfpeQN7YMb7YaYRnIuC2+pqyl4AgmpwYjW6d
Dn32oV3Bl6bW3MtcwVxeGifanGutLHSnrq5AdgUTIOph67yxC/H6sN8FXlPuDtoM87WkrQn2kNXO
Epdxqf4Bi5jiaGwxzD5DES/m8EbPn/bxjJpTE2ppoqFeA2f1xDagWxaTt1d/66O7afKB/FHFyD7P
EMLgzpO3qohZAt3axTKToV6iLuK5XUn/U4MUY64zR4DMGPtmeQV+NZijYBdDkJPkPY5oyHG3kBSA
VNSEuD3qLXP9gQ6xmfZQUfixWbnc2/Z77It02KDUzzWdQTV04SSiv72ErWSjkdLkXWId3jupT9ji
g9PD32FSR6TuU/4PJnctPTBy44hbZtAmZcO3m9CWfmHC2DaS8SOBYSumiHH/CokcfVkJguhyEUSt
bhUbiYK1g6KFJ8Y+EELlXjqgTp9xDNYwAxo2KbGpEqTXd2QlHGCzqiw7m3mU0TAJI8y9awhfIoup
d91hfhq2C7wynRo2Ezf+QZIJyLLuz/SIfJ3Ms3BEiFL2OWQlYtC3PwTMyypIQ6EoNpBdwrjZHlPk
CqMrx6teszWlkshsFFtD+96xShirdK5lVzmVOhlGecF253096QuryHlvqE4kSj6peN2FloS6xC+6
2BKem2ftarfKFPlmYDxmUGZ+zFNW/SGun8NSwYCb4nHw9VutfjilUPdpBEJK8Ynxe5GiDDpPy0pb
RPFloq8jSBVCIaAw8kXLqELhsCJo5Fqnf7gu8V69d3eu0UKBL9DbKyJWjtagWCM1nJGSZnN0lm3Y
5AsasTHsPtu+qis/LuRsgbZIcPafRySgq7xTfr4GG7b3sKY5B0mCKs24MagZRyhlSCMF2pL8nv7T
45h3KbHcCe9o6ZhqJix+oUPdS76KAAFmWqu6NtyC5SEsHnoL/wcyRBmvrxwJX7xRpTE6oMW7HCXU
Eh0663m+GtlJL/4YGGACjLGRU38X87Ew3FISLjqbyyxj5I1omKdj25SjdWORnuQaOnHu271QfY0D
ltfj4YHpwSxBUltCQ090/6yDrCOGPPjJKINgBM4y7U8lxKys334pt7zjE983L71PAOe9ueLkcLEr
Rc792BXX6SD3d0MzjLzWFgvT70m1ZTPCqRKkPbAM8Bcq4Jf6mSey6Wh0PV1jTe20WusUr1s7LHdl
j8DhzRW0aCD4Rcc2JjCR4sAM02mUCnOx8ZLxuIaOC/BEiChF2W7uUzgT1vY4Xo5sUEJMktnLb2iE
aahSkJWdJUKdunc1tgpf5eU8iRBQxrXmow7VfoWh8GiKbWQxUho3FLH91so3Nj2OovHysIP2JSKo
FnFI8gYelp1qU3Mqgv5VN4lFFAthLPmIaZfz+xhzpIS2wAWEviBSQYT8gDykYP2ZpoZ1tGQwPFv6
qHooX05gDS1P/pYQkV62AuocsmtIuIa8P2uMUurPsNuqV0vqpsmzuEN2tlS1KplVy7SV7TbzC5JM
cMeQ+FOIHZaEWcDvQduW83GH4v+S/SwT3mRoNF069vPa9Crvr8qeYIQF5ac4AQv5O4k0tMXA6/l0
mMv6T9g6RKjQ3r1NxG6lUBAofPdn4wQo9qJ864B4Zsx9yYVjlUg2YcTs74F0Zr9vUpGpwtNMb1YK
e/L2LlZx/+WiuvdfhvgQrbRpDq+H3YNZb/x7vvMKjPzssiJmFQ+TblvJJhMAZiusJ+z4dLtQMOxi
wzdPJi6XSL+GlgvTcjATGjbqzVGZ+upwmDHE5m4IKeRFeUiSnjPbJ6xod6f4kYh3xq0mBTuBQaTe
/WeCYL+Yy+lhbcGlQVv7l74qTl/sKPr9IoygGZCIJ90sa6tBCEEiPd/EEt5817oWtkYn3F4MCK+w
4j1so5pCG/9K3enMsGaMtK/0CYYEQ0K7j82H9fLWxBGc71Hyq1fY7CxqemW0INbhcc13QFo8u9+j
QHRJpQP+V4v/ZIcwpafedB9c3tUffvXWRConCiQjXu+FzuitBQkELJGlbvoQF+3A8D9KtwJ0KxYp
3mZb33KPZt2pVNF4/eIB4EwCNTV2//6p4fSebCJ8Tr8CsJs+lKybbT8OYz+M0fxr+nmjBPbcifLC
ydhD2Fqf1i89KJRCYtIBDw2uoue3FRzT3nSrB/A5o0qboenY4QcP7hZHBLk9IVJ8q1Q5dfztILLj
/LLcyWRsF+nadv03vB0fV7RrKbIUEcMDPUroN0rBoGnR4OplugNHttshIEPBx6j1/fEVbA4F2Gw0
HfPBTxLSiIiodq0kH5QBaTQpgBy6ixve+wDf1UyTB6R9sEZjdyV8zE1YSBieN54NZRY/FStgD4HI
OmZORNqkEoy/szUd7Tk1YTro9gIieqtkvROKlKuwjdpLqF2186y+AtNMETomPlJEIg38cncaWQ1H
MeTbbmNBD2ULOUKFwwjXQsUJ2NlfzLdeYH4WeVVyXNJnAQS3aSEVdqAskMs1TZbzFOz2OpwqU3sb
8n0bMB/FnHeMBZBpRN1DRqRazKI9+NJg1oMEf3diUcV++/IyrUQkLWZ6GTNbRGyiCO4LVIT14mbG
nyk+uoglZaXKeMePsojJtYX8noKBkaWnT3SBB2qFso9FySiW34dWCPTpvThzj9YHsvS8wvcbG0Hk
tVMpgamp2YjO/AtxHE9S/Ql8X5eVZCa/8ItDJIJXEREsQF4RQAFmZDBA37/BfnzuydTQ+Tg7QtaF
OtwRIwXGA2ORO4vP0iiNPrpHheK6YgsM6OydT9br/B6NnZFV+7wpARZqHeWXg8l2jsA3hSilgFBW
EbQTQhnULDJFw/zzbgEfB9s+Z2TG0Y8R93JKGSzXHHKRgUki0AxV1BaGayu1WrD/1bMP54YbgaeQ
SVTvOGs0CyW1xoZ+EngIX3Gmwtx4bHPVHpAg9ctUt2M+KV/CzYgY7LLdWB2CAcIvpf6IJEnacf1z
qMmd1CUkwnBR20QSfcmQj5gohdWNiiAy7ndtzlqyhUgqujWTcF99jc4gbKa9btslsjYdsr2pEhQp
59TnMyu33GVBKQa+qj+to/rVu7XPJrG4p+Ovt/nTuLX0Ga0=
`pragma protect end_protected
