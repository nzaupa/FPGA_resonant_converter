��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`ww�	�Tز� �=Z�ApP�>,��5#��T�]7������}�z+�1�h�ː*�<��o瑭�C6V��L���OTm�6�~'�c߫Sҧ@V��KH@����ĚZ�җ�c�b�Dv�ɑ�u�:���
֍��O� ��N���8�Df� x��������=��J�哔��ԟ��l�_���gN� �"I��:Ӷ�>_>�6h[AU��P�iYo�<3���gj!�+E��sʳ�2��4����/F����~�\�)��䢺[G0/��f���0�P/g�'�AU��Ƙ*�+V���1P�g��	�mC)å�r�<�H���c��"��Մv�-9��^�'��[(�����XVӐ���/���4j��1
�6j�����U[�i��r���Жn���4J��AE�=��Ύ7� UL��Q��1�r��8
�L���i`�����g3U���Υ��u;����������4��*������1��C��a?$d�qh��sϢ����5H�����ضl�PO�E
���{�+[��R��V��f����9���$(@�J.�����^]�Ns.�����JW��e��MY��4ֵ�O�}��ʳ�E�WɔR�y��nx�d�����3}��X�~���) [�ȳ7/1�v��2C��E�qU����P�*���썵T�c@�~���w5�pO>�I�ݣ��-H�1a�<��sj�c"��MX�4�A|t�E6^�	4�b�O2���bL`B�I����n��F�ݙ���ξ�u���5�� ��Q�7�׬�5���^Q�I^��2_%�E��St���K*l9�W�r���;��j��2T�zT�j9k�!9Q��'\P�H�Y����Ǆ�	��ۏP;V����MJ�>O>G:��K(��CdE��up�9U�����$H	�� 5���.� ��Og�C�����Fs�0/�h�\ٕ�QI���S��u5�R/�TU�����[���j����3�q-Z1�:2����T&����+�/�R�<��:#;�B��g/�	�j��k80�SeH1rJ|IPq�����N�lI���E:Q�L�I�ox<2��?�v�侲�閜�XɒZQM~Q�
�e������.���Um�[��M%�i�{���OC;aڻv���[��\7�q��2�ɖyw@n,F�+U�|��mj�T�b��ۑ]���P��w��)(�Qz�Tc�@���U	�����L���o�3�I�iq��3�џ\�k���Rr�3;О�)g�)��t�#搄��IȊ��HJ#�M	�ߑ�2dT����z���	��حR�5�@3򥖵6���� 9�3�q^ci���C�a�E���.�9�gu<��n��lx�!6�H�RF�>���2+wN���h�����pT�O�V��� �S�٩��%��B#;���)<@{�j6��i�b������I�MMR��`��->W�f7M���W�y�2A��Ȣ�bD5W�L�1��Z�sdd<��F6qu�ki�~�D���G��8Oc�*�݀�ؖ4��V��"��Zm"��J�07+�M<�4k��_��l���˥�p�~��#��%۸�{'C8FR=���8���٩c����΋ǃ�+��IѸ�&D3�zQΉ��FcO��O��������(�z��oB�O3�6n�n�M�`�0�IErlE:Or�`KCVKU���b��Eo!��Kr��ϥM����0���E.$�:��-q	�5������8T��
�_�5ꄎܰ��6!vQ�-Q\1H�M�Mu�-�bT���w�A%��.����CC�[��OY�nXF�7����H�ɿ��/֜�<���B��U�6!��1z������u�qS�&ۮ�ߏ���K��Iģ2�6�/�/I�#�JcH���[��(�I)����M�����lmZ�h�O�t�Mvk�K�2�* ۯ�x\��ܗ�&Ί�%Z�
֝$,���7���rnVZG5D��F�q~Q�V��?π8���q�G���s���d��Q����ML��ŚnT�5H���hE�?ڙ� YAܰ���ʦ�m����i�=���DX��?6�kB�;�8h��f��S��%�7NL���:�Q���B��Z����@2���tlE����{t[�]b1q�1��Z�!G`��]�T��.Uif���X��3��t�s�
h9�G��J�V�(Y�%=���L/��P��������-&%�~w��2UǦZ���Y�6��f��(�T@fW�#l�.4:Ñpj,���s���R�ߵ_�Ʀ����hK��O�z �Wڃ`Ȝg�DwP 0(�V�2�Ȗ)n�~)�s=����I�Y�����H/�Թ�M�\�W��Ӫ�ҵ�[����jv>ٍL{��A��;{X��3{M�~�&O'�4��0��3���@Ԙ7�dso��W�_t*�U�/+4ا��wE�i_���D<V�����\�5_��vx�T�H�� ��l���x�#�=���(�-���#W���vK,��Oϭi�q��[�p���h��ӹE\�: �*�$���R������u�W�U�.m�r�S��/!A�ٰ%[�u[+L���%��X����i�;�4ɗB3��zS�ǀ���o6 O�Z�
����:�ߣ�;��_� F�(&n(=��t��n���5�$̀�]�dO
�𑾽$K=께�z�Y�Q�f�h���uA��V �t�%̺�.;����O�++�"�ž.]ۘT����؈ �~���%�}>h����b��sn�>�Z\s]}f�܍%�f}������X�V��zկ���݀��OD	�~ $�P4��u��bԝ����5U�a�@N�-�,@�����4?\��� ��pm����J��C�� �Y]]i�r���fNP�,���Ⅵ�e�C"]p��;�K�D8*ܱ�Ī'�F��6R1�o,?��,�ڙ-9��-�� �-���ߔ��PQ�=��t���ͬ�њk䚐�,��� /Ő;Z6��Z��	�X=$C�]_�q����Pk�Y��<�fnػ�v���0S��#�O&m�Ct��Ӯg���o�S�1����R8�CÀŀO��˛�y�fẇ��8fgH(\t�W?J��bX
�F������6���Qd�6�=�k��w����-�1��h!�ܨުY$��H��Qh��	T	 o�[�o6?M�4s}�?}�����'"r�Xi���LX���Vp��!+@*)7�g�T���i�Sv��ϔ�g��������9�c�r���^D�����a}���{��v������&=�c�>t�W���н�'�ַ���s(��]�����l��䩟r��c�뿳+���	S��qg�i�v�e�N�2�@]8��ȷ�8�p ��D��Α,�J��'h���Z;���l�-P��Y�l�W&X���%�Md%ٵ'���G��
0L���M��L�|����m"�ZI�g֠;j�J�F��6n~o�N�ʗ�D��48&�+ٗ3D���TRl`��	-<������#c��"�����px���_��*�+e�G)�#���N�'��a���Km�9�0��?��쐕����IJdݯ؍�q������ݥH$���-d�Q�٤�|�������V��Я�ʜ�!�G�^�µP �E�B�nT��P� ���n�;�L;��k�����	C	o�@[+װ���A�0���̦��ɨbD��܄Y��b����A�S^��' �jU���FD<P��}C��ֱ;�O��'Y;��>-:=�I�A����
��]>�I����q7HEf��g���2NP�,�a�2.����z��ò���"�B��텸����d�O��e���n�E�6�*�'�"a{������(�?rq>h�z����+w�+�4��g)>�S�՛ Qv�п�k�`�bZfF�E#�~K�X��]�M��rHE�����c)ޡ^�J��.a��Q<�O )^�$�cK�|T���Ү�?�^�� ~T��`l^QЁ�헙�Қ�y�\i��L;ӆ+�h1���Y�o )���|5�y�V6k:�s��	9�*�;�c�Xz�7B��Z3�7�e�Q�.*��>r -���ف1�]8���������={Ҥ	�W� �o7�,
��(�e��,1��C�~7I���6�c���uj߀B�,E�{k���O|��3\��pf�g�p��9|��u��ʻ��4a�c�Jy�[c��͍h��]X��<e����0��(��(�ow�(�e��T�VA.��n��[W�Uw��_AbɢI����i�:>�֣Л�Z��t{�kR�e	�չ��Y��-=c|u��ڷ1p��%.����B=�"���R�/����pu'�1�m"���-�0;�?��	�}����Z���d��f>�����|����5
� ]$FzW>� �Ծ_3������[N��+�<d�MHf��w]ʐ��񝖵�/o��F�,��hr�JiN��aw�z�!d��u��G�4Ա�i!v��6�&<��g��<�RH3��+�$ǗeN��UUct�����0�V{������y���
6��P>Y�6'�U��|'�[�9N-RC�Q�kt0 ���f�C;�V�kc�P��|��R��OE�������b���{M������e����`n�&�`��>�<'��4r�P����K�V�2���6��O�qm2Uu�"3�U}/)�_��A �j1��Fp�O3Kl�GY_�i� d&0"�N�ꪼ�5)�ɰ$��@7�"�yԠC�X��"�T��,"�Y ���%�`��'���f&��U�[���J	9�$�b�O<�/lH?��u�{�W�ʗ,�Փ��+n�sV�e�n�0N*�ܪ-5*�sY�xj�$K:g�⸣��`�4�_���6>vX�����s|��\K�sƦ����1He�cd���^ı�}~�KN�k.^���n��jg6 � _��,x����B)���k���&)�����Ұ�ǚG��P���o�RJg�O?2Pg�� �,��o0�*�+��11x/3h�1~�sq��vޭ�d�c�!��e�}�X��V0A{�ҧT�4ݮL+f_����9����8tR�ny���r19z@=���z/� ~ֿ�g[�X�+��(�u7[�ʅanLG�O�7%<P��1W��ۊ���-{x��R3���S� )�c$���w�Go�
7��=�\!����z$�x��M!=s��	E9j\�6(��K�HY��v� p��S��4�H+�>*��ڄ��j���q�����*b���"=�z���rx�j����p�.k�o�������vԺ�ڷZ���4�8(�{>����\N��tc�J ym'�w��y�<5�4.�:D���k�zD�k8�����Xv)s��>����"cSݖ��@ߙ�ӽ���,���'��s������H�z��hz�%����&!ZY��۱������Ĕ�q�hx@;Т�2��K�`��@��D���z\N����y�7���n�a�!e�p��%(g&��9t�~��{Y%uP��,�d�޳��Z	(U��U] ��î�kJd.���ޘ�C,UjǬG�^l�����PO�NDx�9,��D*�f���U�� .<�\��4�є�&��ǉ|�u�N��H��k���� >v
�m��㻆t�px��~!��Q���"�;`�\5f���¢+u�3���u$��}��2JWR$�6���\�PW�D���u�l)���S*�������G�ҽ̻*4�T���TN�D냸��k����skػ/��\�.��Y�n˒ZL�9��uX0��bJA�C�T��_t����C�#>�f_�������>J�op�H��Y>�����5�UO,��Z�"�1��O���{��8�b�\q�^��mt*�fbE?q�
�F�U�������~:n��~ �5��Mn�4���07%2t���
}*�Ě5��º�ۮ��?�"�6n$U������� ��5��g��|�o���I^S�{�tO���QN���eL���1���2h=x
:I���j�w_�����A����JpR��N�=Ռ(P�gcr��('�i:�\^����ba�7�O�Q�m��c�ެ�l[ 9�[2(I4OA�kiZ�����hP��m#,Y&�#�َ�8���f�����S��	2�e�_��>��N�_i��_�n8��y�������O�E�}_��-'BW�EdP%<���*��.s%�V#%kП��Ty���gE�	o�2*��7���ca�h��}@ȟ*VTD4�38O