// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
T/qw3vXNFAn9TQPN5urIB5RN3RdvLTk3y8RW3YK4HYQLFdtBQ4Le8DL5eGLi6P/ZryZHw7r1wb4s
T0/q/AZW+ZViXQTxiWdz57taJJTW+jk/bOiwFU94aQDvtphRnU1+NPHHl8NUx6G2R1E0Umzj++w2
R50/36JeyWEsbmCzLx2FNi8lqUadRaCul+F/azXS4NK2pv93BuF20yO87TwHaVaVTQ8PJxBoLizN
wivpZVUE0hyxuH77aHvwMA3HBO/cYJSjWX5Mb1/xSq8luhAp0slwcafNnIdh/FZNNJZADqlRrV7B
YdM0w+i528ycgotkcw3eH7BM+nOFknvtsZcyKw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24432)
prQJDoMLkXNVL3QhcWN7oVxkfoMW3MzAm5lhtpbBEiZ33rWgIdyKjHBFDR5kJYROjepN6cqlaY9I
5tLrLdMCMdrCCMlRkPt14P3DY/ml9orCaK8A793wmqtoG6yMVDIuKzbPmz+yVnNmg3J/obpNUSD9
ay42dw2RdAJsQG6VJ612mHLEeadgg9JA00o5CsVCSc6vVLCjLxNQgP26HEs1grHVxW9NK3/d8GOf
iLFXZ8CZuQDZeZQmOZzxnG1ptq+2sfW+2gGWAuXkt5lbk2vchlgVasd/1zI5hbMoqzAONEQXWhya
hygxPnnYaO63kjfY2Z2QD7JDsxHxonkY454CO2UCBFQPIKmZuhD1HfOuOOEHzWzZGRMyPnqKALqc
IhGbxj+H9ZDt6CpwS3WlgVIT+h1VV4sonNTJIHDG693T8mx5UO3sJkxGmEVHArV+kWK4F9O8qlmu
hBE9EBTVLbGExujoynuzjPCeqSyZPoWAgWlTc/1m3dujbpFmJED/PefhPw6GEExPm+W/YUSqM4OU
GcM3GPi5HTmpTylVN6f4pHWTuVr9tOh+pzSsD5ImAge01ZxfEGKiimXRLgGg38fqE3vVH3ibejB4
TAPpFSDfHkZHF2SQgXy7SV35g0W+KYKQPqO0gY0886855e1i55Jtf30CUcLGxbiiESIeVlHJModp
zYi/tVdidjfMstFsF0N8lGVOQStfCUQeQncS/ITPrRbsapCyR+HmVZ4nWKE68MEpSol6W/gN/BHP
FWabwpsiYJ0bJi/jmuDqwZtLeCt+AcQwLSWOiMKCNZ+Vmv3qQryu1fe/9UfBKK5hxj79PfyT1gus
r3qKI9qX4mu0oYLn1fEYUSs4W6EWFkTKDzObzfW0DVEiaMyOwNTmnyLTwCSUVmvKHjqsqxaA9CMZ
/yoWY/uxn4J+uJ11bzHvRoDVhGSh2J/DlSk9L+d2x7sD/izODMw2V6R/cTPKPXQVDQ5772SgdAyP
V5IEXeJoDx0pAbxz0KmB0871B5d6py16GHieH9mAH4Abtli/GTVQ6JlaEs9cgCEmOvByzZJ6uEDH
eibomdDU4eUxtwYrzM0w2yDptrHGDQXBE8G3VZVzTyJwZ17nihICkxEcCegxSCwv5xMGn13fdL4z
vPRuVpMBHlJcOEmj/EzCR/isoFqCjAFhJ2iUwlT5U+Y6gR1/sKtf9kMHWeujJ7Da+5KoA99CtEza
b8Fp4DJxN1hEgo0oVBQALKxba8JbuD07dlDl4lLDCH9I3yJdTNRyBX1eB9McBM/qCF7sbwZJJmrk
wWK6W9Ry5shnYwFeys7Qu33rHG0LIYbl9Balyf8m/9z2vt6ROt/JI8MBGKciP+RHt+3GduiZuvGq
MKI5dHt//GCrB52xZn6dl3SegP4dU6ik+iSmyd7UZXTQE6FNNmtOSUkvzeiXLONSdTNRuxkiDQLK
nBODi5C7tadozbhRmYYHcJR7K5EspBVCGe9gHzzcYRtPcfBIvZLqHnRuginCLKVj5axyxYyK4eZT
ClJgPTDg/Ux8SA1QDi8MChZRT+Bg+bMyAdktPFzi1uuMIEzSmzf4NFAdPnmU5UHQh7ZIhw6ZTgLj
nhCWn/ABotaWRXaO0WiswOXdLe6nnnPnsy3WAl1Z6BSQkfXSD9HtEQAqdF7dBSAJzV3VGEpKxhrj
t5lQtM9ZYYD3onrVEWpUv2CdoHZUfNcnMG5qWrVA3MbsK1AknNI6hd+gXlD+YXMytPuTunXdpFcu
xeV/M9myvwiNpqdSLfc/3MMqDVyIN8r87RJjw0PyUzX6iBAAyW6JD/WEgN3+NJW1w/a/x6erTFPl
BXK5q2abWQMUnTWrIGUQxLxn77poBNw/IWEYLfAzRCAYN3qrUqP9jM4+aF02ArpqzLWSW5Tsrbvb
mPHiyMoRyB86m9mC6GH4Z0aP1Hnc9sGeidVs9kG5WBBxGttYiaAcBL6J6u6MCUKwX8Iwe4scUFkZ
wmOSaK6u/iW4mSRNLUfoC3ylEG96+p6P9ZauJBLT2EzFWQB/YMVGxB5I3+tPODeMTleF+nNqNVco
AFW5YCqu01dv2QVGWeQ68DHSmayzvq3rjKp73YcfkN4s43tWwkmKD9p74AvqaW4/WEnTgOUX+CB/
bULK/906CJZhpqpnS/+p0jSI/HfHylRpe6O0bx/j7ZQGGM32n1g4w/cxSBZclUTIN3kdhn/MK9KU
FEy4oyTjNbeiUdC/avmwPReNWKrO9D0AickbVVGqj7YlgC2rwY2eQ52y8OyyBUtU8/klpssmgi9E
B606luam8knwdX91rbqbTl/oDEmb6yP/6hCLjVJASWXEksznlRy/Rhm64pwGvJizQYBVxQS+55S0
insTiBXB+Da6D7QMmO02uF8fEc3aQWylIddV1ipy26LkXm8MFe+ZfzTIbnHGbY8fRH43ZvYQKIj1
7SJmWmvRYJT4Iax9N35HgS5PHP0hGGQzrpJiYqY1UBzXETttog3AVfKO53bLiMZELVaDbeXsusdt
ZXcUbzXIL3/a4+orB75PULXffo1iUiixa07pdm9hS7RgsIaYJG5zWc3P7QhSVGKlXGL24oVHKXiP
4cy73nw2IbdRIngyva2vU1vaZlQkfnBOrnnh8EIC/aUcp8M1pKU4VoK/D2eSHXRrhMbT98l+SK/9
pAG4D/uXhM+l6E5pqbdeZ/q2T3sKQCwitQyYX95e9VqGS5PTBNkK5Ry7TPNwdl3AcZD0xCjXWs3I
yj4lb+1uqVn5x5pWACWzxjAtmJYOm7tye6rGwrbWluxBhf/GP8aKzhy8b+tMgrrZWb7GWtm97i2m
a5YFKCvIA61NRhHLm+pxZypP05eioV4zdf/pCPbjx13+8QEW4UoSKbWV5IP0/+1etA2bVJzH8f3h
UG2g57T2hgtrEQVu3PNYbadsJS9PXYMAT3FU299txh/DEOPq2x9opBeX1NUhQpA2hIjU5ZQk63QB
S2/YHEr1UvLM/7kdnWz4yyk/FVUp2suUbJnCiqbabs4lXWgqBZgch8nEe3hVVUB/VCn8yt7sgomg
atPSPSdXysovwepKgUZNbVy/GabU4ZPKhrJe/7DXkGmcHHzTfwBEUOZQKlc7oYMW/ESIM09Ral0i
6U3HNEx07lOrVZb4KGpiIl/6uAEwXZA5rqhKCeWbA+d5P/3JL3Rum/FPTKBCMDPSZzC7QQLjWuyH
mOxXRu8IXrCESHEGUs8aCsNaP0lOaSUUsrJn8NDKTFOtLaRYIgYNt3OZq4dmWXVbEhQRJy3aCF48
Gs9JxYtecZv7i8lA0Q8eEcjzwVHeutK8EgRxf8CBK1cMSPSStYlJXik7iefMa3qjJMXbKDz4Vah5
kCwsqqp51uSGzkVnq7+EMuNENHZfeltGOVar5NwfTk0bVEQBXsOgdeEdLhD+1TEtWl451GX4TEVh
wHLzowHIqsEdTKjWzQFayZhJ2ZKkuuOP+cB0GMQXCxFo9v5vs7z66smuiP4GgqcunH12hdZe9WUl
6+VeY6IK7FN5VcKRN6GgcwrlHtmmw4LscBLvrnrWc3TjJtFrZ4abBYsXNc7l2XsWQQMKqsN2pDkK
OPssRl9qSPniBDR5WYFS/5fG0DUH74l0M2KhPT80dTIPzQpdZzLFZWo+jUZhMU44+3yNLZvT0iR9
DkAf+kvgheHMbS4ZETBWIxhKpuHFYC3mJHCtpyrznssBHaUCimLMXvatx078kT6zPEx67BW8VajX
CLh24chjkZ3PTEawRczn8CK8k7HPHgYZEDtU7/OGU4gWNOqCIjDIrmojT5+u/MLy4kjnMVsMlQ+O
XRAdrP1JKNflLov9ZLAd2ZyVCtOlPeBY7NU8fa+mjbalr+y2OsiiHB42OufpeBnPuaIFp6vfcFep
s3qbTQjUzd7SaOL3rRhDK2S8LsLcvPP5bh8oqXkrFovG0srFMhs2AdkqZ6ZBD9NWAq8Vt2qCyvEd
nNQUgPOQ9PaOp21UrcWH0xhJSZMgrubMcXcNHH8Cn7QSybEjxULdKCUspdEFduqFzhSuGukd28sR
X8UtW8OHamQHPnKuyq/YTTGdydS88KZUdSbLw8TYBHR0R3FtLzoFxtlRFUkic6pT1keslWdtCIHV
I7pGmpKK5KYt9oUurb/dlAl7sugXxOr5E5LUOK9Ca+BsaL+yD6RH5agigK8gpICLm7kPYW5Ne0iP
Zj1JVhRR7+HbS8a4YFQj8anE+0joHKPK/8VyHyvglWS3ohSw5FaMVTKy0J4VXSbUbR0dw/Zb0y2e
zlQKB8s8InuFhYHNuXHCiRmXbXLmvWMWXcWiua3AXhHUPJeRtCQIjpPTgfsSH2RX0hXUk9E+4OtL
96cU7G3nGbOSq4ymm9vELF3F72UJ6fSTGJ4GjH4dMS2o3mrl4PWKW/AQ3FGSsb1mebEtiQEGyBtQ
+pg49s+Mx3QChmfMu58cksTTvbvbrOFx/2YUuNpVbr2CtMdntJcFJB/dIotRJDsE3aNj6kZxDgez
kHIsmEAA7LUzGcuQ0/1xZ+RSL+Ix0uhdenvTdG2c+OE0WGFpL/G/xjPAFUjiEmfepvDIt/dy/3fx
hAqOM6vl3sy9BQxOi/d4gqrCECoKzQrED42XNyeseXZzcSRJz6hVTPKu4SbGBRxEreEVt48yjInV
f3ewYTxJeQwopYtiA+N/UZj71CzKwojdb7kz4AqBB2aCUnOcWbgHAwvCXIP6HwQH8kHJBLFYDzuE
XALYXppAx7pzn/qjy1+A5KVqsc6m7fvTBRHxI5LCIvi66h7bxG53L35DG7UlwRUG2qdUaogqAaNw
C30kgkTjHpMwfVfTpF4mDlvSXZMPCiq7q2VkD82/QCK2BxDReyB3MMF/foz5FI53bnhtb2c0Ajj0
332Vl76xOR1CXrZpAuFgdlvAkfrpg/i4coVf4+fowyQLiMU5FVfxmE8RmKkahMWGr6/VRLsdGhPb
cgAVGSTcgU31iXToertdexLItrVOjBkmh3atvDcKsUxBX+uBkTv0TWcarbTRj/WPYujNmFMJ+2OE
Vsts2F+XaNLO2Uw2fboXXJWPkVeYPe+07P7FgQYNNBgqvCYyoBXp18d2OeCjMfE92LLqQg0rzvAa
KHyXz4dcJIw38Yzcy7EhMbtMkxZTV8Mbm11Nj3aXX5suGAd4s10aLwPVE81E37y+SFjBRwnelBB/
IbQIBycg960YlKl3m7SN222rVZq7PilvKdAaHf6YLDkOdFDz8brKbqIgNJBmXzzf+uCGG9msIyAK
zalHPzwQZCvRvYFUrTl7C3FrCazSlWFbZP4cB/qbKGaN8G1srXS/S8mux6DMHDKExU0vkB66YYL9
pJ7yZyFlDMtIMndNi2kDTnaE9D6CmB62E7pl6ij3t0LbSuV5bdtY+CNLxQcAuAKZmIzOCaIAvYfh
STc2rlj4ilDqSzievM4jC2xViliao59boDw9wqkuApjBGwIbnJBChVVfdvpSKQRvJHwk71TTUW7w
bFdPoi1cYEmiOECqydbLV84zT2XtgF0DzkZryu8Y5IL1Gkoe4qxEZgFvnVma3zasqAAJ3DToxa2A
zDrltLXnztyAut1tQo63OVfyAlZbQw1BRA0Dcd9OYc38UhQ2n8qFDtBHiJgkj6KUWsxCCxt2LohO
JYYI0phfl1NFHSQREbm7WQEFIY7SrG3jHppZ4evlMzf6qeKEKlLR81t3n11kOSFXKFNPywgMBfWg
OUER/2biQODUqGMwMW9t9lTTqLcdEZOtjSlbPvoWAKbgF/dGrBFXDY/Bor3XDIPydP8EBeTiugkm
9LLjqTnmTFDks/CiSqSjUcwCKanutVEYL2Vb0v/+3MYIeah7yNw0mrX7JFUQLhjQ41wns2P3XADw
B33Gku0m5xJI1Gr84xUevFlBW7LEX/rVNu9zc3tZvVMIHYtjwvvlJ7wpdIOAlB8cZ4kaJz/7liDF
ol/YmoNZnepL272HTuIUHABr6cC2A7/hjkVpgd/vjecCm7Kfb5wda3ERCBEgfNIfj9rD1eUmjoiD
eHWhdnbFDUGtOi7wDCT9lQ4NVB4hiUWNHaIsVuHOGSRAueViTN52k9TbuI6f2zgNTXN3qHiNmTp/
xJqciq6/tW73v4CbLKZzr2PiUZ55acojRMJ5K3savM4JV7kRNBfZ7dS0ed3N1oTUjvIQ4YnSboQd
XVPsSYXzFL4n1OmxgN0ya04gu/tU8QNMdO8swqre1YQciw/VTBkM8AOPE+2f+T05waD5OX+6/Clm
SAe80x4fbhtHa6OtAyAP2+67jycamtiPcbCBepPIVzLxwWE81TFjIN+gTszPCiA0dqJItBoXYKFx
gap72hFVxcVETME9xl0l0rEILdQjKxvZ1uqOk3nopfQIq9zfAvblgm1NKljKvDaLqUpt/Rc7UHWo
lgwbbEIt3kg8fXOiW5w1ZBeqGNZ9qu45KMaWpYefqwunNcV0sq53QlxTY9iLYp9SyWNbDJ+X2cs8
sScLHWHQHCjg4/YDP4X9oqOSJ9suYo820SiSqZ09gdmhi4bE/ztnifQWdjTQVu76VWL6umI1JPCF
mL6aUfdchVN16MTYx78gZIWcYSBPorFh+3YdQ4GoC+wf4n4FSTSz71vVk2aSbOXvmkgYu+cgLCuz
fnnx+ES2Js43fmv3PRAKBhmtD28hevR7eGXbLlI0U7tCaQUushg/cG0mg+h/E12G8So20Kh/aJk+
EZqt7IvGGsaKLrx+VGaa5+p41dVHS2kA/EGO84+FbjCkQghx5aKApBPYpGeY+4QfKCWD7aknzxwo
PRTmcCe5n+305P1v9QWRrp3DyKU1D61ajyRTsnvUZCIC0kD7k7+CRXWxLvwq4RfiBK8YRPWyUmdS
gkDv9XXjJUg1wUMm0YW1lIj433blPRQqRmajqr5oa8uthvD66X3iEK9t/Dzb3v4swrKX0ugCv/qM
9H4Ypi0fpLdCgqPchEFfrzHVq48CatxATCqvghDS01gphhBtmOJvKtkvXBROYQdHcpRaO+hPq1kt
hCssvQjTmWkI4mrmAcu820VyfKn/O8AOverER+DvV7E3O6qgWnjAAZVpBjapeMue1mxVYMCdCABd
qMhh8W8A+MCRp7Ze25PIIeC67/aNDi/3sCLCsVOP0WH32stmNrO9rP9C84Z9SRxwRICRUoY8axEH
k30+zfAARHvwQuAM4DLHumSGvS23A8mqToJo+7mT2L4RxWUKhiyXOzjWkoJNdbV/ZvmIS6f+P2PG
ErJ8/hhaRbcNywEHgIY3u2fzgiUCADryOg09WYxNQsMi3YpTx91MVgeJYYpNBwMBlfqxrZzyAHDu
X9G0cCjcismdi1ksGlPWLvFr3Dou+sSuDHXs4usael1eECec23Q65LRYNZbW8BdbxaCT6+Xbx4Gg
yrI3hdn9p2FlUp2kBIW6xFtvUChrY2BPJlGm6SqDs0Zl8hhrImUrt28YH5UeZjRcpiydFwx3sPLq
jg9RQlkEnQ9yQg1gHji2bVIZ9cxVKOQ5lc/BLJXDHhCgwNVK+w2hbpHNKp4XB9jokQWySO0Ue1KE
DqRCzUhQTltwRKCSuKi5sruRhgnOdKmjwCYdPJ6Hm90d+gBtTq2Rnkm9Usvsfw8C23yjRnIczbj8
EPiQfEPSf8Glwo2no1bv6zgorsc5+3nNQsxhHStgielacFEhnvwLEwZOoYcA5QWAh8ilT0hWpvH7
3d3RY91b8VOBXR1qz+1tQAMo9iEiZ/cYv+5gj4WPah8UHS/cfgS5tpjbsb9Va3LO6rKdZSoz9TIT
pvcqrJaETfThV+9I62D8Vqh+r4IUdYz+M9RT46QLAHztamRTmaX9BbCv0OcsGKnjX/tvLUh/7fAY
NXWVbJCNolneusP9a7xLhj47zpdKtikUmjwNiXhKpEsF/WmUUfgPi68MozZI5tFwBreQZUq3+n3X
xJsYptKawyvaNM8o1ibXIfTsRlUgCrO4iSCzxQPRPr16p7l15qYwXsHozpJseqfGYc6sz1cf5Pt3
uu8UA+muc8tPIVLnhWnsL2ZeTiUe6d3h70pQXWWx7k6luck7ecNiLAwnxli2zf7ODd1cfksmI+C4
k7LEcNsoeGDfkk5UYs8DkDRtrDoSxY8SwOS2SWLvX8NejKzrfb8TE6lRmJXl782bu+L9ROpa2vxJ
e7JJCkY3LjvlNXz53QNYnowk8LwnP1ZqHaLwPFuhb9Jb033IG9UUNeDC7nP/vXUPciDGy8PIXD8U
0ywlSehzgOrjwkPExaqbBnK3fuvetUM4O0R94NfG/yLgghMHxReWAGNCcGbDFK3Krx458eVBgQI5
hLpql9TrEXCZfut7YcT54P3hra8hqWVXVci+EwxyEp0u5WDqzziegVHaUDGM59uXIiso1OIEICSU
uiQ0QJ+84fVBpMCj/bTNYNo3XDpBRdSHjDQ8ypzuFWa1dHnpRyRMvvN2mKbFoz47mojHf+kaZsTK
S6+ipl3aNPPl9+JvGgm0V6bVp37bW1nhh3JnOndLnUEcBOWN4wIEgl5F8HG6nZaHnkKh1iJ7fn4h
1GgAZFXFRamhKUX+i5mdpLjHrim51vGUDaH0WACmd7429qi04n/Hm5sVL+jvuq7Yj4VxKPf//iFu
Jf+VKpvx1x9R2QG9nb7LfwY0MH020+83xa0RUHLn6MuiRmti7St/3wbexJeCTs1+mZMT2zeFI3FN
W8LXFPvuW+8B0bJmXYvynLgD5v6bFtm3WeQcGDyGdmn6W4ilosWmCfiPEiJ2Sb/Jx2KuH6K1hgbL
GRkv3BbJEaPS3Z5nK/arXSu2WBztBznCEQofNd6CM93aEVc58fejVpSs/w46qwUa6U5b0WOqmmTM
xWwDzRgNVYP3aV/ZVOND4lxDsl70WSQLc2AShMjiWFULKyxZAtcP9oMN+K730Hj9WWVyZEGxygB/
5l8JteVpelpaqHLTlbaRqQ3MwhqVCiH5wnLgwRkV6y00QiV4RcOaIL70t87vG/wcusuwXZzsCVw3
8Br/3dTxHPip/SxJHUw1XaotwcKHN10KhYSzE1D9CurdzDmAPa9QwdNjSt1DVt5GtKmeTEqUTU7r
yeb81qgjzjEQJhTlRAtr4UcGYQxBCmyN63x9BRzAJjK6hc/8absVA4eJIHHwHkEDYINgxMLWHxwi
/jGG3+oQtBg3bJjvtKNjVStbDzKPKxD0qxGna9rHnQlFqAFb4TMfnfWKQNFvZGPSXDWPofinCUri
nx8hduAjPwpuc3hH2rgga/YTzSfvmret2fyIxXusXYo/laRMYmRrqMVcsZ+87ZFyXTx5QUoF8ixK
Gw0Fm7BmDYttUaBQBZUVYw+QHIAZ0sVduDF53L5hW93fGdonWS+74Y0PaHiyObIiqC76+13xwXoq
VVUS80ht4TjNqGAVNTUNwDsUuIrOo0kRA9ZA9VO2zcAEGojT/z2uCnWrX5xEUP2+uvTeWns2efQW
kttOYq0+yXi5zfSA0OKSlQFKFohqYkcze1BgzGTA69fVW20OZkkkSFeG9HYODyd5JjkXOTIKhIyC
9vbWFuzJ2NBXTKlC1zqE04AIGPScW/926N8BxeuswglUZziMAl+GlF+y8ygwkBNl7ppK10JrPlB2
Xo0rs80Acel2gudqVqs6VTlKUzLb/RXVEWG4xkzL8hWI63Q1+XH6g/7gxLvdrZ+G+GnLYtq3sLpM
CO/8REd2YExHC7cF9hs1n3rZ3yYJQhBZ3R/oTXFYv1X87zH+NDrMWdtjdDkZrl+hLDvFgb5QlsLF
RROjZc2IUEqb/Ep11XLbYQEjiAdpnT9j9vjxPEwyJrDA4xw5PXjlnTSuTiySx4PkJYRSdkH/Uilo
NRl46byh7L+dOXu6QWhJy3AyAqhcIspkeabV/0aLRKZFKJDrCW8ENfUcrK386e7PjL8iwP+uB8cD
fxjVJbgLUp7rnLewPSwmfz+03Bq1eLCnsKmg+ID8Dj/lxPaH4sJrmFJSlZWUgLeW5LrYu0LV9lp5
s0AqooInzdElUa2Pjk0PEUv9U4RsULaNJ2nuihK2xda+d/nu8c2ufJPA/M/eFxNoZ7+WtkFeQOPq
qElJ410cI8CZ01m/8jwAJdzaudopKrcg8FhkgV+dj3oCCYTjCh0SBcEiBblFngBDFMRxeoPOtCMD
awMbDKajokWsGhL1tsrCXrPyyvAcK8xZj1HvLzl6wagrF2YDbHtZ76Sgblhbk4nQLwqKgYs8xQFP
kE6JpuRKS5NK4PZ3H7+jXkaFzLQ02moCt5ny1pw/htHwFn7pmANE9GPYyAs0bA43fdVSENqWch8E
4Rm/Y6rM0lqFA29h//3a7wN0ectSNWtOE2mFn4wn0gNihDIPRQHW5KLo5tgWrGFlcaBr5r/IEdV3
MctIb12qBIk+QyHUUDUlNMPCxtwNQlLP4N42Zs89z9Evk/tTRRTF7MOijq3+ZoFUGbKzliEKx00S
B5PfbkbDXpOBxKT/qCAnrevVtR1e8kpv8EohWtiUQF1t0Xk9CQa+gI6nvuQe/LQ5VP8ts8SCc7A6
2CI3C+GWYApZr3atwYrfdStlNMZt7QGfwbVodVMTncvYNQs3eBWmR/OZwsDa7FynQzWs+N3cINke
bxLtgyvdtsQ0WIjKAMzrJJD3dP92S7YQfxs1+HoG5BtHBArk/xrlb5t2EDoYy0kkOSRCLNJhiZe1
JG7QyCXwQwsaQXVoTVQh5us0Qo/02jTWF/t/5wp7WLykHQ20Gx7v6soP5MJx4BK+cTSvrYht0Eqt
WI1ew/QWPpHREYheT3GeeG8PjFH/Q1nOqfJfzT2tld+i7GFO4IeV9JAQppLcpB547E+Ki8b5A/z7
F3SgEmA2b4qw9xI5eYIyjI1ALE0PfmIamYEI7HthCjQSabyQY4QC3KNKrS+s3oPgswi/zXCCqkUi
skQN25vB0OAZ/2ZYp3ATVGXncUNMLD6aeqLSi2U3nhvB/oh6a+FOtrSpurvkzW9qM7lUa3ig/5Kn
gf5Nc7DwkOaQFYPrUYP6z9dzPPI6LSRWmj4khIQ82tLcHO9mDleqprY6I1wMW1Q3lcNPap+mJuo1
6qgrshyPP5JvlZHG89A5HCyo7gLceX8cPuvAcz2LtL0+uRgoL74MkCUs3DkP3d4G/HEi4XRDyyLa
8lpJJ9LjbRKmIC6RBi1GNrY7DiubjjE78/0qAwEZsYuOY16H9y+p+SjtmzgTqkkDsFJOfTT9TabW
thT1q/wPN71KW+qHP4E8bzydIPM9qlZgGi9iARKMtOib5hBHsNYwDl3G+DTVY1l5JzefD0V0Ayw+
tRZeX622rBN3vChbGZ2KVdZqXQj6cBobMjQ5dsPDylh9Bn5HVrmqIcxwci3vXJTsag5dRjJsI7gX
9Zn0wEiOktuoqeIsE+LsLv+/7fb2tGQaAORkmxqZyley3MHyk4epwmwobytsXXXBQGNedm6j2TBo
8mImgNEYvXyJZedKMDWjsDyfy0vv0bFWAy0dNHh1+FMD/1FGbVnAjmins/FbzoxRfG1sk6eQiWJj
kaV3KIPgPXY1znX+ZTkcqK4PnrOwUReiNzXZp3NNwqSKx/vIt+X8Wk4mXwGspFDiL3Mj54pVqHQ4
IRDco+wzJRRSIy+r/TXCsO+hAtBMyMCE7rbuOCJyjQZUngxLQLZbKpv+XEHh0BWFVWTcNJw1mCUo
bNlB8E5icKXPRw+pV0NSSKJIgnc01i0nxOKrCjNUqdIFX4YcUuUOeffxgq8iZCRu0piPW2K6c2MW
YCkcREr5D9xr7D1fvxAeaqmzWde0jRVf4/sia8QHSZ8RKvQ60pVYvst2hXYNNlGatskAhzDWjveR
rGYaIxKf+JQ7gNNeYhPliuigbnbDpnFuCVRKrAjq3EX1/JdrsXhxW1OM/lalgf72hGVHJ1ECP+/e
1oo7TML8A1cPBvZic04VCTZ2bE046bM21giBa36QpgKoJywekRp12A3b+vfIptSp/BH4YJ69RXOG
EuxfpdH7SRdtMiNIoaHJYATEzgjn6UQdRbQr/nLC1k3qJKHN1wb+Y9s9zE72EipJbpzVjJG8hRSS
v05fZ64HAyYAc1vjnbDUk2l5qfwumGhaJstvHsGMIWKP4CHiR/2LlhD92lZ9aAdifdhHD6u5lqkW
yPMK86GrZrTYXEQowP7j2ZRstK2S42JWpJcE/9yLmyqEIsQUlkpJXqQveMf0/BaFhzPsoQEoQt0e
S35AsJDggavU8L5kzvshjWWRZBzWgyXZZxMzD+W9q77vu/zA5EaoYpLTGZ9LzlwiFU9ls3Vzscqt
y7bH6XZhsJVvxWvURYcjpj0dsvwiHZ/3bcOY65tGIZ7EEI1Jvmtn0XICk/FObFWhECgI5gacMDYG
KXt8VXLc6ZAdFGXYbjD7rB8Pstv+1vqhRow4JH9uuHiFWdltnIBfM7SnQ7pwMKZpZktoeXXcmjsp
URhtIXz3nEOqdWgfYu5VNDoeiQnobJYV3CV5xQu6Ng5cu+u+WGlPuY6PPoBAfIj1P4VBFCf1xoFK
wjWeX8V+IxxM0O1hGL+hQkX9bH/PWqPJOB2IAwH/4Ih5Vt7fHLxNHBSZtLRz+y+pCVo9Gvrxz2mZ
JyWlaCOA5/w/7VPoRvsObGZAIyVBHt4KLOqyiBnAewGOq+Ru0QdERAJWTeLBBA3Y5/vANtnbE3KC
r1fcGFQ08hcZfsf2mq9+yq81RZ9lTLKZ7YiGtoyzspDA/ftD1GPSPLVDG9pdM7APzm0mSsgzAME1
o7NNKpDDtgP+nCHtQVnEuUSxIrhUjqScz5PdmY8x0Zt1wOa7f/p21/2/pWl++fGcqyU/PywPGXYi
/+FcO+c05V+ENDySDT+RFE6Z0o2n+N7BrraykPfsGZwXlSg5HL94H3jKx5oeaoirQPp7/fdauc7G
yBLD/uwSwWIRkC35ipUvb9yiY2AKkLlSzkSzZodNpxF4IxLLj78+qsDoLgUDePNmFcscMk+GxQ82
mlGh8fv5aod3G2F3a9dWj5x4kYaKTyIGckdA+vS9ABKlqTx1Sq4NGZeESjNJAQbSbCiXaxHmmoz2
RmMNdzeyUBpTQJqKsqFCS762kB0NZuKRiljYjXzspi/If7VB+4yMYka6iE3Fmf0jPjx2GLRLNDW8
9QGFIucwkuzypzG9y9l7zKzJitAOG69gjK7XYPDfy7VO1sIFSQZTqNT5bYayvjomPRvFmQRebm6k
9fj3NwafMSJfM92KpHksZdzmmq/3aVLDjkYqKc33XevtuImkNzRjzhpunrqHIRCh2st9IUkpHbJ0
dfad0Gsb3yQCP5sWCzs3fV8kArJntSPpCXcm4+qPkPH/dgf9HMnODHqB+Ns6FbWYg0UD1egnimTu
i9iCWR87wq/4p8a20zycgrw3iSr+sMt6PYJntLb8Tma/zhZcstYvfAuSqCBxxCw5yl2WjVKVZFrY
diQTzIM/HRapiGzdjSAO+wx6wPMACocN+48qSByH9lfzVe7QjnKxAvZR1zBFCidhTRnBl1sbxcAf
Fwb4Yo+2hanMZY2uMqmS6/TWdOqdNqLI9LnwBKgfWtgHU7hRmfzLk4MKnlxDVOe3dY2jryNGbJtT
cP1UY7OkSJrh1zc6/3VZsP7xFla+RqFnvk7d9u4Fm1JyxZwNcaFIcWbdbZv21cnEbEmEvWrsWcxc
TlyKyvLp9nE+GtYGpmtUmJ4IrIxdDGcPMtPD9lo/IZzN7nrLY0hz6gSKuFZxqKAgxqCmkk0/bT9y
4+O7rN2mbTce8Kc0QzNUVVzI3g/aFCApdmi3ihwCOK9ResTtEJ1371v51k9jBo9TsFp3HwmEHPwC
KkI4k6NjtouMUbOnKmgwpPT9dvyiv3A+NeyMTBN/9nGsS8AkB99PkQdJRouvfXF2ClZRWHlZ4uMn
T8UcnzHa+/h1SyLqqSZc6b/umzUOVK9j2gsF1794TRVi3KWQ3S3e00sfSXWwGoa2VlE5YhVbF7/L
wRjIs1AWUIzgS1W8kWx3Yk9/kEl3ASnjafkgQXbEpZF1uEv8Iv92V6uJJBqHQ9nnA1MQWprLLHqi
hak/6Nhr6swGGAzVB1OXvLrZrZK2R+/ENzvCQHLB8ra16uDq7Qh99zCMddq7kzzpn59kEGJi9yiF
6DvzKEUmDoINQrdR71k6BoRFDGE4foE5espwu56pnEMjMJOOSQHyfmomuOCzzkAvWYH6j8zoz8BC
D11s4swkB6I2sL7/bCZBwsO5dMIpbmr2gT08hm3zZEh8T+YohzSoniIm4CZrnCq31MwYeoVeLg5t
yQi5nM0cQ5iH8+9izpHlxyMpRvGoCimK3dc2cjOuZcJW/NWGHeADJcEzhZhVLV8EnwguR81PpHhu
XNijawdFsFKtC1Aw3sRrXqQE01tz22SeJU1MYi6D8DsIEIObc4e/fpaR7zklphILxmyyfifeahn5
ABvnFRfHsPtZCt/2Yk4cj3zFzaR9ooZH+VP+PzNPamkvPrs8+ZBz0QSbyXw78N8PYJV9x75aHnB/
vkYbvsHvfFfXRMP5hQ4DXHaeX9T3vX63tk8TsW8UapEZdbi1JYeSVYqjX06DChRxw9dnN3t+Vkbe
a4CwE+yTh1Dch3DMnVgHfebAs2l6iRQLMp76BGnWFFSeZ838AGsFVxIBtXiS3GrhqTJ3zf5gb2J+
FV9xWJFle/S4diBeGzgVzZY7J2wG5jkX5O0rmoChxBclBWPmXcotEnFziAKaqCzO+YCvQWAOQ9d0
6QSCgrSAeL07hwpi4XeLcNkuUS8eJzA6U3J/QYIqONQ756bxroUOkyj4IZ6fxeQavgg/MdJTsTIK
86CjtaDWgGJbBhrchDT8iUrU4/FOk3GZpBQf8EB7haqFVxQ2Gu1GIXYHOkOHH9cz3yOWqVpUDkvY
P4mRx5XGoEFgyrGdPqh2PGVFwdGkp2GfAQXojfR1bkKZEEvRA6duzE51/XgSUFkMtc9f0wdW6JI+
E8b92ta+irA1Kj5MoaPtDQJseOk+FBIMYfYj4binSlYSwF8fiaWza1hHpJgmEXvb9x/Qt//V/gyD
5SAycZV95NvqdYD1vamG0THYrIH+SNy3uJI/7m3MRexjJj6qvlkjJXNBchZzFfqkT77FFnmiSKYZ
SQuxqFugY0Xllshp6QqhLut4fZZcex9vmKx8hmp35VGJKRs54ZiIetH0Tb5dn0uHj1A1RWQpw42L
c/Lke6YvEXmhBNiJgk70Sfwz6aFCc374PcXKVvEWhEB9v0q25X1BAEavklzeaTuuqXlc+ueuukLu
C2DTmlUuHJ62FD4U4FJ9OQTv9inzGerhQ0YeXWiyCq7245PqukJXx4bq1oeWg/3xc+Dx0jbvtfpj
JS05PTKtXPvRcj7hvsTCFx5tBK/ndFbKRzmKP435RwObLKX0ENuIyA6832Cd14FPrSWyPK3qyXhl
aU8eFcH3dVTUA5cLQ3ki0cMEHnYC3wF8S+FDCUyvactVoqxzpnMvUMQOesTcBosM0zzL3lq5PnXl
8k1YhwBZQqk/XoCzTA/wriVpwJ6tWrcnIfRodRMOawzirOOB97N3TFwvAZDKtCPqrxRyj3NJFg3t
lNWIeXvcZ0rP4N2OaRK9hxRtWfjEKjnGqtfb59TdDH8jfhcxByfrf6EVzdv95emDN76FWIefumaB
GW/RFTdxAxeM4j71Al+sbCF6GiqqqANfUShTLEsB7tVUb+orpP8sBVwIaewQqCmVZM2X8at7FOSq
xETB5DBvZZQ9pCNCqTtjXS1g9H7zA+sQZRCE3UVHhyt83DLLkasJdXDDCe4KZPdkEwJZK/3FZDB6
GhGPlEUSYw6rHmVwyQh4MY/Bm0EyPMpS1abakeUnVLa6UI7+9+739m36XIfwscBeTROPz/efyct5
mpY2UIroRzKcQLMo8suNeMB3o2VCO974rm3BCB/ehfRaiyRpOJWJkkC8Ht80V6U36jRIMplLJALP
tzd1FIdzR53ZjbbYnhZEt0IkaLf0xY8hcarpUpOdBw+EVadscGoOzHx39RWPC1wOEvYiJbOzx0WR
voHMZQZS1iTwc1vhd362jn7sBAxNVlyov0WXi3Ao2LwxLq+OhsPTYtD5Z4iqBHMmKVlczpEGStaE
z/HZfph0NhhK93OgF/T5msdM+pAkCDngMYrkkFDsWy70iKzyyScZ+6sYT6l5Cd1Rbcz8CKdQoJod
RT0HKp78KEGCXhRVawsXiKE49ioPR4eRukYnSBQ5At23QRIOGzo9ntywqKU4witXqgBRpnxqvONU
SoJkgGm/UwFGReZJswLW8hD7I3aD+kFLk8KV8eypz4HvtiewmWqEfOoBItro79HetOwcxhmVCoTV
mNtX6+YDulstyu2lv6dlP6ZQ77Qsk61yxHuP5D9ZeowbnEb3EjZjQAjW2j+yb1DNjYo3Duj3yw8Q
fR/o53uH+lVMPh/QMrlY9wGVINrK77aF+SMEFYg8EBHm+uAZ7kpwm9J8QdJ9NYXAk4hdtYf0eIcd
5BaSvfXS034X+//nZQWc23BaEDa1MkKboPmvzzVBCW2ZXGiZsSpzrSC8SNiP0RyvQXh0YU7YW3c/
zmXpKM0KSx8sXF1SONykG5l7tmb3XiE9hxp1ia4tSsrf14f7KdSBI9IspvtQDt46sxWN1ZMXsINZ
mJRg0PZRxtsGopgAdWYSi5PX6hSnoiskpHyj2qBE2VX3e/cwhKChGnDl49pnqOFgA6f1bh2a0dZJ
Fv3Q0NnJ+ImUyWzyB0jZK3VeP05Mc7hO5b7GYM2T1tEbwLBLbwgGB7daQS/GD/B8QPSAR1XXXTCw
DnnOPUG8FOle8cNopcZF3u4XlAbs1qnK8tb63yrF1eDkyeax9UUciHktFR7fSPCNHpl4kEpoviYq
v1vLK9V/mHT3yFaxAfG7GmI45bKY8ncH8QtQtKcn96ml7qXj57vFD5KwO4Rl9AnU7XxiAKyz5zem
JM1svOAGW8Zlb9JuTD/lKQeTs3T/iqSPHyeqXbxXtzirzIKW1qRhez4n+GtjAA4+oTkSmnvHrfGt
KHr3/ye04pf1qTDSIl9SQvNp2s2eYktD1L1XEZL4qEqP0rJtFXDwVlU7DBjSrLgjvJ5xcWS6p9pn
cZBJnOjoRbtw9z4pXvLCMcU3jvHjZDCI+QXh0YvJ8ufHzfmbYeosXAspRCo8tux8AQfAkFKyAr/z
xwtgJpmMYoPPKLY/hRzp+KhfAPo8e4W06WHf3lQFeMnZYGKa96kIqnTGc6s0CWLpPHlPn+/dk5WR
eDNvlycbXTH/ZvYVT+NvIZQsRW14NWpWc72PJ7Xf0/fvemM/B2y1KUv6QYmnK4Ux7p0ytCvQclwl
Mu/olc5re7dgKCWo9PKRBHFsMt6zofZ3UMpa5nHMk1QTRDXiiObgRYBB5NXf/bxG3VDRP4mZbK4y
F6x1bAO5ooBjhKdYA1phBasN31KTxkgjH0qzD7PgWBk4eybcGvreyTY37flNo2mMVuguuE+G+J7z
gcMJDXiYCTA5vDAAQN+CFtQxr6NgpbPFPkR/EiF5f+2yMABNW+mg4T61BnV0wvjSEwJV3OWWOSEL
HU3heOLFBIrfzn5kmthy1GCLuvOXz9dIsO66KHMatgTWtysXN0pcrE3+m3yBWVRCzdix05zU5HpX
xDTdLCQEerqHIw6OM4cFOixU3+VyqS3hpHjFG1X2l/C0bIlShLkMyK90NZGlMZ4A9YsdWYUi7mj5
nI6pmPGfKXOOvnlvi9ke94OwZXR3y7uoT5hF/yUybeXMO6zTpnphOa2XhTjSwbGyJZZq+KDaxVlR
MJWLv8Kw8Gj8anSZJsBkOp8E/yt097iOinbzChrYWkgcx40TRyF417McfX3Di45rmvYUmYEHBvl2
VNiKTKbrr2k62ycyGLBEpoofBXDTLTnBeo2yfXIWjSDZRkj9oCQ8o7eYqqXv/EaKeG390n9raw1d
RuJxmzHooygZwMnCnscjS0tOYt1hKZRiBNyD2gNFG9NyN5gVOhprBg4+Iy95Uo/qz4qW+JPhVyiR
MSwYOqsjn5XJ6UuPHKqdBlPhuCXMeG73yHOS3oc2q0MkLvdL5MA662ht9GaCzJOkhc93Mpoq6B1y
ZmqevvwUrb+eIwOkVhVhoDcVueLLisXajzR1szIDVPRp08EW0DisOQI6fmSudTIKuilOaKdtm1LZ
NFY6B9mx0mo1Xr40U5mmV/uEksN+2fX8Nan6XI7l1ayNInEIwiWYpN20ApboJLXPb5AT5Vij2PKJ
rDvUPKrPtrQQBYGKNxbRYw1mX8T69tHAKtuoExCAZcgKen1Tv1sWGHFrVfaVsySk/PrVFaXO7JB5
aNY+Du/LXtas91qOsVY+IE0GsChMEKbd9nkuoxyPL5jFgW6rDdNiuEvaKz8ju3z7xxrm6g15UZRc
oUYEIahJTZq4mTIM+P70n6+VskieNX0UexlyIxC/BzRmDPli3/IFs12VU8hix9FoZtoYJ12b5gWg
pY/E5QELKMTJz4IJDct9xU+5VSIU+VZXAy5db7xgTfI4oqh8V64nOqLVu6d2meDE/TAykMA6IcrA
gKcKkz2ia6u6HVfXnXxS8bfETyK6rSmk1jZ6v5psWH2Cvc5CGuKoweVAQY/GSZP19mF5/GHBBPyM
RLXft/BDBoGVDFBVbM0sD4p1CNA23LcZU7eO7I/GfZs8jb5rplneI+vtD6n/26Lny06zf3JIRYYI
5kq/zLuDilG4x3aXlyZblqJ6F0LAiRx1e/WtLaNp+GRRcOHfULzenUhSbv+wr7xpWNfeEDUGQIvB
pjxalcWZ2wyyTuw9C5IEyAAtnkmoUb1gkQeoF5iBj3SslJGL5MgrapVwVJ573nuD04LoRSePdz+Z
1bySsJJ544FJ6TxiMdzGFaun4xtHgbq9HMarmwB54XheuEEN+YEymQIlPiCt3m77T4yWIOoMShYc
Yb18swH3nKDzA5anDXkjhmCtGpIthE98dWxGpNHI98PxfpEFzP/JkTfx/G/POSeLANeFTUs9YyLe
4mxvBygjgbuEWfFfGEL1hPAyF2HIsb6mbvbHagAeQTwHfR6+Mkc1kn9aIByG467I2PcA7IF6NN/n
GmOZOvjK0Cbw9+N0rPsP/+T7nkElNS/DqaxSytkkgfrh9GunL7o2XYXIsyxPpuMlc1aBUqZ92QLI
HXnBagMKhOc4FGxhHsE1V2/brXLiRUzzUwlQPiapAjI0xWh0NC3VxHNgiLRlhVN6lbuSpuBOvGGd
/PU268cqTCxHsdEhzTkRfYxj3VxPzG/cN+aQD18iP9lwuYqOp4yR3ux3vQh4YamH+RmBaQpkbO0m
0kVyoSX84HjHxlLVl9Xzm+Brz9XBJcPTCSSdIZRdFbmESF8d+blqTzMBcSIL9lRUaAyEn1QH/UWl
7/ceRUgACC61wMdlFPepRN91Uhd6Z9ZfZUuzekAS9AL8BLR0cJ9zSOYPzOAfkS4RbbSmncZY7ksJ
OKyjwixQpALY9RnfoSH0HLnWagQ02mRJiYOZNyErroG1x4uGQxuFcTVDFLyM44+EjG8MHErXKHgC
4mtNqt8H/o/RaYaAUXhjcELYUefaSDd9R3eAClQqaU7s0yjBaSAslWc3EZet2gAR+2R9rIXbCnjr
2/aU5Rdv2PjMmOo+vtVikP5qQfeNY1l14WwqOWk1r5oC8QeG/giti1zI87dQ7VECPiOFwm8TTprk
MOGTRyJBrafTE8amxfWclXGVRZ+dVhO6C6yXctwWzwbrqmR0kg3LgKR82k20nvXlVOiltVljG1gS
TYJ/t4uyq14fNT2R41NNlUyBx9mf/nQ5e6n+FZ4MklEghene1Zo34gu3v45xYQWJE6nHpDwGAt5G
7+1Nm0lDY10d8xxWffWGIHux8NnWVTYf9fHf5hvZBg19qndi+sJlMNyaAawmAYMtLSSkZRyz9dS8
FB+giSWbor6xnywf2uqHwgrq6m3eTLpzy+CsGoVZqBS+IyV5HeKxFC5lIYODBZWroy6MTOn4YEpn
jHR/Gt+JYc+T0F3MdGac/tlOekgX894eCMmKCuhxv5XMxC3mZYoCgkBzQB8sfiDe2B/IIDzNU9Bm
4/tAbqdBQySHEYx+UWSs6SjFLDPe/jsUmQ7Z1AKVNjqvGP0touovslP433MVymFi23BK0IrQ+diC
hSRHuSRzqjW3fomA9+EBKnZ/2Nf46lRzGF9Xo/4VD8sKxbth5+YnYBUXxzzRvm6z4BrmOWofHN5O
HQMqT6R/aKZGhkvKi2g4R+CLScVe0E+Whri76afppDkJD7y+0lEYyTHQJ/5zcqdruj+OAnYkLJB1
rN7k6dHKbgNAAbQjw/TEryy1opQ7XBpS8QK9za+QAH1zQ5q4izt1uCSVoOrIBzCxbzAizK20bayF
CL+bXly9N6yzGq+x3N5Yygw5MM/zg37J36OU56a2jBD6lDquwLGqkOaUqWZw/KLDMEkba1+ELESp
bDtKm5a/ZcT3HOQDZQB062rBNXH1lVAW6wErbALs1E9DO7OMmrcq8ajKmTUlo6u8+6BSt/yMKguC
Dz80SiZWm7N46Ar6amOPzq4zuryLS+gOdcB3nXPs4V4lM5j2MKDhAzne0G3GxNADcPu+ZqegGrct
01x3knBvrba04kcj2DC6rYCdARTiHry+XNGttXn5ahoERrBZieZjtn6a3FL97bcZ5NZ+LTebjiOy
cgNTLtbkmkiEr8QV4QXRduOwcJbdgOrtwE7iQJumbxEIpD2PO+LljoywiQa0OcfS17V5/MAEW1oI
oFdMCw3g3pDzvU96dTEPnhSP0zZIx1JksA0QZQtNSx6uelKgv1TCNelYvpTVezeNEZaOcU26sTox
ompcAysqeQEYifPToiCcjP94EumIC+E89xJZCcltSVGk80xVrcHdv3wbsKiofHOsG/0yNSy+/Dkd
hQcNNWw9xTeniAgd88ZOiAb81xSKDfGvENqHo/xRhUQ6KtPxKw/jNXrmiS06MMfWS902fk8KWUgu
8aaDAOzjkDFRudE/Y1fpiQRnIGURN+2V82uoLl3HJshQVnyuOqtp6kp2H4m/saHBoex25WvEWDqU
8mXbqpbNib7ggn3YJasbNam2pW7m8zwoZh0CEQefSiBG5/8Ya3ThijOrKswuBuCtLRjT8HVwUXiW
3LEUb3zeEZ7KP6HTnQPgANYQN1utSBVpuXvMBoxuRvs8PKIUQOVSgcUjTkIQmBVTjS5kqeOW1ep6
JBVRVRCOoBL956OPSXoWbWU9uTeJwBfdWvvsJLv8FXJCtWhlqlx4lWiWWGLk+Do0kG/Kyqa5Cx/6
gkZBeZlIVF78pQAdmobDbbB/iyF356VfT1sLQZ5Te8ag2X96N2Ql0DV6gl8BdWwfWvDZiVWPjjT/
pOgTGcxpPVxnlLvioOR9EQjoucynRfBlJClW/4bBo/TID4Z0KfvTs7b8wYy0ajrq+a+cvNCqxsJR
q1bi2hjUpfYf3NABgbHkZQSkFGw+WWAjcSA0gqScYb4fHxPPvKGDxYeEV4WKd2GwwQPDJO5F+NbN
XZJjb1axvHMcSab7Rqu57lqx6SDXXf5H0vGGLP2zyLEcb9FBnh6t8TenceMcW+AaKzi5FxY0uE3f
mc7NbHIOOj6R3xdc6Co+nAwMOPZV6zBcgB4xlD7C9qPuBJhS3/O20mqg6PBHtdG9UnVQqbr7sYOg
qT5+Xa0g3YE9Tc9cIEB/RqETAcW3/FpLtmjWT0i/+lNfEmcCzaaGm018VkUV26IR9MnyDUHndK7c
g7MH/DZC60e1I19iLrHXDmVJCpi5aJ9HnkAfbmmSTR9Zii83YC465d7qYvxN6j6l+ey4+Ze3a9dL
UtLcNa0j4VbRbCrGVrx1wmoVzCjBMOJ6Mi0h1hgi5jQjG6KEsyO/1yTr77gQNazHej0DWnOwDYIl
D/oPCOLplF6vnCa3XNXUHPICjU/ZT6t8UlbhjajESfO76c8k85N9o1ODJWlt+YoZtp/oOQNh2LHP
KIbKfrSeQwFl2j+bbbtDJrapGeinH+UGSBQSE6gutjp9/mVG3tyN4+MrEbUtw42VDb30wb+cywIT
rkq1spohVZyyZrB2kNKYdG2Qau5DVhhiI1eo2EL/LNbmOOdOJK1PI8gvKOOubwkBV/D/hcC7e9nX
9ptEp7WbuTpGclk4PQ9TMCg2yr6nQ9IMpSeC9yR+vtOHAF85GHCY2nDWkkxO6utKmqZ2oZg+gB8C
G3BGr8bdMSuZrqaFtHA2ewPVikonGKBM7zugQxQIQCeUiWShMeBI1z1yuWiGeC3gpvehPn8hDrGR
NMCXMqjf5LhPAqVyMxP3LmFtq1m35f5Kgu+V1AFrbi0WrM/P5PoYBBQr3c8OxoSXw0tu8iNY/qYl
75J+BtJpCx4LTagljps/ZJGguvbGJo6ivrio38INom8yDMPvK4q3QX+ISEfW7j030mHg/dSLwris
n5/MYMcrJZdK22KYlc1K7NXnx/iIMjMHUChBZ8pqc6QJio8FY3scs/H9RO1SiYdL0Q/gJzlXSaA0
2Y+n62e84hl9O9Qqj+UmwJ7KoB+qh7jMdmgLw431KY1GZLKlxMedSrjvOlp2SiJtzWYj40UFk3EP
LCfUhKWiMxj+97MOuXi5Zg4UKH0mnb7gocPDHXKV2e281XKjJtThRaMIHj7i15pygUoKGm3lWK/U
rCsyOkzt1RI9JLtZ4UXWdgpK1t/mNTSVlU+jGl/sGgigMrr0IPjLWYTZo1EgXZhFJfYnKiITdNi2
QAySF1F7uSKgXKi+N4/BlajJZgjxLbz8zsrOl/hJjqQ4sVFIzRcVeZpwQ1AXxufmptUTTRyv2DCd
6agc3BfObOIU+9xo5HiF25bnL3KgJuT+Rj1kIhrGqDLKdgFqGyx9TUaZXxZVDr1GdRh3Ex8YMQWT
fUaQGPQHE44s1JAvqdXAkorX54fXuzdlfIgXmHqGvmKwY+OMsc2WBcBrCPuFqmK3xuErrYQiXZOx
l3sMZXp3iEHFEJQ1a1f/UIUZe1L5+6ZRP9PkMXJiZUSqlrH+HWTluS+MJCvoaSZ8CVABz8KgyMzg
Ac+yvtad+fXXUGRuC8yAldQxySnjvEaBz7fgdRqPHh9LAW7W0u9SLPHebpxpOUl4D0raBWv6fw9u
AsigwhvUpuMXWWrOzde4hCChqv60e1nHJL/N8xxxpUUqbtyI2t+30qqeodAPMt6wB9qLKuo8Y/TU
F122d3svOKp/xeQJuwUmZDv+fogOcFLhwZsM2VYlcS/1fGAS5RVTSsiypTgo5M2/jxhurkXbwKX9
KOgKDrTRfdaZDxZL8BvBp4QTyNc7PnMXQ4FP3MSAWxsUc7oCpibIQ+MJ+xElJGd+rK7gEx3jut/E
IIu+0I0trOl/3YsaHMYkSVXA1ZfUIQoPbaJVp62TPx8ySF37+sOhQTkUuXb0SuClwD9gcgrS7st8
gsOmEkscpbCw8lo7rPnxB5YR4MDhlCXVP1ZzIJP5RhS8YU7OZHNsxCaceOfpNX/cytjJKHl7t1Ge
hCvONegRVF2eE95HrDkeNwiN8zDoQZHGUAZkBm7HX2gTYtl0GPH73RVpsoiCYikFLzlgefpyFzUk
mI8FLXSj0R0DzeGCGsYIJMPR6pnhEv2Cc3b9OzIYWCK04coeTJgFRwQpDW+u15HoyM+FnCCfcCdv
R5dAdvQlvkWZgEe/Cs2Aco1Xn5JmN17Inf2V66eJ9/1oGFxgfNBzSLesldK3F0fTCJR2Sd3PKd+n
vhHPcl1jpYXirVAqPphqe0mRsXFrge2ZuqRF12GvZP+ZiafP3ETWMfkrc1vTRsmCSfycJxs3lssi
b5/bYu8ZIjF7W9GGh4FBgQGGfjL5P2i6nE0rtiOlKmHHO7cJdr71SkkO1y/0kwC2/lxTFdWUWKkN
0O5Via/AaLtr5YWjBueWcbRhW4hK+I6Tm2+I/+7XsUBj30ThWTCxq+GJ6ULVynpYPx2xV+UYeuqH
hr/KIxOpWGrTYe0Mkf/VCckgEiPpGx0iU7kWDUj6HsWmmKFQTzei5T31rLexcT2vIX3A2GkENtIv
woEZI0YEEEYTO17QMKHHe5U6CRsdW463ry73S+Xz2arDvAJEZdi68NicKHP9ystFMiAEmw+Q/MYj
h76Dks8stmVED9oEV6W52iJC66CylH4klpCPOoOXdFsHc8KUKaW4r62HoMvb+kmNcP7Q3yZY7ic3
APKbaOfKc/X2u8dN5nimPORCWEqGRnNjtqQBJ1o5mGsA3zVVh2PZOaDUzsQMbv2kwlx0EmjWb7uv
+qxaPchefF6yel9id1Kn+E92I2uCAlWRAqTmbSGydP30Emn6Nj8YP7nbsJoICq4nvLnC6DBpRHXm
Imz0vmwGmpg+AQW//yYUpycZyJVUyUipRohwp3IPrDZJpuh8JSWqarQgqqDU//iNy4afCdrZ+YlT
9MKNKcx0YR5MO0Ku1nWt2dWrA9rvID5muA7bjVjJRYelc/pBnNyOT9JJpCcDKLwWTYu/yv8k9UX+
CvIxtVOPSeHS3Eshm8p71Bg0FEun/WGQvG5eJWhatdWXoLxMazvzhjqvSgqSo+eOlEXzqmd9r68a
Fmms6axV2bNxtmPUKsZWXAs3UXqjC3bkfIKffqaDBrOOn3XQVoeIKwZtJgIDyW3WlF4OObKu9tny
LUD+mW0YINvf4AMguPrmjzvQbsO9RaDd2fKppOS1Q1Bp5H36C9ibTMtjcIzK5P45HZCqAPmCLsV+
TdoX28ysuR3hntc1q72m0hberz32umKXs/A+bDlnji2KPTAVw7RJJgzmwWgOMDkZjwdxD9z0pVK0
oSaUBt8eqY1lV4n52QjgB9XvjqDEfRo1yf5kmdXxjNLaaEvlgzgmVY2n5BAF97KxLWR9AVK4HJSk
Ib4CLoepSkobqu+1GMhMBQPl5kLrtwvWpG6mHUNlFGscFnH8FQ19Zf8493kIXob1X+4VeHK6QFvs
BPJcx3iii+3Zfn7dxV2XPNpR3CCDtWCXHcE+S9HINogQau+fMy4g/OicN5SZ9+i4LKln0j1G4GOE
as1hIInNXH/R8yXV8PLWp4yzzWfC1KvZ8CE7wacqvE79/m8ZBnQa9lcY6djkF7bZmBZE4X9d1vPf
Y9Z3q5qszbtdsZDYTBGDdveF9WbbXVeQI+yPLG3sYSQMCIpOAvZb/Ryz3Fq4cDPJI7cOS11FZZmy
6xh2L7FqXSuwFg+gogE9VcqTa0wiGhAn5QJo73+N6j4zgRaytgR6cq7glt53k8jy0BOvohXiAoc1
tRq5Uuq2X1WY3G8cdYXcVDjWUX2RC2Syf5+8rbwgWkCiaQZUhIBi3atmGjZ6wTniFEjj5e0rOIYS
/ydVyLpHHZWLsgrazVOm9EDN+f3ObOufpIcoF5cZnsQgI9wfxMrabhL9s9WWpSXXxL6cfrju4Psl
qFfWcSzHBzL6p6JRb1H6CNvH+y7fd34W711Cpm5HIrEr5XG0t8MMaGTh4yHhnSv0nPQKqXv3qhmK
lxx3lT3xw15aTA4fjrs0lRJOiigSC0NJ/5dcEclE2gXfLUM+9nNFdQnMDpr1GdcoAEIyJvbrH7DY
jM8ehKXDef0y5RYoDP06uBZtkw6PG30CUwzY7kg5qvCw2It6RfiwU9GXdVMEr+6EuftFo16Y3gE/
J2wGKY3ETPc8yAndlibH1S+dtaSyKnq1wYe1FM2PI2I4ky+efZ6VrV71Dl3SAjSa+UzKpzOQ4wle
B9eipFhRCEhFiOxYNINJL+F2jY6YW/XsvEInqkQdvfnRx2ZpA3EuRi0bJJropVxm85ESGeE2yV2K
RiL/hWQFntU5ZV9dVkK7D1cdY7KK7w1nHMc8qTK0tlJh3errzv5z67qFeZscdmSwmrNavYqXHiAA
iRxo1+4E7UhZG5HpjAtfGoSrvELoZWG6SXfj+fc76c4G1IFGTa5TpzzflF/45+wBKKbEbMd0RTkT
6WA2geCPKHpp/0S20ayc+3JbDXEcUfuBq2nr+9mDsclx8Zw+AqOl8QI4ZpuuGzCwtmYGsBQe/DBQ
OOuyaoPu+FpN6ugwAU33WkcmjhQMJsF6SzfKofPmlgpG1PRDYD3POIMuHfviN2ZbYYTGH5VBu/KI
d27IdSErKa4JRNdBAsdF9Ec9GhaKDncQ+e9GFl6VSfPq+qAgN1pfZkzlDfmLWuBf/zTAgIH4egAC
sq4OY1Shof/cGJZQ6EkAPZe+YFzumCkNMco4j2IgMj4wZ016mJpyaIuMiBPXlmwRfP79xC46sed0
XSQGrMQumMNnZUKjGdTBws9GvrHRegIUJrwVYf77LDuZrle5T7eNmDhTFLJQE6dL+LKjjxyHn4hZ
/8TU8sEk+gcmcAYToGKjJCpKPoGG0gUTdlgcCek9CwGRgqGMhVM3zD1q87IhhB5rLxKB6N/IyigP
Wjas5rHz3Ne1Cg4xsIeaRxPA0o1YQ/DhelJNU1p3Ypw06m8N/x8ITbYKbZYBp06RQk97Bd/nWXoB
7wnoL9FJRLZ9aY9Kec1UbSW25tlQHU3NHLiGAwj+g43AHLMoDdsxtbspkVh9tbqNYa987EsDAe3T
BUQOOzmkcvsINTTfXzhJ4AKocDn2CkycBE2koLqyu3MpqqNP9dMvDtsCkMWdibRVCoLDppmM5qQ2
wnAkBEHkuDfiK6upYmPLWqh550NXlEUsr+ZMJlaLThmUf97K+51XrVCLENQN9CMnP7be0Zdxj6y6
1ugnhR4sFaCDLLrhv/u1sHzEkySi5voLvOf+v4aZbapF4qPNoKbgiEuutYfWC6Die5uZkL9nZjBc
CQSnCg40oFqbAkdZ1ZJwK5+ZuLpy/eZpnPwCEzMoxOACEAqABCql7d8sXakOPXyxqZKyKvsqnYZS
KfD/Mc3ZAi5elUfWO5L3OfcoT6d+1ZWJosEnQOe4j8j0oVV+V/vICrBagbr8K8n07ReXkERxBc2N
aELQrL/Yr3UaEp4L0ecSMyQnbAr5PF7NWvONCweuhUVX86Bs1dk18Jg6jmI+q5eXCKR/qcPzerVD
EfZnr1OTo3BTgR+7UYFAO+hzwMshsTAX3YoUndkMDCCQ/ylsZIhHoLkPdei49dUHJDgebtVkne8H
K4ldnZeic6S3EbQOT8lvNh3pTPS9ZHYr9hFQsfvCNeexYk+IZNHRkMGx4ydppJbM6QqZ/6JNAqNc
zKEPEML6jOerslp577DI0mGBvLEOFW5cqT/jMJZRpx375NdRjHfs6ZLdEmdzernJiRfrKu78hU3D
iHySF3beigy4sYHnRFkrwULYfZ0SZCrv7RyeRHDF0I6wmjtUV4RoTAQC2TkB0/Sa5A6k6mIVY73e
0W7ewAlsCi6rgTYdjMTuAUibl87QKvxGQQ3daGxp6Dax4iH9qBGdgtFrRIM5vzQVlp0uSltFOcXP
BqwGchbaYMMeFEeCSBP0t9EHFdSccckYsZfjuq7QtqiEOFCvfnRAfiPIGQf2yTWppYa3XNSFwqSN
KF/SI9r1qgbK/VviNa6zylVjvjnUtztdM9QWbkjglnD4PkKceXLfjzEekQQ/Xm1Mc0Gj6wlpzHRs
VTgxChH/aaO+mQJ7u3bGBQynbDy/hFnf3DMhJ2e6fw3rlaszIOioXoNMG8P1r5/FQ1Bhx8yNt7dF
ZyiPk0MnQBkvW/1QlZaIcIgXzsGm0vvIoRcbMPiJitsdXiLOG80LdvYU7Otc1Nj5Lg5FqoTcKTAO
YS148NvOUnBZd16TDzYx3Zt8RQQUfzQeo4eAWfPbyYbDi254/Z3qiKH+EhaWYpfQHz2dSyVx4/P0
IEcSfwnfHiFyPiERi1ZfCKV1RKjPGMK35Y8dFFNYyoreyMsvsbd8zceqdZsfNtV/ZkLkQ9xaVCYA
WOUBrBI5kUG7vZdd9zhjgyGE81xx8tymQY8Tw3VsLpij49GxLo4OLww/IIEE62RVKwKhsMFOSDLI
jcdrxrA7Thka/NIqQiFAR8sEh+YlUt8pX4R80QMrkMkWXFpVq7K15haPt2RKwZqFAgCqRV4Al2Xm
YqOTItdTfAx/f3+BCJM8P8OAQKO0TnF1TXZqxlbGjSSzTGNJDETU9bbrkdBGetkK00+Mkzu+nVSa
7tj0tsBvW1g51cxlK6cSt2Sx0h2Dr9+iYxUihowwKNaE64FMnFb1F2PJ/MhmomL/adEQ0AVBuuXj
dvSrhtS5xU2p9/hOyPcFfyTue7aQYGrKslg5bmIdPl7+fcEX4ZTBUQ2pcPFNKQ/PMWVi6EjBsy5C
9uHghFRTR4IrvVn2/yl3OgW0yuoBUCTG53+2TAwRpByImluBwOaHc4LavxOjPYHavaShdIPuZDUz
Yq9EcY28GwgKJYJ9WRDLjgu4Gck4WbX+yaUCA1eZLvZNG39tnBMd5BTl/eB7ESCiRxevTmDZy4cc
gTPxGcgmdU2D22v3JFxYWzOOg9dfU4dLpE68MXDas7s4glXTL7LaTLhB01GKJkDGNXyffF1InQr4
5CxesxFovuhRPwmeNZceQrcrl67Fd04UL+k1zP/REkbCme3eALxAbKx9tjzZpRoFPJNtTGJpdm9Z
4IOpPPJJMMixDxTt6BUy70Vz9NKFQQqkhEouuQK3r0sMr97FoyDj1A5VaPDcKf0NGhV53FzKE5lz
SY2NChkA1Sz+xw5NPvOe7ZzwNdaUOT3nmceHLADsyU6LqA5gOQ9DDY+j7GVHxt2333Hph6/AnsYl
daHZIRdnd8cQMQAmsqpWIiWnDCUqm2YRASOeRfbTmdP5BWNnY1otPOPQBmrZIN4pIvTCAu12bXOo
UMDE3u9quvMCI/b3xObhgop1Ax2qfOxXSD75EluWa6hfAB/YNnB7P9sqKhgu77P+j5uCOwZTfh4A
i2kRgj/NDf0QDKOWIaXUdWntbIKDawUtuBHVwsAd6d1GKYB2s9Dd4kjHvTNtipw2Rk92uz4L4u68
V8Maaf/8jFnWmlJbDuOdtLtRiCL3cMZvyyizTUdnSt3AKZz2jzQSHe6o8OwpG8aZZGw7dXtNEN//
C7GfkNpqVOvwuJSago71zQOszonAEv7oZutaLzJXmzqpwp9PKYu2D7isHAomr+1BzSG9+lWHehBi
xFqEu/NQRLUj1x5dOhG92pMvJwjNG14TGITTzCntYFz3hxV80+KVjxsNKal6BeU3oN3girHVpTHQ
+BaIr+VgL75CpYZ1R2eQp+ozhXlsxi5v5Uce5k9IUrBiav9Yp0PVF4bHzSlEsNm/6ZmcEh7Ff+Zz
ynJIwBEwsXN7JMwvAPxSKhOak1i9XuWHnZzzr/uoA/QYDHiYYKVzSiBF0UC3LRASqikX81VuEwcJ
7RsFDTR06g9ClhCg5MO8oWwn9drOdxnca8r9FSIXdetwJn08PHVdHhR6h3v+h/oZhIZ5lC54OLSx
tpbUu2vnzKCOWZ4+K0jfpFkHywJjDayuYcyZeM9X2QbpNNCfuyKJplcgdkASAwjkwF9MB4c9tgmY
S8OeXVUtXsTTlSPbU7hIljHrBJu8dxju/J53jwBIJjKEAolU/3h5PLKWsWXZEcWnufqLp+JNQxvz
HTJiekOXbhVAUiEUgYGRrFdPS7HKpxpPO/ff1JplECD13AL2qV+26uvfDM11cS4yIzAfaazY5lXe
Zsn1kosZ62uEYcj6b5ybqkST0xpZGkbc1Cwq4ymSka7yZ6BV622kW8Ke65zU+RqJeg9w0TX9D2cr
p/qJVGFb538Nq0bwS92smDOpjZNBfYqZIE7jbxWnjgyLuSDLLlUG1xhuBRkT6c4kj/cUAXTRn1LF
9OZ2IME25JorttPW09tMXRuePvbSFqW4ihjB0XlJ1k2a4pCCbrAZqonn3m5Tq9aGpWInVSaQQwfD
/eY4IWbJWSnHen7LWLfU664j2Ieb7VSbP92oBZycJFRwkRVxJLWhLm125RlxuXP6uxOzAfz/vuzA
FmIoy/7OiNWr5iuGTDopALwpN5s1XVG8CGFg8zGhFtKG0q/7kpFIjAl6n6J7WRsg5tjhczZ5rEhj
AfAaTA3sVriMu8XM5qAtPwm+W/4ZiFSseB+0pL2It2fcz3G2EjpIJZOS6pwr+1+HoYBVEoggBJ+X
eRsgWFJR5x25A3D7UmUPB3Zv3QzFIRK/PgMJpz/2vrzLPLuV31HDdRWKEgeIXd287dFIyJb2l9JA
X4cQIpMTeLJbTWnFEm3H++qA4hXgRXdiOHiKHybAMDGb0ZgB17Q2Rz2wFLc3uBZHNI/u//tUHF64
qM2hztzMCWX3RbLGjIz8dtfSmeuFMg+CY0nKb9yZBFsTQmzUjqSn2FHoWzG8tE1ZxDUBW/SFv8NE
10YYnc3L/w/Epn18yvJFiu39oWtG3qCe/dA43anY+YCW0hLHJ/WcP7EKxTDsAUndT7rCDC9z0NUy
g65OBKJwiCsou1tjad5Kd0X8fNTuSSjiHwjOwh4HCGHg9TrAV0xiqgPrW0p78IAc4qgiMmYuuzqm
ias/aVvaeief2mbw/FFfPvGmigEhaT4opn7CHXUElcWv9EUORKIQuZeXa9WfgoKHl57vHBnpGWTA
OcAvEmgWAr+gEsYuSn9RiLvBP1ZgB6tK8sng0vOCLFrM6vFXZWsSxCsgYXfOwEiyOrqgx7IftMeN
S//Pj5ZL5Oqr78P5+Tn9aYw04J2ueRdsfxMPnRb1iw2NvYftHYfMkntQihzEZlKIjfUi67lxjihV
iWI8M83xftVVpftqkARGbvH6JrrOHeJabAzB4n+GN+w9LjBDgX1bQ4+K/xskLeIoJcXQhZSmC/8t
F2b7cPP8pY4AhQAav41eXAT0hxk2lpfFrLropYNrcEo3wtQbZxjfqGwzhHKpiMuE8ruQPe7DlG4p
QOrfFgBn278C8eM5/OtB7+SHCL7gmof0AG+D73E5FsF8ImG5VVPC/qphNHoeMAqc8JbZ5BbkpUny
Y4wzBKEY/pVY7qAwAXZgIdKZy7i3r5NNxla2maLPeGmGeVGBiKDfkgKhpSxFk9EsTtzHoE495tbo
PQJ3IM8tkOsmBTffeoZyWj3X11zcCANMRS9WL8C9nVWkom1jw30W1+BKoZBJCys+F/nb4Gnngh+W
JZ1c2WGYOlhmC0kfEFRrIJboB4TQcz8sqKJrWg5mEP00mRpIa0pNCrz8DqZqryx5alpjChLNodx2
NT3J1MyHku57PNcFTk3N4564/Xwhg+TmwkqRCK5uijaEQaNOrobZl4wiwfac1SNk72z7NWLcd0Gt
5jqm6EDQ7ui/KMGYBsRJAWaJove/zrM54Rucgu9fNoTyCGHfgH/Uo50/1wt1AU4L5kEAQxomQ4Pe
oMaiMymO583MvumQCukSbj18uHN4onrfu1cETD1r0dV3z9n2XMwhSVbHdU/GK2QdWpQLkUHLTUOZ
jEibWldThmzn0FIR+N+tN1satIF38HrY5OptceXGbzrIQeyzn7jHblW28V7XofUShAbCEsrn5PGr
SWfOU1bo9rKsjSF+uhQm6IkKbESm8dp7W+7s4qrwkHF94RyNT/t+2vhAaFe4mmUjEcw5Phklp6Jo
0AALrmdaQdy/T9p95QIlpuubRaTvCTCP8HckI+od+mIRNllzrc4urNuiUXij2jC4RcngedhbNCiS
RFeVz5B7yxcJytA/YzSzgpQwdDVRmeaXZk/GDeuB5i1kSg4e2ley67ZVquK7+9nz1FMVHDX3WLMo
XAZNaJ9qJrz/3DK+3b2mZIJ35gZFm+HyaPc+YkLb53zAwqjxIuir6yoyOkoXETHASaZNxndosdXw
HMeBirjvYHgNvYkVeI4QUyVIE6S4X/cHhVRL1BREoTyNvJEyLUM//xRDPvhawM7Ej2wyX4pJ+UJl
lYPAtocz9oah0CJTyvOawAP74GcAz10PN25U86wh36+GM6EAVHlbuj398NccAiO5fQwsPwNgmGpT
sCuEv9oCZrzqp50QivSk0Eh2Wi6UJFU60/zOhrH7X9VTO/7s7hwXI1jvT6NTRS6Z6MH3XcLigXZa
oX//X2Ky/0Y4QyXXBtA4ERUvcBEvg6Lf/HSH0sAM18ZuBQ8mRGcmMMQntNoENrnQ+HCBNIpZfw5t
uoSrZIU1EhanHECGqKZA3LNSL7aRIitosPOKBMtqWcXoW+A0vT39aYQI0eAAmk9bDto8DnOKfg3I
fQm37xJUR42GIyw5rnNJ/13i/HSVaqDy3XA8kqjyVDs7izxzBJ4RZ7RekAWSCQGPOpII7vdE/w/W
eKWTiMLt7kDShZHQ579ojjnjoNzAuBxF4N1YCw9v7ZWOdwvJHKZSOtnFT9rdyiIKHKKhaCA+rczq
tledAefcJSu0rjwt4Pny+aRZjjeq8vFSMhEPG82GlbeRDWfy6bvvuJQuj9+A6b4xdauenqzf/Y+W
btE/Wlq5mTPMWk1HJ0t7PISXdK9SBVbpP63YXg2jfnEfW+2cAh+l3c1CYlzPGM/MtS1qQVh7o5/J
IJ0mk/K8SKUQsu31V5WPPlxnfhiovLh66JmkJSuT8fYPW+8JOdYvJ3SipOsYyzy6hNY7efDF/vqT
j9A66/GpJT5ShADb/u/O6f2wXeNN7nH7b6va9i3NMgi28wV+iUsGWsRZGNjNTENWjusQUhnaGtxB
709LS851PiuaFQHwpxYSeQMrGPC6L4MlDC3pQM/0BEJzRHDoYeV7n0j6vXjqtzcVs8sObUGxeyT+
nRphaMTdNqm/4fHiA0R6VbFGivF5W2btC0VT4fkqX8ORBQNM
`pragma protect end_protected
