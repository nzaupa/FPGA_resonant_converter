��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�=D>�ͺ��z�E�����D���2"��Nތ�3O�w���P�
��g���U���W(k�fL��2����P�Ә�yт6�K����q�n�˫�����eIX��£d5�(��h飂6�,�l�g�����;���J� TkЯ�Lr�?j�E$������s���%�MT�(�y�Zĺ�	��x,52�h^��}��E�~k$�?�ʍErd'�J����b� ��W���t���J-�fB|��OQ6;w�������B�hb���C@�l��j��P���E(���N�crEC�� �
J���S�{�nA�g�ScȀGM�̖{v�D��a��_�e�v��-�G�Jf	K���K����nLi�k;^��/����T����ʎ������ Mۑ���^�6��?*U� w�p;�6��X�T��m����<��I��#�^�o��p9�/O��`����WNm�P�{W"����&��/�A��\[�B��t5>ڴGcg:w6~2�[H<����F��?�ޓ�߶G�l��@�f�_��G�f,��Γ)$�"Ib6U0�Re�ʰT�74Ƀ�A	�"L,��EwoѦP�:<,^8�ѭ
�B��nxn�)@�DyY��������G�V�[�G���˖����"�X�R�>Va��"2lG�6�2���PP��ޝ��I�ިVޙ�l>��;3F���Ҟi�D��su�B\J�*Ō���=��f�g���		Ku�J`Q%ʊ�NeW��a�����qiޗ����s0 �0���3�iˊ���{5��)t}I>ƌ���{	��zQ��h�f�I���.7�U�r��o������Q��"ܚM��i�{�rs�ݓ�|�6��E�]���~����z�v�:�̼ۭ�I� ��&.G�GG����L���9�ؑd����8)JP��aFꬎ�g=2���'���}����j�s!wG�e�._�������ݯNc��o�M ��A�jL3�������g�pg��h�4���_�{ρ�/��WŶ�K$V�_ߩ(���`{
ił�B3��c�\����y�aGN��3��*V��T�VR��s�/���Ǌ��<+��jPޠgTLmL)�ʽ�I]�='�};G䚺�ㇳ���<d�"��5��Z���pt����
�\ͅ��Y���by!�ǆ3�`�xtExܫ��V��`�%h��g��Yn�Y�.��QZ�=��I-o��*�~�HG:���PZM�����d-
��Gmn!3o�2����������a��2�U�Ю<�,,P3 �Pue�Z�I߬l	������]�ۣ"=�42�r!��]��܆�pZ���v�x\L>���fj5=>�J��������������k��jߊ��������l�
de���?�p�d��d�0�ӆg��(�lح\�P�=�ӘO�O�Z4R����a�\�Y�鿻%�,9E�В�w�q���qXz�Q�Ǳ�����GLL��3e�i�:�À _����VR��+���Iu+s�Z�l���U�����h�ԧ��:��pԅɗq����N�&�T`^�i��B�U��L"VQ�L:��;��H��H,0�S�A3Ւ��>��s)"��n�#u��~�`�'�k_�ZO��e�Ջ��@�s�>�������j�K���y)a�?����߼p����/�o��Jf��ө)����KH;h4<b��O�._,�=�EӜᵶ�0���T䉡���qQ��B+����R�Y����������)�rZ�q�8�ִ-�}�)"�cOT�_V��aU�h� ��|���
=���J~�k��-o4��f,Ū��_Z�dg�o��|��i~�&�r��m�Jݫ�geM�>Y�~��+A�pc=��|���B����Ӓ��ۗ�8fM.4�@RP�H�XE�Y[F6w��ܔ�������9��3�0	AҖ<�]>e�����ԛ�z�ݨ�|^�9��<�3yz�`&��� �5~۔���A^�7��x�Z'����b;,ܵ��jG𼞐i�"����"�Pi��YO��[�6���U K?��d�O���^�wc�1�@ڝ�*W���U�V=^+I��B֝���s��ݢp� �ϸ�Ŕ�����>��aEg��`*ͦ0����^��4(bI�C�AB�%���n��aD���{
 �gW@�)�j�vq�#��6s슼S�,��@:}䫭��d�H�tK��ï�m�.�Sy�-Ov�����ӭ�"Z�\%j��>��m�Z�.��i�˰' KMG����W�5s�$b��"L�J�o�h����� d�N�%�����?0$�|�g6°7W�`��
��X���~�8����L8��<RL�T �u�gi�4�U��=������e�I��_Q��i�tvd7o���G�}��Ґ�
��̼ ��?���2�k�_E�B^]$��\-~�.��_ �5����������t�,���z���B��t;Di, n�,`>mF�����L��ڢ��ݻ�PP �,����R�����8�*��)�1�0x�p\��C�J8��LwL���p.<�~��H��J{�����Cb~Ʒ��\��D�z�|Wj�0�No�r�;��.����C��FkUn'��~�Vg��l�wZ��−�l�C|oU|�o�bधk��$z����1�R��N�5a���6X�C:a5[%(Α���ί��pi(�Pmۧ����C������H� �eN�emZ���*7��O^�ǲZ���� 3����}���&!j���- ��qmz����B|T"�lYg`�	�f��z�΄
�`�m��O����OGt�ؠ/���u`��DX���n�J`���\,DO�{�g?�Z��6j��:L=�1ߒr��:!�$v���<<*zN�,��{0f�	]��K�7
p,cnػȞ�޿D���Y�����uÒ����l#����
�:�g����\�3�M��*�0w2�F`x}�*�"T'�ޮ�-���F��MJ����<#��[�����24����,1��T�ӻ�s
�ށk�m� 2�z�yt��p"���|��
M� �0��-�����
8�Rd��|u�^7��7R��hxǑ�^6�f��'_�	�$�-�'�I�5 �>#��7�j��f������v�efz�͕��Q7��/�{�~��}v����E���G�,�ƭ��٩�����������L�ҷg��֌�D�|�T����秬�ӥ�;�Z{~Fȸk4h1�n�b�ߺ�:q8����j�>�����WiuΏ"9�$�]�)��5Q���xW��!�I#
k��V^��-��tT�hǴU�Х&�p��ig'�� f�hN�����N�Eө�-�{@�|�y��ˉ�ń�Q�wʷ�6��:���8����ʃ7�{4&LҮf4=7j��Ƶ���x���~�~���Z����k��(m�g%����V���ZJH���ʿ�� OL_�F�V	�ɎҖ�n�Ir�;!�ޭ,����N�m���#[�e Pܻ��7�~WJ� _��.$W9u8hy�z�=�m�W�R�a�R���%%��Z��}����7�gc}2�`�z6�3��xӿ�G�c4��p}?��)*�\��XP��]�Ez�8aa�R�q!�IRi�ĥ�;*g	��s�a�&�@y�9F�W٪�{�����q��[�B�<����s�o�;)�l�Q�ޓ:5�/(����p]S<�ة�֜�@ (]%��z�c\s}|�h���I��^n"d(�7�̌P�ǝ�Bp6>?�(��L��?4���R}�ĹU�1�j���Iuf�I-�@���&�����'�;��8A�&5�n�^6=ϝ�4\~̎ �>wle|�՛���2Sm�
$n�o;�/(+�VZ�0Zvi�u�}�@�5q܊�ܠ*Z���7`\��n7���ص}"�÷��/��a3]�P��Y�q�u)I��sw5\����o��爯�*��{�!e���}�l�i^V���N��jr�w�+��؂������~�r%�p�+t��?mm�_/w�b�=-��U�����j�\]Ҟ	�%|EY�$��a�|w�Ԏ���B*�2�/c�tm���9��Tx�Fq�Aπ��&T:/I��ϘQӵ�ER�8d�ᯫKb��� [�/Q���ɩ�%�:�V,7�\Y�d7�7�q�)E��؍��Q�GK�|� 3��J ��nӃ����/�&���~��'�U��?�o5�W6��&�(N�\�b=��l�X�a�a���S>��=�� ��q�:wb�%b$^b,3�����*�*�!�'�LU@�A�TQ&�2�5�%�B��