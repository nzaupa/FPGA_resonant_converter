��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l��ӡ;h�>�s��j��=U�߻*"���A�T�t(��05Y-٭!�Iu�Q7��|C}�r��b�}�l{�����8r$P�14eWw�Ϣ:ej�)���Ӕ[��T��
I�3.d�'A8��-����g�kW���ڇ�����,���0���N:�Zd2�W���!���	��_�1%r���Ҩ41¹]�a Oć���','�p���Ew�û�ܟ+��B� :]��O�O�������t!�O����lV�.�<7CJR�^����4h^˼�b�]��rc��"�0�Fu0�u!��Zpո/g�E:�0�[ Z�Q5�,���(5�O#Q\��E�����d���ĝ�W1��Rbv,�K��̬Jܖ�k���Ye�2]B�.2��5�����A��F�������q�f�E��`��ǥ�� �'vNɭɅ���	BB�D!��ش�o��7>����U�'E,'*���'��,����I<s��2ُ��@�!�]wy��ݘ�?���wߦ���d�:H�B�F�_����H��`�
t\���W�+�H�R� ]�0&�|"�^���\�me/���r�\����@�o��ZJ�>:A]�"�ހ+a�K�(���g�L0�׌Ɓ��.����%��m��b� �5�ٻ^�as ҩ3��f#�;�Yw��w��'���q�B��i.���Nð=�I9��[6&�W���M۫�V(� /	��T �i�{��Ba��^��Ό��~9ۃQ�~} '��ӌ����wZ�,��A%�;ۉ@(Y��������bR��N����Բ��9�SE6Df�Sk\|�$6�4��A���gC�*��/�:�/`��F�����~i��_@е1�G�2���Љ�\i�@59�Z#-K�pYuc��[�N	ǆ�1�1���̌Bc�ٴ@8~m�N�?��m�3�&�RC�'6TRb��!b�j�|��c�KEt׎K�R�w�y��lkbof��o响���tbI)�̸N1�{oJI7	y���iqQ9�"�+V�Е�p�k1=������c2�vl$>����/����D�<��.�.
Jt1J��2+�M`�y�(�+撖����n-</��f�""�f�&ʑ,�vyo�4MY���O8�,��Z�g���p&�p&X
r�Dq�������rx����7HI��>е4&�-(�U�"�JR��Ѥ�9�K�j}e�\ǟӟr�'/&���.R=�1r9�������9�8�9��o@6�8�1�� �^8������i˼ewU&���-g��w�|��mV	x1�+���+��YI�:P���^q�u�$2F@y�w�!`�r�gX��"���:ʸ3cobW{�;����E1��jcM}�gp��Ѡ:�KQ�m-�vt1�h�a����Po��'�����,P�c��潎�_n�w$.������&0q!\����k�cl�@�|ۓ�U�)��p�B�f�cu�a8r���n�/��*���q�@`
������C���
T��(<���z��q��oSD�I�͛�F�i>~8�e�}��E�g���S}��+���s�]:Q�����=���Т��"4ҕ��6�-�I�œ��(��NN�wa(��ΰ /�atu5H��Q!ۡ	oj�n�Rd�g�:��v��;{ӥ��n�<�-#�u�D �\2:�N�L.�����&��h]b�� y:L� FK^]P�:��1|ʧ��l�Զ���{r�!J���ہ�\!�ύ�ߍV%](�XЂ�0G{�WWu�̩+�6�hI��	7�@�4<n8��F�3Y}��&����We7�Ⱥ_��5��_��,�--���;p$��8E.NxH�8L��J������4V�?������UW�U��K:�:�e�*��-s�M��{k�n���@�����Chϳ�g�6�1�Asn��h�����'�&P�>*���q��"w�=J�<v��@��@l�z3'�挭��k�����%ժxV�N�~��b7z񽯙���SRb����n���y�w��J���Y�;��\'P>��; FC�D�0�9�{@R:<��{H��b���	�)����H*��d����� M;+��,�\q$S�X�&��Y�>hJ���� ��Ds�[I"�辐kt��]G�OQ\e�����<z��M��5��l�?�2<}��H��������[��"13��~�S�RQ�i���/�QQ�,�<� R��bLel�L���f������R��<��qE�BS�MZ���Tlu	��a��9ٲ\太��t)��3Q!�2�DsJD�X��;R�L8Lk�*�^�S�6e�ܼ��{�m�ڕ"I~n�Yb�Q�)4��^/��u_Y{h�;��t1�-�EJM,f�	$�ˬ�@��״��D�a�8^�'8X�y�׊�(��C�'^17A�+[>}0H�knER��P�������z����+��>8�/��@ֳPJ�|�_�56Ҽ�t���?��˅@|Sٍ����B�"NA;e�t��C���qu�ͺ�m��H��L[F/;�|��r`��
r��P	��_���~�c�:QU$k��By�b%��$GUE$X�y���V!�ڢ��uѕ�A��s@�T�%���N���y8��i��ƭ����U��(^˺t�^����(E�хc�&Ɂ܀6�z+�-.��-\\����f0��1��P���;�M6����0�zc
��M�>�W����,�v�io��+9����/�C��������mMP���7�}�ܯ'�cv���LP�U�1��Ia��'�2��h�Sg%}G�$F&E�;�}�yCeQNN