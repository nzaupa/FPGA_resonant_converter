//------------------------------------------------------------
// Project: HYBRID_CONTROL
// Author: Nicola Zaupa
// Date: (2023/11/08) (16:19:35)
// File: tb_hybrid_control_theta_phi.v
//------------------------------------------------------------
// Description:
// test-bench for the simulation of the hybrid control block.
// The idea is to test the proper operations of the state 
// machine.
//------------------------------------------------------------


`timescale 1 ns / 1 ps

module tb_hybrid_control_theta_phi();


reg clk_100M;
reg [13:0] vC, iC;
wire [1:0] sigma;


// call the block to be simulated
hybrid_control_theta_phi #(.mu_z1(32'd86), .mu_z2(32'd90), .mu_Vg(32'd312000)
) hybrid_control_theta_phi_inst (
   .i_clock( clk_100M ), 
   .i_RESET( 1),    
   .i_vC( vC ),      
   .i_iC( iC ),       
   .i_theta( 32'd165 ),   
   .i_phi( 32'd5 ),
   .o_sigma(sigma)
);

// call the block to be simulated
hybrid_control_phi #(.mu_z1(32'd86), .mu_z2(32'd90), .mu_Vg(32'd312000)
) hybrid_control_phi_inst (
   .i_clock( clk_100M ), 
   .i_RESET(1'b1),    
   .i_vC( vC ),      
   .i_iC( iC ),       
   .i_phi( 32'd5 ),
   .o_sigma()
);


simulator_LLC #() simulator_LLC_inst (
   .vC_p(), 
   .iS_p(), 
   .Vo_p(),    
   .CLK(clk_100M),    
   .RESET(1'b1),   
   .sigma(sigma)
);

// create the clock signal
// always begin //100MHz
//    clk_100M = 1'b1;
//    #5
//    clk_100M = 1'b0;
//    #5;
// end

initial begin // generate the input voltage and current

// samplings of current and voltage


clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110110; // iC=   54 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011100; // iC=   28 
vC = 14'b0000000001110110; // vC=  118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010000; // iC=   80 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100001; // iC=  161 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111001; // iC=  121 
vC = 14'b0000000000010111; // vC=   23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110111; // iC=   55 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101010; // iC=  170 
vC = 14'b0000000001010000; // vC=   80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110100; // iC=  180 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011101; // iC=  157 
vC = 14'b0000000001000111; // vC=   71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011010; // iC=   90 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110100; // iC=  180 
vC = 14'b0000000000011001; // vC=   25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010110; // iC=   86 
vC = 14'b0000000000111111; // vC=   63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110001; // iC=  113 
vC = 14'b0000000001110101; // vC=  117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101000; // iC=  168 
vC = 14'b0000000010010011; // vC=  147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000011; // iC=  131 
vC = 14'b0000000001110111; // vC=  119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111111; // iC=  191 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010110; // iC=  214 
vC = 14'b0000000010010110; // vC=  150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111011; // iC=  187 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011001; // iC=   89 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001100; // iC=  204 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010011; // iC=  147 
vC = 14'b0000000000111001; // vC=   57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010001; // iC=  209 
vC = 14'b0000000001101111; // vC=  111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111110; // iC=  126 
vC = 14'b0000000001110111; // vC=  119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010101; // iC=  149 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001001; // iC=  201 
vC = 14'b0000000001101101; // vC=  109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011111; // iC=  223 
vC = 14'b0000000010000000; // vC=  128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111100; // iC=  124 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101111; // iC=  239 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010010; // iC=  210 
vC = 14'b0000000010000101; // vC=  133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110001; // iC=  177 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011110; // iC=  158 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110000; // iC=  176 
vC = 14'b0000000000011000; // vC=   24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001010; // iC=  138 
vC = 14'b0000000010100010; // vC=  162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110000; // iC=  176 
vC = 14'b0000000001110010; // vC=  114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001111; // iC=  207 
vC = 14'b0000000010001100; // vC=  140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011001; // iC=  281 
vC = 14'b0000000010000000; // vC=  128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000101; // iC=  197 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001010; // iC=  138 
vC = 14'b0000000000011010; // vC=   26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001011; // iC=  203 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110010; // iC=  242 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011001; // iC=  153 
vC = 14'b0000000010101000; // vC=  168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001000; // iC=  264 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101011; // iC=  299 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100101; // iC=  293 
vC = 14'b0000000000111111; // vC=   63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101000; // iC=  296 
vC = 14'b0000000001010101; // vC=   85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110100; // iC=  244 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100101; // iC=  229 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100001; // iC=  161 
vC = 14'b0000000000011100; // vC=   28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100101; // iC=  293 
vC = 14'b0000000001101000; // vC=  104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010101; // iC=  277 
vC = 14'b0000000000100011; // vC=   35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110101; // iC=  245 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000000; // iC=  256 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101100; // iC=  300 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111010; // iC=  250 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001111; // iC=  143 
vC = 14'b0000000010001100; // vC=  140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100010; // iC=  290 
vC = 14'b0000000000011111; // vC=   31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110111; // iC=  183 
vC = 14'b0000000010011011; // vC=  155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001001; // iC=  265 
vC = 14'b0000000001110010; // vC=  114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011001; // iC=  153 
vC = 14'b0000000001101000; // vC=  104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101010; // iC=  298 
vC = 14'b0000000001000100; // vC=   68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100010; // iC=  162 
vC = 14'b0000000001111101; // vC=  125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000001; // iC=  193 
vC = 14'b0000000010010011; // vC=  147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110010; // iC=  242 
vC = 14'b0000000001110100; // vC=  116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001011; // iC=  139 
vC = 14'b0000000000011111; // vC=   31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111110; // iC=  190 
vC = 14'b0000000000110000; // vC=   48 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011110; // iC=  286 
vC = 14'b0000000010001110; // vC=  142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100001; // iC=  289 
vC = 14'b0000000001011111; // vC=   95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010100; // iC=  148 
vC = 14'b0000000000111000; // vC=   56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000010; // iC=  130 
vC = 14'b0000000001010000; // vC=   80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001011; // iC=  203 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111011; // iC=  251 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011001; // iC=  281 
vC = 14'b0000000010101111; // vC=  175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011111; // iC=  159 
vC = 14'b0000000010010111; // vC=  151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100000; // iC=  160 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000000; // iC=  192 
vC = 14'b0000000010110111; // vC=  183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001101; // iC=  205 
vC = 14'b0000000000100001; // vC=   33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111100; // iC=  188 
vC = 14'b0000000000111000; // vC=   56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001011; // iC=  267 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110011; // iC=  243 
vC = 14'b0000000010001001; // vC=  137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111000; // iC=  184 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011010; // iC=  218 
vC = 14'b0000000001110110; // vC=  118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001100; // iC=  204 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010011; // iC=  211 
vC = 14'b0000000000100110; // vC=   38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010011; // iC=  211 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011111; // iC=  159 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101011; // iC=  171 
vC = 14'b0000000000100011; // vC=   35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001110; // iC=  206 
vC = 14'b0000000000100100; // vC=   36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100100; // iC=  164 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010111; // iC=  215 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010110; // iC=  150 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110000; // iC=  112 
vC = 14'b0000000011000110; // vC=  198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101010; // iC=  170 
vC = 14'b0000000010111100; // vC=  188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110111; // iC=  247 
vC = 14'b0000000010100100; // vC=  164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110111; // iC=  119 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011000; // iC=  216 
vC = 14'b0000000010110110; // vC=  182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001010; // iC=  202 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100011; // iC=  227 
vC = 14'b0000000001101001; // vC=  105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010000; // iC=  144 
vC = 14'b0000000010001001; // vC=  137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100001; // iC=  225 
vC = 14'b0000000001111001; // vC=  121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001100; // iC=  140 
vC = 14'b0000000010001010; // vC=  138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110010; // iC=  242 
vC = 14'b0000000001101111; // vC=  111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111001; // iC=  185 
vC = 14'b0000000001001110; // vC=   78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101010; // iC=  170 
vC = 14'b0000000010000001; // vC=  129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010111; // iC=  215 
vC = 14'b0000000001011000; // vC=   88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110111; // iC=  119 
vC = 14'b0000000000101000; // vC=   40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011011; // iC=  219 
vC = 14'b0000000010001011; // vC=  139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110001; // iC=  241 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101110; // iC=  110 
vC = 14'b0000000001110111; // vC=  119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011011; // iC=   91 
vC = 14'b0000000001100000; // vC=   96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100000; // iC=  160 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111100; // iC=  124 
vC = 14'b0000000001111010; // vC=  122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010001; // iC=  145 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010001; // iC=  145 
vC = 14'b0000000010001110; // vC=  142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100011; // iC=  163 
vC = 14'b0000000010101011; // vC=  171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000101; // iC=  197 
vC = 14'b0000000001010111; // vC=   87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100001; // iC=  161 
vC = 14'b0000000010101100; // vC=  172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000001; // iC=   65 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001011; // iC=  139 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010100; // iC=  148 
vC = 14'b0000000001011010; // vC=   90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000001; // iC=   65 
vC = 14'b0000000001000111; // vC=   71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011000; // iC=   88 
vC = 14'b0000000010010110; // vC=  150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010100; // iC=  212 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111011; // iC=  187 
vC = 14'b0000000010111100; // vC=  188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001101; // iC=   77 
vC = 14'b0000000001111111; // vC=  127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010011; // iC=   83 
vC = 14'b0000000010010011; // vC=  147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011101; // iC=   93 
vC = 14'b0000000000110100; // vC=   52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100100; // iC=  100 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101000; // iC=  104 
vC = 14'b0000000010111101; // vC=  189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111011; // iC=  187 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111000; // iC=  184 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110010; // iC=  178 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110111; // iC=  183 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011001; // iC=   89 
vC = 14'b0000000010010111; // vC=  151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100110; // iC=   38 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111101; // iC=  125 
vC = 14'b0000000001111010; // vC=  122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110010; // iC=  178 
vC = 14'b0000000001101100; // vC=  108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101010; // iC=   42 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111111; // iC=  127 
vC = 14'b0000000010000000; // vC=  128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011011; // iC=   27 
vC = 14'b0000000010111011; // vC=  187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100110; // iC=  166 
vC = 14'b0000000010011110; // vC=  158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011001; // iC=   89 
vC = 14'b0000000010101110; // vC=  174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111111; // iC=   63 
vC = 14'b0000000001110010; // vC=  114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010100; // iC=   20 
vC = 14'b0000000010001101; // vC=  141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110000; // iC=   48 
vC = 14'b0000000001011100; // vC=   92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011111; // iC=   31 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110100; // iC=  116 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010110; // iC=  150 
vC = 14'b0000000011000110; // vC=  198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100111; // iC=   39 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000000; // iC=  128 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101000; // iC=  168 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000011; // iC=   67 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001011; // iC=   75 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001010; // iC=   74 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001001; // iC=   73 
vC = 14'b0000000010000001; // vC=  129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010110; // iC=   22 
vC = 14'b0000000000110111; // vC=   55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110001; // iC=  113 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001111; // iC=   15 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100011; // iC=   35 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100100; // iC=  100 
vC = 14'b0000000010000100; // vC=  132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001100; // iC=   76 
vC = 14'b0000000001110101; // vC=  117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111111; // iC=  127 
vC = 14'b0000000011001000; // vC=  200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010001; // iC=   17 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100010; // iC=   34 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100010; // iC=   34 
vC = 14'b0000000000111110; // vC=   62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000101; // iC=   69 
vC = 14'b0000000001011011; // vC=   91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000010; // iC=   66 
vC = 14'b0000000010100101; // vC=  165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001101; // iC=   13 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110001; // iC=   49 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000010; // iC=  130 
vC = 14'b0000000001011000; // vC=   88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111001; // iC=   57 
vC = 14'b0000000001100111; // vC=  103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101001; // iC=   41 
vC = 14'b0000000000110101; // vC=   53 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100100; // iC=  164 
vC = 14'b0000000010110001; // vC=  177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011011; // iC=  155 
vC = 14'b0000000011000111; // vC=  199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001010; // iC=   74 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001110; // iC=   78 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000111; // iC=  135 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101110; // iC=  110 
vC = 14'b0000000001000101; // vC=   69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000010; // iC=   66 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111001; // iC=   57 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111101; // iC=  125 
vC = 14'b0000000001110111; // vC=  119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000100; // iC=   68 
vC = 14'b0000000001111010; // vC=  122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101111; // iC=   47 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011000; // iC=   88 
vC = 14'b0000000001110110; // vC=  118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010001; // iC=   81 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000000; // iC=   64 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100001; // iC=  161 
vC = 14'b0000000010011000; // vC=  152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000110; // iC=   70 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110110; // iC=  118 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000101; // iC=   69 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101101; // iC=  173 
vC = 14'b0000000011000011; // vC=  195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001100; // iC=  204 
vC = 14'b0000000001101111; // vC=  111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010011; // iC=   83 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000100; // iC=  132 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101101; // iC=  109 
vC = 14'b0000000010110110; // vC=  182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110101; // iC=  117 
vC = 14'b0000000010111111; // vC=  191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000000; // iC=  128 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010000; // iC=  208 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011011; // iC=  155 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100100; // iC=  164 
vC = 14'b0000000001001110; // vC=   78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010001; // iC=  209 
vC = 14'b0000000001011101; // vC=   93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010011; // iC=  211 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111000; // iC=  120 
vC = 14'b0000000011010011; // vC=  211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101011; // iC=  107 
vC = 14'b0000000010000000; // vC=  128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000000; // iC=  128 
vC = 14'b0000000010011001; // vC=  153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100010; // iC=  226 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110110; // iC=  182 
vC = 14'b0000000010011001; // vC=  153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111010; // iC=  186 
vC = 14'b0000000011001011; // vC=  203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100110; // iC=  102 
vC = 14'b0000000011010011; // vC=  211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101101; // iC=  109 
vC = 14'b0000000001010010; // vC=   82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100100; // iC=  100 
vC = 14'b0000000001111011; // vC=  123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110111; // iC=  183 
vC = 14'b0000000010010110; // vC=  150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011011; // iC=  219 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110101; // iC=  181 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001001; // iC=  137 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101111; // iC=  111 
vC = 14'b0000000011001001; // vC=  201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000011; // iC=  131 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101000; // iC=  168 
vC = 14'b0000000011010110; // vC=  214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010000; // iC=  144 
vC = 14'b0000000001010011; // vC=   83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001001; // iC=  137 
vC = 14'b0000000011000000; // vC=  192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010111; // iC=  215 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110100; // iC=  244 
vC = 14'b0000000010100101; // vC=  165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001111; // iC=  143 
vC = 14'b0000000010010011; // vC=  147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110111; // iC=  119 
vC = 14'b0000000010101010; // vC=  170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010001; // iC=  209 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100001; // iC=   97 
vC = 14'b0000000001001110; // vC=   78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111011; // iC=  187 
vC = 14'b0000000010101011; // vC=  171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000111; // iC=  199 
vC = 14'b0000000001101100; // vC=  108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010111; // iC=  151 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001000; // iC=  200 
vC = 14'b0000000010011100; // vC=  156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100011; // iC=  227 
vC = 14'b0000000010001010; // vC=  138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011001; // iC=   89 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101000; // iC=  104 
vC = 14'b0000000001010101; // vC=   85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010110; // iC=  214 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011011; // iC=   91 
vC = 14'b0000000011010100; // vC=  212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010010; // iC=   82 
vC = 14'b0000000010111000; // vC=  184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101010; // iC=  106 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101011; // iC=  171 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010010; // iC=   82 
vC = 14'b0000000010111001; // vC=  185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100101; // iC=  101 
vC = 14'b0000000001001111; // vC=   79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011001; // iC=  217 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100011; // iC=  163 
vC = 14'b0000000010001110; // vC=  142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100011; // iC=  163 
vC = 14'b0000000010001100; // vC=  140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101010; // iC=  170 
vC = 14'b0000000010100101; // vC=  165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101000; // iC=  168 
vC = 14'b0000000011010111; // vC=  215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000101; // iC=  133 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010010; // iC=  210 
vC = 14'b0000000011011101; // vC=  221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010000; // iC=   80 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110011; // iC=  179 
vC = 14'b0000000001101010; // vC=  106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011001; // iC=   89 
vC = 14'b0000000010010110; // vC=  150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100010; // iC=   98 
vC = 14'b0000000001101010; // vC=  106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010110; // iC=   86 
vC = 14'b0000000001010011; // vC=   83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111000; // iC=   56 
vC = 14'b0000000001110110; // vC=  118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110011; // iC=   51 
vC = 14'b0000000010111111; // vC=  191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110011; // iC=  115 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000111; // iC=   71 
vC = 14'b0000000010010110; // vC=  150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101110; // iC=  174 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001001; // iC=   73 
vC = 14'b0000000010111110; // vC=  190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000011; // iC=  195 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010011; // iC=  147 
vC = 14'b0000000011001001; // vC=  201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111000; // iC=  184 
vC = 14'b0000000010110110; // vC=  182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000000; // iC=  192 
vC = 14'b0000000010100000; // vC=  160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011101; // iC=   93 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101110; // iC=  110 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100111; // iC=   39 
vC = 14'b0000000010001010; // vC=  138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001110; // iC=   78 
vC = 14'b0000000010111110; // vC=  190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010101; // iC=   85 
vC = 14'b0000000001110111; // vC=  119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100111; // iC=  103 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101001; // iC=   41 
vC = 14'b0000000011010011; // vC=  211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011000; // iC=  152 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011111; // iC=   95 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110100; // iC=  180 
vC = 14'b0000000010000001; // vC=  129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010010; // iC=   82 
vC = 14'b0000000010011011; // vC=  155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100000; // iC=   32 
vC = 14'b0000000010110110; // vC=  182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010101; // iC=  149 
vC = 14'b0000000001111101; // vC=  125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010110; // iC=   22 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010000; // iC=  144 
vC = 14'b0000000010010010; // vC=  146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100010; // iC=   98 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101100; // iC=  108 
vC = 14'b0000000001111101; // vC=  125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011010; // iC=   90 
vC = 14'b0000000001111101; // vC=  125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111001; // iC=   57 
vC = 14'b0000000001101111; // vC=  111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001111; // iC=  143 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010001; // iC=  145 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100010; // iC=   98 
vC = 14'b0000000001010101; // vC=   85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110001; // iC=  113 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011010; // iC=   90 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111101; // iC=   61 
vC = 14'b0000000001010111; // vC=   87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011100; // iC=   28 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010001; // iC=   81 
vC = 14'b0000000011011011; // vC=  219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100100; // iC=   36 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111010; // iC=   -6 
vC = 14'b0000000011100000; // vC=  224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010000; // iC=   80 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011010; // iC=   90 
vC = 14'b0000000011100001; // vC=  225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111000; // iC=   56 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000011; // iC=   67 
vC = 14'b0000000011011111; // vC=  223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001110; // iC=   78 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111110; // iC=  126 
vC = 14'b0000000010101010; // vC=  170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110010; // iC=  -14 
vC = 14'b0000000011001100; // vC=  204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010100; // iC=   84 
vC = 14'b0000000011011011; // vC=  219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001001; // iC=    9 
vC = 14'b0000000001011000; // vC=   88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011110; // iC=   94 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011011; // iC=   91 
vC = 14'b0000000001011110; // vC=   94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101011; // iC=   43 
vC = 14'b0000000011001000; // vC=  200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000011; // iC=    3 
vC = 14'b0000000011001111; // vC=  207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000100; // iC=   68 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111101; // iC=   -3 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100100; // iC=  100 
vC = 14'b0000000010000001; // vC=  129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000100; // iC=    4 
vC = 14'b0000000010110011; // vC=  179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110011; // iC=  -13 
vC = 14'b0000000010111000; // vC=  184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111010; // iC=   58 
vC = 14'b0000000010010111; // vC=  151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101100; // iC=   44 
vC = 14'b0000000011100010; // vC=  226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101101; // iC=  -19 
vC = 14'b0000000010110011; // vC=  179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101110; // iC=  110 
vC = 14'b0000000010011001; // vC=  153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100000; // iC=   96 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010011; // iC=   19 
vC = 14'b0000000010101000; // vC=  168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011001; // iC=   89 
vC = 14'b0000000011001011; // vC=  203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100011; // iC=  -29 
vC = 14'b0000000010001010; // vC=  138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101110; // iC=   46 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001110; // iC=   14 
vC = 14'b0000000010101101; // vC=  173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000011; // iC=   67 
vC = 14'b0000000010000110; // vC=  134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111000; // iC=   -8 
vC = 14'b0000000010101100; // vC=  172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001110; // iC=  -50 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011000; // iC=   88 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001111; // iC=   79 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001100; // iC=  -52 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011100; // iC=  -36 
vC = 14'b0000000010101110; // vC=  174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100101; // iC=  -27 
vC = 14'b0000000011000100; // vC=  196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001111; // iC=  -49 
vC = 14'b0000000010001100; // vC=  140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110111; // iC=   55 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010111; // iC=   23 
vC = 14'b0000000010011100; // vC=  156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100111; // iC=  103 
vC = 14'b0000000001010011; // vC=   83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111111; // iC=   -1 
vC = 14'b0000000001101111; // vC=  111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110000; // iC=   48 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001101; // iC=  -51 
vC = 14'b0000000001100101; // vC=  101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111101; // iC=   -3 
vC = 14'b0000000010110111; // vC=  183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100101; // iC=  -27 
vC = 14'b0000000010011101; // vC=  157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110000; // iC=  -16 
vC = 14'b0000000001011000; // vC=   88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010110; // iC=   22 
vC = 14'b0000000011000010; // vC=  194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000001; // iC=   65 
vC = 14'b0000000010011101; // vC=  157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110001; // iC=  -15 
vC = 14'b0000000011011101; // vC=  221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011010; // iC=   26 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011010; // iC=   26 
vC = 14'b0000000010100000; // vC=  160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001010; // iC=   10 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010010; // iC=  -46 
vC = 14'b0000000001100000; // vC=   96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000011; // iC=   67 
vC = 14'b0000000001010101; // vC=   85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100001; // iC=   33 
vC = 14'b0000000001000101; // vC=   69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100011; // iC=  -29 
vC = 14'b0000000010101000; // vC=  168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100100; // iC=  -28 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001000; // iC=   72 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000001; // iC=    1 
vC = 14'b0000000010110011; // vC=  179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101110; // iC=   46 
vC = 14'b0000000001111101; // vC=  125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000010; // iC=  -62 
vC = 14'b0000000001000100; // vC=   68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001000; // iC=  -56 
vC = 14'b0000000010110111; // vC=  183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001011; // iC=   11 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100110; // iC=  -26 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011000; // iC=   24 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011001; // iC=  -39 
vC = 14'b0000000010100010; // vC=  162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101000; // iC=   40 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110101; // iC=  -75 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000011; // iC=    3 
vC = 14'b0000000001011100; // vC=   92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001101; // iC=  -51 
vC = 14'b0000000010001101; // vC=  141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010111; // iC=   23 
vC = 14'b0000000011001001; // vC=  201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010001; // iC=   17 
vC = 14'b0000000010100111; // vC=  167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110100; // iC=   52 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101000; // iC=   40 
vC = 14'b0000000001010101; // vC=   85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001100; // iC=   76 
vC = 14'b0000000010001011; // vC=  139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011110; // iC=  -34 
vC = 14'b0000000001110111; // vC=  119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111100; // iC=  -68 
vC = 14'b0000000001011010; // vC=   90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001100; // iC=   12 
vC = 14'b0000000010011100; // vC=  156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001011; // iC=   75 
vC = 14'b0000000010111111; // vC=  191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000000; // iC=   64 
vC = 14'b0000000000111101; // vC=   61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000011; // iC=    3 
vC = 14'b0000000010100101; // vC=  165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000001; // iC=    1 
vC = 14'b0000000010100000; // vC=  160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100100; // iC=   36 
vC = 14'b0000000001011011; // vC=   91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111001; // iC=   -7 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010010; // iC=  -46 
vC = 14'b0000000011001010; // vC=  202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101111; // iC=   47 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001001; // iC=  -55 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010100; // iC=  -44 
vC = 14'b0000000010111101; // vC=  189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000011; // iC=    3 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110111; // iC=  -73 
vC = 14'b0000000001111011; // vC=  123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111100; // iC=  -68 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000010; // iC=    2 
vC = 14'b0000000010101010; // vC=  170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111001; // iC=   57 
vC = 14'b0000000000111110; // vC=   62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101010; // iC=  -22 
vC = 14'b0000000010000011; // vC=  131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000111; // iC=    7 
vC = 14'b0000000011001011; // vC=  203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100111; // iC=  -89 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101001; // iC=  -87 
vC = 14'b0000000010000100; // vC=  132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011110; // iC=  -34 
vC = 14'b0000000000111001; // vC=   57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000001; // iC=   65 
vC = 14'b0000000010010011; // vC=  147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101011; // iC=  -21 
vC = 14'b0000000001110110; // vC=  118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110001; // iC=  -79 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001011; // iC=   11 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001110; // iC=   14 
vC = 14'b0000000000110011; // vC=   51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001110; // iC=  -50 
vC = 14'b0000000010100101; // vC=  165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000101; // iC=   69 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111111; // iC=  -65 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000000; // iC=   64 
vC = 14'b0000000010110010; // vC=  178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101001; // iC=  -23 
vC = 14'b0000000010001101; // vC=  141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011010; // iC=   26 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110110; // iC=  -10 
vC = 14'b0000000010100111; // vC=  167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100010; // iC=  -94 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111001; // iC=  -71 
vC = 14'b0000000000101101; // vC=   45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100101; // iC=   37 
vC = 14'b0000000010001101; // vC=  141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111101; // iC=  -67 
vC = 14'b0000000010100000; // vC=  160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110000; // iC=   48 
vC = 14'b0000000001100000; // vC=   96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000011; // iC=  -61 
vC = 14'b0000000010100010; // vC=  162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110101; // iC=   53 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001111; // iC=  -49 
vC = 14'b0000000010011011; // vC=  155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011110; // iC=  -34 
vC = 14'b0000000000101000; // vC=   40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010100; // iC=  -44 
vC = 14'b0000000000100100; // vC=   36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110011; // iC=  -13 
vC = 14'b0000000001110100; // vC=  116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111000; // iC=   -8 
vC = 14'b0000000001110111; // vC=  119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110101; // iC=   53 
vC = 14'b0000000001011010; // vC=   90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100011; // iC=  -93 
vC = 14'b0000000010111000; // vC=  184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101111; // iC=  -81 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110100; // iC=   52 
vC = 14'b0000000000101101; // vC=   45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011111; // iC=  -33 
vC = 14'b0000000010000100; // vC=  132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110110; // iC=  -74 
vC = 14'b0000000001100111; // vC=  103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011101; // iC=  -35 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000001; // iC=    1 
vC = 14'b0000000010100101; // vC=  165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010111; // iC=  -41 
vC = 14'b0000000000101111; // vC=   47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110101; // iC=  -11 
vC = 14'b0000000000100101; // vC=   37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001111; // iC=   15 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011001; // iC=   25 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111011; // iC=  -69 
vC = 14'b0000000010001001; // vC=  137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100111; // iC=   39 
vC = 14'b0000000010100111; // vC=  167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011001; // iC=  -39 
vC = 14'b0000000001010111; // vC=   87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001000; // iC= -120 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101000; // iC=  -88 
vC = 14'b0000000010100110; // vC=  166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100110; // iC=  -26 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100110; // iC=  -26 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101110; // iC=  -18 
vC = 14'b0000000010000101; // vC=  133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101001; // iC=  -23 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001110; // iC=   14 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111111; // iC=  -65 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111011; // iC= -133 
vC = 14'b0000000001000100; // vC=   68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011110; // iC=  -98 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101000; // iC=  -88 
vC = 14'b0000000010000000; // vC=  128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100101; // iC=  -91 
vC = 14'b0000000001000001; // vC=   65 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001000; // iC= -120 
vC = 14'b0000000000101011; // vC=   43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100000; // iC=  -96 
vC = 14'b0000000000111001; // vC=   57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111011; // iC= -133 
vC = 14'b0000000000011010; // vC=   26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000101; // iC= -123 
vC = 14'b0000000000100010; // vC=   34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010100; // iC= -108 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100011; // iC= -157 
vC = 14'b0000000000101110; // vC=   46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010001; // iC= -111 
vC = 14'b0000000000111111; // vC=   63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100101; // iC=  -27 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110101; // iC=  -75 
vC = 14'b0000000010100111; // vC=  167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011001; // iC=  -39 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010000; // iC= -112 
vC = 14'b0000000010101100; // vC=  172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101000; // iC= -152 
vC = 14'b0000000001111011; // vC=  123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100010; // iC=  -94 
vC = 14'b0000000000110100; // vC=   52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101111; // iC= -145 
vC = 14'b0000000010100110; // vC=  166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101111; // iC=  -81 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110000; // iC=  -80 
vC = 14'b0000000000111000; // vC=   56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011011; // iC= -229 
vC = 14'b0000000001110010; // vC=  114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110010; // iC=  -78 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100110; // iC=  -90 
vC = 14'b0000000010001011; // vC=  139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010111; // iC= -169 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101110; // iC= -146 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101001; // iC= -151 
vC = 14'b0000000001101001; // vC=  105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100110; // iC= -154 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101111; // iC= -273 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101101; // iC= -211 
vC = 14'b0000000000101011; // vC=   43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101110; // iC= -210 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110001; // iC= -143 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100001; // iC= -223 
vC = 14'b0000000000101110; // vC=   46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011111; // iC= -161 
vC = 14'b0000000010001111; // vC=  143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001000; // iC= -312 
vC = 14'b0000000001110010; // vC=  114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010110; // iC= -170 
vC = 14'b0000000000101010; // vC=   42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000011; // iC= -317 
vC = 14'b0000000000100000; // vC=   32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000100; // iC= -252 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011000; // iC= -296 
vC = 14'b0000000000000001; // vC=    1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111110; // iC= -322 
vC = 14'b0000000000101001; // vC=   41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100001; // iC= -351 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011011; // iC= -357 
vC = 14'b0000000001101011; // vC=  107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010101; // iC= -299 
vC = 14'b0000000001110100; // vC=  116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111101; // iC= -323 
vC = 14'b0000000001111010; // vC=  122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010100; // iC= -236 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000100; // iC= -380 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111101; // iC= -387 
vC = 14'b0000000010000011; // vC=  131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110000; // iC= -400 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111101; // iC= -259 
vC = 14'b0000000000000011; // vC=    3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110011; // iC= -269 
vC = 14'b0000000001011100; // vC=   92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100011; // iC= -413 
vC = 14'b1111111111101011; // vC=  -21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100100; // iC= -284 
vC = 14'b0000000001101010; // vC=  106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111010; // iC= -326 
vC = 14'b0000000000100010; // vC=   34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000010; // iC= -446 
vC = 14'b0000000000000011; // vC=    3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110110; // iC= -330 
vC = 14'b0000000000000100; // vC=    4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111100; // iC= -452 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001010; // iC= -310 
vC = 14'b1111111111101100; // vC=  -20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011011; // iC= -421 
vC = 14'b0000000001101101; // vC=  109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110111; // iC= -457 
vC = 14'b0000000000001101; // vC=   13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110100; // iC= -460 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000001; // iC= -383 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110111; // iC= -393 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111001; // iC= -455 
vC = 14'b0000000001000111; // vC=   71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110001; // iC= -399 
vC = 14'b1111111111100001; // vC=  -31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001111; // iC= -497 
vC = 14'b1111111111111011; // vC=   -5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100011; // iC= -413 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100000; // iC= -416 
vC = 14'b0000000001011100; // vC=   92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110000; // iC= -464 
vC = 14'b0000000000001111; // vC=   15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101101; // iC= -403 
vC = 14'b0000000001010000; // vC=   80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110101; // iC= -459 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001001; // iC= -439 
vC = 14'b1111111111010101; // vC=  -43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000110; // iC= -442 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001001; // iC= -503 
vC = 14'b0000000000110011; // vC=   51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010000; // iC= -560 
vC = 14'b0000000000101101; // vC=   45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111110; // iC= -450 
vC = 14'b1111111111001001; // vC=  -55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110110; // iC= -522 
vC = 14'b0000000000000001; // vC=    1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010010; // iC= -430 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001110; // iC= -562 
vC = 14'b0000000001010011; // vC=   83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101111; // iC= -465 
vC = 14'b0000000000110011; // vC=   51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110110; // iC= -522 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110001; // iC= -463 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011101; // iC= -547 
vC = 14'b0000000000010011; // vC=   19 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111001; // iC= -455 
vC = 14'b1111111111100001; // vC=  -31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101111; // iC= -529 
vC = 14'b1111111110101110; // vC=  -82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110011; // iC= -589 
vC = 14'b0000000000010001; // vC=   17 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101011; // iC= -597 
vC = 14'b0000000000101100; // vC=   44 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100011; // iC= -605 
vC = 14'b0000000000000001; // vC=    1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000001; // iC= -575 
vC = 14'b1111111111010011; // vC=  -45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110001; // iC= -463 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010011; // iC= -621 
vC = 14'b1111111111010111; // vC=  -41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111011; // iC= -517 
vC = 14'b1111111111000101; // vC=  -59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010100; // iC= -556 
vC = 14'b0000000000001111; // vC=   15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010101; // iC= -619 
vC = 14'b1111111110101011; // vC=  -85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000101; // iC= -571 
vC = 14'b0000000000110011; // vC=   51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110000; // iC= -528 
vC = 14'b0000000000000111; // vC=    7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011010; // iC= -486 
vC = 14'b1111111110011010; // vC= -102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100000; // iC= -608 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011000; // iC= -616 
vC = 14'b1111111111010010; // vC=  -46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000101; // iC= -507 
vC = 14'b0000000000011000; // vC=   24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011000; // iC= -552 
vC = 14'b1111111111011010; // vC=  -38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111001; // iC= -583 
vC = 14'b1111111110100110; // vC=  -90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110011; // iC= -589 
vC = 14'b1111111111101011; // vC=  -21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111110; // iC= -642 
vC = 14'b1111111110000101; // vC= -123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111010; // iC= -646 
vC = 14'b1111111110111111; // vC=  -65 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100110; // iC= -666 
vC = 14'b0000000000010100; // vC=   20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001000; // iC= -568 
vC = 14'b1111111111000101; // vC=  -59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111111; // iC= -577 
vC = 14'b1111111111111100; // vC=   -4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101010; // iC= -662 
vC = 14'b1111111111111101; // vC=   -3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001000; // iC= -632 
vC = 14'b1111111111010101; // vC=  -43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000100; // iC= -636 
vC = 14'b1111111111110011; // vC=  -13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001111; // iC= -625 
vC = 14'b1111111110110111; // vC=  -73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100100; // iC= -540 
vC = 14'b1111111111000100; // vC=  -60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000110; // iC= -634 
vC = 14'b1111111111000111; // vC=  -57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001110; // iC= -562 
vC = 14'b1111111111000100; // vC=  -60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000111; // iC= -633 
vC = 14'b1111111110100101; // vC=  -91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010011; // iC= -621 
vC = 14'b1111111111110101; // vC=  -11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010101; // iC= -555 
vC = 14'b1111111111101011; // vC=  -21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010010; // iC= -558 
vC = 14'b1111111110000011; // vC= -125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010101; // iC= -619 
vC = 14'b1111111111110010; // vC=  -14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110111; // iC= -585 
vC = 14'b1111111101111110; // vC= -130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011111; // iC= -609 
vC = 14'b1111111111110000; // vC=  -16 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b1111111101101100; // vC= -148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100100; // iC= -668 
vC = 14'b1111111110111100; // vC=  -68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110111; // iC= -585 
vC = 14'b1111111111010000; // vC=  -48 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000011; // iC= -637 
vC = 14'b1111111111001000; // vC=  -56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001001; // iC= -631 
vC = 14'b1111111101100010; // vC= -158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111101; // iC= -579 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100110; // iC= -666 
vC = 14'b1111111110100010; // vC=  -94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110000; // iC= -592 
vC = 14'b1111111110101111; // vC=  -81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010100; // iC= -684 
vC = 14'b1111111110010100; // vC= -108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b1111111110001011; // vC= -117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101101; // iC= -595 
vC = 14'b1111111110010010; // vC= -110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101111; // iC= -657 
vC = 14'b1111111110010110; // vC= -106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011101; // iC= -547 
vC = 14'b1111111110000010; // vC= -126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b1111111111010001; // vC=  -47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100100; // iC= -668 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b1111111101111100; // vC= -132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000010; // iC= -638 
vC = 14'b1111111111000100; // vC=  -60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000110; // iC= -634 
vC = 14'b1111111101100001; // vC= -159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100101; // iC= -539 
vC = 14'b1111111110111101; // vC=  -67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000111; // iC= -569 
vC = 14'b1111111101011100; // vC= -164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000111; // iC= -633 
vC = 14'b1111111101010001; // vC= -175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010001; // iC= -623 
vC = 14'b1111111110001001; // vC= -119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000111; // iC= -569 
vC = 14'b1111111100111001; // vC= -199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110100; // iC= -588 
vC = 14'b1111111110110111; // vC=  -73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101011; // iC= -661 
vC = 14'b1111111101101100; // vC= -148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001101; // iC= -627 
vC = 14'b1111111100011000; // vC= -232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001111; // iC= -625 
vC = 14'b1111111101111011; // vC= -133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111111110110001; // vC=  -79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111111; // iC= -577 
vC = 14'b1111111101101101; // vC= -147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001011; // iC= -629 
vC = 14'b1111111100011100; // vC= -228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110111; // iC= -649 
vC = 14'b1111111101001000; // vC= -184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001011; // iC= -565 
vC = 14'b1111111100101001; // vC= -215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110010; // iC= -526 
vC = 14'b1111111110001110; // vC= -114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b1111111101100010; // vC= -158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010000; // iC= -624 
vC = 14'b1111111101101011; // vC= -149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000101; // iC= -635 
vC = 14'b1111111110000110; // vC= -122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000110; // iC= -506 
vC = 14'b1111111101100010; // vC= -158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001000; // iC= -504 
vC = 14'b1111111100101011; // vC= -213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110101; // iC= -587 
vC = 14'b1111111101010101; // vC= -171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110110; // iC= -522 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011001; // iC= -615 
vC = 14'b1111111100111110; // vC= -194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011101; // iC= -547 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000101; // iC= -635 
vC = 14'b1111111100001011; // vC= -245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010000; // iC= -496 
vC = 14'b1111111011111010; // vC= -262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010011; // iC= -557 
vC = 14'b1111111100011101; // vC= -227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110101; // iC= -523 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100110; // iC= -538 
vC = 14'b1111111100000001; // vC= -255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b1111111110000011; // vC= -125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111111011101000; // vC= -280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111011; // iC= -581 
vC = 14'b1111111100100110; // vC= -218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100101; // iC= -539 
vC = 14'b1111111100100100; // vC= -220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010100; // iC= -492 
vC = 14'b1111111101011100; // vC= -164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101101; // iC= -467 
vC = 14'b1111111100110101; // vC= -203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111001; // iC= -583 
vC = 14'b1111111100011000; // vC= -232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110000; // iC= -528 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110001; // iC= -463 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111001; // iC= -455 
vC = 14'b1111111011111100; // vC= -260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110100; // iC= -524 
vC = 14'b1111111100011101; // vC= -227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001011; // iC= -437 
vC = 14'b1111111101010100; // vC= -172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000011; // iC= -573 
vC = 14'b1111111100100101; // vC= -219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010001; // iC= -495 
vC = 14'b1111111101001011; // vC= -181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011001; // iC= -487 
vC = 14'b1111111011101000; // vC= -280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011010; // iC= -486 
vC = 14'b1111111101100001; // vC= -159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110100; // iC= -524 
vC = 14'b1111111100111111; // vC= -193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001110; // iC= -498 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110001; // iC= -463 
vC = 14'b1111111100001000; // vC= -248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001100; // iC= -500 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000111; // iC= -441 
vC = 14'b1111111101011010; // vC= -166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010000; // iC= -496 
vC = 14'b1111111011111110; // vC= -258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100101; // iC= -411 
vC = 14'b1111111011011101; // vC= -291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010000; // iC= -432 
vC = 14'b1111111011111101; // vC= -259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111001; // iC= -519 
vC = 14'b1111111100000100; // vC= -252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001111; // iC= -497 
vC = 14'b1111111101001111; // vC= -177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111001; // iC= -391 
vC = 14'b1111111100110101; // vC= -203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111101; // iC= -515 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100010; // iC= -478 
vC = 14'b1111111100011110; // vC= -226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101010; // iC= -406 
vC = 14'b1111111100000010; // vC= -254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001000; // iC= -440 
vC = 14'b1111111101001001; // vC= -183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111001; // iC= -455 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100010; // iC= -478 
vC = 14'b1111111011001010; // vC= -310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101101; // iC= -467 
vC = 14'b1111111011100001; // vC= -287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011010; // iC= -422 
vC = 14'b1111111100111101; // vC= -195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110100; // iC= -396 
vC = 14'b1111111101000001; // vC= -191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000100; // iC= -508 
vC = 14'b1111111100011110; // vC= -226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101001; // iC= -471 
vC = 14'b1111111010101111; // vC= -337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100110; // iC= -474 
vC = 14'b1111111100100111; // vC= -217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011100; // iC= -420 
vC = 14'b1111111100110001; // vC= -207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000101; // iC= -443 
vC = 14'b1111111011100111; // vC= -281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000010; // iC= -382 
vC = 14'b1111111100110101; // vC= -203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000000; // iC= -384 
vC = 14'b1111111011101100; // vC= -276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001001; // iC= -375 
vC = 14'b1111111100000000; // vC= -256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101001; // iC= -471 
vC = 14'b1111111100110100; // vC= -204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000010; // iC= -446 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101101; // iC= -339 
vC = 14'b1111111100000101; // vC= -251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101110; // iC= -402 
vC = 14'b1111111100011011; // vC= -229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011110; // iC= -354 
vC = 14'b1111111011101111; // vC= -273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100011; // iC= -349 
vC = 14'b1111111010001110; // vC= -370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110110; // iC= -394 
vC = 14'b1111111011100001; // vC= -287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001010; // iC= -374 
vC = 14'b1111111010100100; // vC= -348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100001; // iC= -415 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000111; // iC= -377 
vC = 14'b1111111010110110; // vC= -330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010100; // iC= -364 
vC = 14'b1111111100001101; // vC= -243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011010; // iC= -422 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110011; // iC= -333 
vC = 14'b1111111010010111; // vC= -361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101100; // iC= -404 
vC = 14'b1111111011001000; // vC= -312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011110; // iC= -290 
vC = 14'b1111111011101011; // vC= -277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100000; // iC= -352 
vC = 14'b1111111010100110; // vC= -346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001100; // iC= -308 
vC = 14'b1111111011111011; // vC= -261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000011; // iC= -317 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111110; // iC= -258 
vC = 14'b1111111011111110; // vC= -258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110101; // iC= -267 
vC = 14'b1111111010111101; // vC= -323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000010; // iC= -382 
vC = 14'b1111111100000011; // vC= -253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100111; // iC= -281 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101000; // iC= -344 
vC = 14'b1111111010101111; // vC= -337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010001; // iC= -303 
vC = 14'b1111111011110110; // vC= -266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011011; // iC= -357 
vC = 14'b1111111001110010; // vC= -398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010101; // iC= -363 
vC = 14'b1111111011001110; // vC= -306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010111; // iC= -361 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000101; // iC= -379 
vC = 14'b1111111010011101; // vC= -355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100000; // iC= -352 
vC = 14'b1111111001110010; // vC= -398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011101; // iC= -227 
vC = 14'b1111111010110111; // vC= -329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110111; // iC= -265 
vC = 14'b1111111010111101; // vC= -323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110111; // iC= -265 
vC = 14'b1111111010001111; // vC= -369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110011; // iC= -333 
vC = 14'b1111111011110001; // vC= -271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010100; // iC= -236 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010001; // iC= -239 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101000; // iC= -280 
vC = 14'b1111111001110101; // vC= -395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100101; // iC= -283 
vC = 14'b1111111011101001; // vC= -279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010111; // iC= -233 
vC = 14'b1111111010110000; // vC= -336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110011; // iC= -205 
vC = 14'b1111111011101011; // vC= -277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000010; // iC= -190 
vC = 14'b1111111011101100; // vC= -276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010110; // iC= -298 
vC = 14'b1111111011010110; // vC= -298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010100; // iC= -236 
vC = 14'b1111111010111100; // vC= -324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111110; // iC= -258 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000001; // iC= -319 
vC = 14'b1111111011010011; // vC= -301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111110; // iC= -194 
vC = 14'b1111111010000100; // vC= -380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001101; // iC= -243 
vC = 14'b1111111010011101; // vC= -355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111100; // iC= -260 
vC = 14'b1111111001100000; // vC= -416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100100; // iC= -220 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010000; // iC= -176 
vC = 14'b1111111010001101; // vC= -371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000001; // iC= -255 
vC = 14'b1111111001011001; // vC= -423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100110; // iC= -154 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011000; // iC= -232 
vC = 14'b1111111011011001; // vC= -295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010010; // iC= -174 
vC = 14'b1111111011000111; // vC= -313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011100; // iC= -164 
vC = 14'b1111111010101111; // vC= -337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100100; // iC= -156 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111111; // iC= -129 
vC = 14'b1111111010000001; // vC= -383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011011; // iC= -229 
vC = 14'b1111111010000111; // vC= -377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001100; // iC= -244 
vC = 14'b1111111011001100; // vC= -308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001011; // iC= -181 
vC = 14'b1111111001110010; // vC= -398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010100; // iC= -172 
vC = 14'b1111111010001111; // vC= -369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000101; // iC= -187 
vC = 14'b1111111001101001; // vC= -407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011100; // iC= -228 
vC = 14'b1111111010010111; // vC= -361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011011; // iC= -229 
vC = 14'b1111111010101111; // vC= -337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111001; // iC= -263 
vC = 14'b1111111011001110; // vC= -306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011000; // iC= -232 
vC = 14'b1111111001010100; // vC= -428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000001; // iC= -127 
vC = 14'b1111111010101101; // vC= -339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010100; // iC= -172 
vC = 14'b1111111011001101; // vC= -307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001111; // iC= -177 
vC = 14'b1111111010101001; // vC= -343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010110; // iC= -106 
vC = 14'b1111111001100001; // vC= -415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010011; // iC= -109 
vC = 14'b1111111011100010; // vC= -286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111101; // iC= -131 
vC = 14'b1111111011010101; // vC= -299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001110; // iC= -114 
vC = 14'b1111111010011101; // vC= -355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101011; // iC=  -85 
vC = 14'b1111111010010110; // vC= -362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010000; // iC= -176 
vC = 14'b1111111010001100; // vC= -372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110001; // iC=  -79 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110011; // iC= -141 
vC = 14'b1111111010010011; // vC= -365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111011; // iC= -133 
vC = 14'b1111111001011010; // vC= -422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011011; // iC= -165 
vC = 14'b1111111000111011; // vC= -453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010100; // iC= -108 
vC = 14'b1111111011000010; // vC= -318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001010; // iC=  -54 
vC = 14'b1111111010001010; // vC= -374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001001; // iC=  -55 
vC = 14'b1111111010001111; // vC= -369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101010; // iC=  -86 
vC = 14'b1111111010111011; // vC= -325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011100; // iC=  -36 
vC = 14'b1111111001110111; // vC= -393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000101; // iC= -123 
vC = 14'b1111111010010000; // vC= -368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001011; // iC=  -53 
vC = 14'b1111111011010110; // vC= -298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010101; // iC=   21 
vC = 14'b1111111001100011; // vC= -413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001011; // iC= -117 
vC = 14'b1111111001010101; // vC= -427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101111; // iC=  -17 
vC = 14'b1111111010000110; // vC= -378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011010; // iC=   26 
vC = 14'b1111111001100010; // vC= -414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011111; // iC=   31 
vC = 14'b1111111010010100; // vC= -364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000110; // iC=    6 
vC = 14'b1111111001001110; // vC= -434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110110; // iC=  -10 
vC = 14'b1111111010000100; // vC= -380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010110; // iC=  -42 
vC = 14'b1111111001111101; // vC= -387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011110; // iC=   94 
vC = 14'b1111111000111111; // vC= -449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010000; // iC=   16 
vC = 14'b1111111000110101; // vC= -459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111100; // iC=  124 
vC = 14'b1111111001010110; // vC= -426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111000; // iC=   56 
vC = 14'b1111111010000110; // vC= -378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110100; // iC=   52 
vC = 14'b1111111010010111; // vC= -361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100101; // iC=   37 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001001; // iC=  137 
vC = 14'b1111111010011000; // vC= -360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100101; // iC=   37 
vC = 14'b1111111010110001; // vC= -335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111010; // iC=   58 
vC = 14'b1111111011000110; // vC= -314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011011; // iC=   91 
vC = 14'b1111111010100100; // vC= -348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000110; // iC=  198 
vC = 14'b1111111011001110; // vC= -306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101011; // iC=  171 
vC = 14'b1111111010101111; // vC= -337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001110; // iC=  270 
vC = 14'b1111111010111011; // vC= -325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010000; // iC=  272 
vC = 14'b1111111001110111; // vC= -393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011111; // iC=  223 
vC = 14'b1111111010011100; // vC= -356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111010; // iC=  314 
vC = 14'b1111111010011010; // vC= -358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001110; // iC=  206 
vC = 14'b1111111010101000; // vC= -344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101010; // iC=  234 
vC = 14'b1111111000111110; // vC= -450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011010; // iC=  282 
vC = 14'b1111111010011010; // vC= -358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010101; // iC=  277 
vC = 14'b1111111010010000; // vC= -368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000000; // iC=  256 
vC = 14'b1111111010101010; // vC= -342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111001; // iC=  313 
vC = 14'b1111111011001110; // vC= -306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001101; // iC=  333 
vC = 14'b1111111010010100; // vC= -364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110011; // iC=  435 
vC = 14'b1111111001010001; // vC= -431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101111; // iC=  431 
vC = 14'b1111111001010000; // vC= -432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001100; // iC=  396 
vC = 14'b1111111011011000; // vC= -296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011101; // iC=  477 
vC = 14'b1111111001100001; // vC= -415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011111; // iC=  479 
vC = 14'b1111111001001110; // vC= -434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110001; // iC=  497 
vC = 14'b1111111011000001; // vC= -319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100110; // iC=  422 
vC = 14'b1111111010111111; // vC= -321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000100; // iC=  452 
vC = 14'b1111111011101101; // vC= -275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111000; // iC=  568 
vC = 14'b1111111010111010; // vC= -326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010111; // iC=  599 
vC = 14'b1111111011100000; // vC= -288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101110; // iC=  622 
vC = 14'b1111111010101100; // vC= -340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001111; // iC=  527 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101101; // iC=  557 
vC = 14'b1111111001111011; // vC= -389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111011; // iC=  699 
vC = 14'b1111111010101001; // vC= -343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010000; // iC=  592 
vC = 14'b1111111001100000; // vC= -416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100110; // iC=  614 
vC = 14'b1111111011111001; // vC= -263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101111; // iC=  751 
vC = 14'b1111111011010110; // vC= -298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010100; // iC=  724 
vC = 14'b1111111011111111; // vC= -257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010010; // iC=  658 
vC = 14'b1111111010101001; // vC= -343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101001; // iC=  745 
vC = 14'b1111111010110111; // vC= -329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000011; // iC=  771 
vC = 14'b1111111011111011; // vC= -261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111100; // iC=  828 
vC = 14'b1111111011101001; // vC= -279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001010; // iC=  778 
vC = 14'b1111111100000000; // vC= -256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100101; // iC=  741 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101100; // iC=  748 
vC = 14'b1111111011110101; // vC= -267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001001; // iC=  905 
vC = 14'b1111111011111111; // vC= -257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100110; // iC=  870 
vC = 14'b1111111001111110; // vC= -386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110011; // iC=  819 
vC = 14'b1111111011010010; // vC= -302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101100; // iC=  876 
vC = 14'b1111111010100000; // vC= -352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000110; // iC=  838 
vC = 14'b1111111100011010; // vC= -230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011000; // iC=  856 
vC = 14'b1111111011000001; // vC= -319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100111; // iC=  871 
vC = 14'b1111111010010100; // vC= -364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100010; // iC=  866 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111010; // iC=  954 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010011; // iC=  979 
vC = 14'b1111111010011010; // vC= -358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010010; // iC= 1042 
vC = 14'b1111111010101000; // vC= -344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110100; // iC= 1012 
vC = 14'b1111111100101111; // vC= -209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100111; // iC=  999 
vC = 14'b1111111010110011; // vC= -333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001011; // iC= 1099 
vC = 14'b1111111011101011; // vC= -277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110011; // iC= 1075 
vC = 14'b1111111010110111; // vC= -329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111100; // iC= 1020 
vC = 14'b1111111100110000; // vC= -208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110101; // iC= 1013 
vC = 14'b1111111011010100; // vC= -300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011111; // iC=  991 
vC = 14'b1111111011110000; // vC= -272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111101; // iC= 1149 
vC = 14'b1111111011101001; // vC= -279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001100; // iC= 1100 
vC = 14'b1111111101000001; // vC= -191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000111; // iC= 1159 
vC = 14'b1111111100011101; // vC= -227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110011; // iC= 1075 
vC = 14'b1111111011010111; // vC= -297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001100; // iC= 1164 
vC = 14'b1111111100001010; // vC= -246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011000; // iC= 1112 
vC = 14'b1111111100011000; // vC= -232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101000; // iC= 1128 
vC = 14'b1111111100001101; // vC= -243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011011; // iC= 1115 
vC = 14'b1111111100110001; // vC= -207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110000; // iC= 1136 
vC = 14'b1111111101001000; // vC= -184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101100; // iC= 1132 
vC = 14'b1111111100010101; // vC= -235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000100; // iC= 1220 
vC = 14'b1111111100100011; // vC= -221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101011; // iC= 1195 
vC = 14'b1111111011011100; // vC= -292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001110; // iC= 1230 
vC = 14'b1111111101101001; // vC= -151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011100; // iC= 1180 
vC = 14'b1111111101011111; // vC= -161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b1111111100110110; // vC= -202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010001; // iC= 1297 
vC = 14'b1111111100101111; // vC= -209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011001; // iC= 1177 
vC = 14'b1111111100110111; // vC= -201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b1111111100000010; // vC= -254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010111; // iC= 1303 
vC = 14'b1111111101111011; // vC= -133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010011; // iC= 1235 
vC = 14'b1111111100100111; // vC= -217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101101; // iC= 1197 
vC = 14'b1111111101001000; // vC= -184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001100; // iC= 1356 
vC = 14'b1111111100010110; // vC= -234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101100; // iC= 1260 
vC = 14'b1111111100011100; // vC= -228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111011; // iC= 1275 
vC = 14'b1111111110001001; // vC= -119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010001; // iC= 1361 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010110; // iC= 1238 
vC = 14'b1111111100111101; // vC= -195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100110; // iC= 1382 
vC = 14'b1111111110000000; // vC= -128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111110; // iC= 1342 
vC = 14'b1111111110101110; // vC=  -82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110011; // iC= 1267 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011001; // iC= 1369 
vC = 14'b1111111110010100; // vC= -108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111011; // iC= 1403 
vC = 14'b1111111110011001; // vC= -103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110001; // iC= 1329 
vC = 14'b1111111110110001; // vC=  -79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001001; // iC= 1417 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111011; // iC= 1403 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101000; // iC= 1384 
vC = 14'b1111111110011010; // vC= -102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010001; // iC= 1361 
vC = 14'b1111111101101000; // vC= -152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000110; // iC= 1350 
vC = 14'b1111111101110010; // vC= -142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010101; // iC= 1365 
vC = 14'b1111111110000011; // vC= -125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011011; // iC= 1307 
vC = 14'b1111111101111101; // vC= -131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110010; // iC= 1394 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101011; // iC= 1387 
vC = 14'b1111111110100011; // vC=  -93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011111; // iC= 1311 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100101; // iC= 1445 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010011; // iC= 1363 
vC = 14'b1111111110100011; // vC=  -93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101110; // iC= 1326 
vC = 14'b1111111111111011; // vC=   -5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110100; // iC= 1396 
vC = 14'b1111111111110010; // vC=  -14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000100; // iC= 1348 
vC = 14'b1111111101111000; // vC= -136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101001; // iC= 1449 
vC = 14'b1111111110101100; // vC=  -84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100010; // iC= 1314 
vC = 14'b1111111111000011; // vC=  -61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110010; // iC= 1394 
vC = 14'b1111111110110001; // vC=  -79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101000; // iC= 1320 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100001; // iC= 1441 
vC = 14'b1111111110101100; // vC=  -84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100001; // iC= 1313 
vC = 14'b1111111110101010; // vC=  -86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000101; // iC= 1349 
vC = 14'b0000000000000101; // vC=    5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000110; // iC= 1286 
vC = 14'b0000000000001001; // vC=    9 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011000; // iC= 1368 
vC = 14'b0000000000011101; // vC=   29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010010; // iC= 1298 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011110; // iC= 1438 
vC = 14'b0000000001000101; // vC=   69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100010; // iC= 1378 
vC = 14'b1111111110101100; // vC=  -84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100010; // iC= 1378 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010110; // iC= 1302 
vC = 14'b0000000001000111; // vC=   71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010000; // iC= 1424 
vC = 14'b1111111111000111; // vC=  -57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001010; // iC= 1290 
vC = 14'b1111111111111100; // vC=   -4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010101; // iC= 1301 
vC = 14'b0000000001000001; // vC=   65 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000010; // iC= 1346 
vC = 14'b1111111111100110; // vC=  -26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110110; // iC= 1334 
vC = 14'b0000000000111110; // vC=   62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011011; // iC= 1307 
vC = 14'b0000000001010011; // vC=   83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110000; // iC= 1328 
vC = 14'b1111111111100000; // vC=  -32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000000000000111; // vC=    7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100101; // iC= 1317 
vC = 14'b0000000000101001; // vC=   41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000010; // iC= 1282 
vC = 14'b0000000000110111; // vC=   55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011100; // iC= 1308 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101011; // iC= 1259 
vC = 14'b0000000000110100; // vC=   52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110101; // iC= 1269 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000110; // iC= 1286 
vC = 14'b0000000001100111; // vC=  103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101000; // iC= 1384 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001000; // iC= 1288 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000001; // iC= 1345 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001101; // iC= 1357 
vC = 14'b0000000000001011; // vC=   11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010000; // iC= 1296 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100011; // iC= 1315 
vC = 14'b0000000001101000; // vC=  104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001110; // iC= 1230 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111111; // iC= 1279 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101100; // iC= 1324 
vC = 14'b0000000000111011; // vC=   59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001110; // iC= 1230 
vC = 14'b0000000010000001; // vC=  129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011110; // iC= 1374 
vC = 14'b0000000010100010; // vC=  162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001010; // iC= 1290 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001001; // iC= 1289 
vC = 14'b0000000001111101; // vC=  125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111101; // iC= 1277 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101100; // iC= 1324 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111100; // iC= 1212 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000001; // iC= 1281 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000110; // iC= 1350 
vC = 14'b0000000011000011; // vC=  195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110100; // iC= 1332 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001110; // iC= 1294 
vC = 14'b0000000010000100; // vC=  132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000000; // iC= 1280 
vC = 14'b0000000001011101; // vC=   93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101001; // iC= 1193 
vC = 14'b0000000011100010; // vC=  226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011101; // iC= 1245 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110101; // iC= 1333 
vC = 14'b0000000010000101; // vC=  133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110111; // iC= 1207 
vC = 14'b0000000001101101; // vC=  109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001110; // iC= 1294 
vC = 14'b0000000001101011; // vC=  107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100100; // iC= 1252 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001010; // iC= 1290 
vC = 14'b0000000011011001; // vC=  217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110001; // iC= 1201 
vC = 14'b0000000011011100; // vC=  220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011101; // iC= 1309 
vC = 14'b0000000010000100; // vC=  132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110100; // iC= 1268 
vC = 14'b0000000100000110; // vC=  262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101010; // iC= 1258 
vC = 14'b0000000100100001; // vC=  289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000010; // iC= 1218 
vC = 14'b0000000011111100; // vC=  252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000000; // iC= 1152 
vC = 14'b0000000100001101; // vC=  269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001101; // iC= 1229 
vC = 14'b0000000010100111; // vC=  167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010001; // iC= 1233 
vC = 14'b0000000100011001; // vC=  281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111111; // iC= 1279 
vC = 14'b0000000011011101; // vC=  221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100101; // iC= 1189 
vC = 14'b0000000011110101; // vC=  245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110101; // iC= 1269 
vC = 14'b0000000100111011; // vC=  315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101110; // iC= 1134 
vC = 14'b0000000100101010; // vC=  298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100001; // iC= 1249 
vC = 14'b0000000011000110; // vC=  198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101110; // iC= 1198 
vC = 14'b0000000010110110; // vC=  182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001111; // iC= 1167 
vC = 14'b0000000010111001; // vC=  185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011110; // iC= 1118 
vC = 14'b0000000100000001; // vC=  257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001010; // iC= 1226 
vC = 14'b0000000100001110; // vC=  270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011011; // iC= 1179 
vC = 14'b0000000100110111; // vC=  311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011010; // iC= 1114 
vC = 14'b0000000101001100; // vC=  332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111110; // iC= 1150 
vC = 14'b0000000011001100; // vC=  204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000101; // iC= 1157 
vC = 14'b0000000100111000; // vC=  312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011101; // iC= 1245 
vC = 14'b0000000100110101; // vC=  309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010100; // iC= 1108 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001001; // iC= 1161 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101010; // iC= 1130 
vC = 14'b0000000100010100; // vC=  276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011000; // iC= 1112 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110010; // iC= 1074 
vC = 14'b0000000011110001; // vC=  241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110111; // iC= 1143 
vC = 14'b0000000101011011; // vC=  347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110000; // iC= 1072 
vC = 14'b0000000101011011; // vC=  347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101001; // iC= 1065 
vC = 14'b0000000101111101; // vC=  381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000000100010010; // vC=  274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100010; // iC= 1058 
vC = 14'b0000000100101001; // vC=  297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010001; // iC= 1169 
vC = 14'b0000000101100110; // vC=  358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000011; // iC= 1155 
vC = 14'b0000000100100100; // vC=  292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001100; // iC= 1100 
vC = 14'b0000000101110100; // vC=  372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101101; // iC= 1069 
vC = 14'b0000000110001110; // vC=  398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111111; // iC= 1087 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101011; // iC= 1195 
vC = 14'b0000000100100011; // vC=  291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011000; // iC= 1048 
vC = 14'b0000000110001000; // vC=  392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110000; // iC= 1136 
vC = 14'b0000000101111010; // vC=  378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101011; // iC= 1131 
vC = 14'b0000000110001001; // vC=  393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000010; // iC= 1026 
vC = 14'b0000000100010110; // vC=  278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011011; // iC= 1179 
vC = 14'b0000000100011100; // vC=  284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011111; // iC= 1055 
vC = 14'b0000000100100110; // vC=  294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110111; // iC= 1079 
vC = 14'b0000000110100001; // vC=  417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100100; // iC= 1124 
vC = 14'b0000000101000111; // vC=  327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110101; // iC= 1013 
vC = 14'b0000000101001000; // vC=  328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010010; // iC= 1106 
vC = 14'b0000000110110100; // vC=  436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100010; // iC= 1122 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100001; // iC=  993 
vC = 14'b0000000100110101; // vC=  309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111110; // iC= 1086 
vC = 14'b0000000110000000; // vC=  384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001111; // iC= 1039 
vC = 14'b0000000101100001; // vC=  353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001011; // iC= 1035 
vC = 14'b0000000110010000; // vC=  400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000001; // iC= 1089 
vC = 14'b0000000111011101; // vC=  477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101111; // iC= 1071 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110111; // iC= 1015 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101100; // iC= 1004 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100010; // iC=  994 
vC = 14'b0000000110101001; // vC=  425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011101; // iC= 1117 
vC = 14'b0000000111101100; // vC=  492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111100; // iC= 1084 
vC = 14'b0000000101010000; // vC=  336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100100; // iC=  996 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000101; // iC= 1029 
vC = 14'b0000000101110110; // vC=  374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110111; // iC=  951 
vC = 14'b0000000101100111; // vC=  359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000111; // iC= 1095 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001101; // iC= 1101 
vC = 14'b0000000111100001; // vC=  481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000100; // iC= 1092 
vC = 14'b0000001000000001; // vC=  513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100011; // iC=  931 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100011; // iC= 1059 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001001; // iC= 1033 
vC = 14'b0000000110000010; // vC=  386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000110; // iC= 1030 
vC = 14'b0000000110111010; // vC=  442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111000; // iC= 1080 
vC = 14'b0000000111001100; // vC=  460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110010; // iC= 1010 
vC = 14'b0000000110011001; // vC=  409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010110; // iC= 1046 
vC = 14'b0000001000000011; // vC=  515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000110; // iC=  966 
vC = 14'b0000000111011000; // vC=  472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001010; // iC=  906 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000101; // iC= 1029 
vC = 14'b0000000111111001; // vC=  505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001110; // iC=  974 
vC = 14'b0000000111101000; // vC=  488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011101; // iC=  989 
vC = 14'b0000000110101101; // vC=  429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010111; // iC=  919 
vC = 14'b0000000111111101; // vC=  509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110001; // iC= 1009 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100000; // iC=  928 
vC = 14'b0000000111001101; // vC=  461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100001; // iC=  993 
vC = 14'b0000000111110001; // vC=  497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101100; // iC=  940 
vC = 14'b0000000111100000; // vC=  480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000111; // iC=  967 
vC = 14'b0000000111101011; // vC=  491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011001; // iC=  985 
vC = 14'b0000000110100001; // vC=  417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100001; // iC=  993 
vC = 14'b0000000110111001; // vC=  441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011011; // iC=  859 
vC = 14'b0000000110101100; // vC=  428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010101; // iC=  917 
vC = 14'b0000001000011111; // vC=  543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111110; // iC=  894 
vC = 14'b0000001000111010; // vC=  570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110000; // iC=  944 
vC = 14'b0000001000010111; // vC=  535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010000; // iC=  976 
vC = 14'b0000001000100011; // vC=  547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101101; // iC=  877 
vC = 14'b0000000111101001; // vC=  489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011001; // iC=  857 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110101; // iC=  885 
vC = 14'b0000000111010001; // vC=  465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011101; // iC=  925 
vC = 14'b0000001000100000; // vC=  544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011011; // iC=  859 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101000; // iC=  936 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100100; // iC=  868 
vC = 14'b0000001000111011; // vC=  571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001111; // iC=  847 
vC = 14'b0000001000100111; // vC=  551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111100; // iC=  828 
vC = 14'b0000001001010011; // vC=  595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000100; // iC=  964 
vC = 14'b0000001000010100; // vC=  532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100010; // iC=  930 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010101; // iC=  917 
vC = 14'b0000001000100001; // vC=  545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001110; // iC=  846 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101001; // iC=  809 
vC = 14'b0000001001001000; // vC=  584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110001; // iC=  817 
vC = 14'b0000001001000000; // vC=  576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110000; // iC=  816 
vC = 14'b0000001001110000; // vC=  624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000000; // iC=  896 
vC = 14'b0000001000101011; // vC=  555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011010; // iC=  922 
vC = 14'b0000001000011101; // vC=  541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101111; // iC=  815 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110100; // iC=  884 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000001; // iC=  769 
vC = 14'b0000001001001100; // vC=  588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010010; // iC=  786 
vC = 14'b0000000111110111; // vC=  503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101110; // iC=  814 
vC = 14'b0000001000000001; // vC=  513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100101; // iC=  869 
vC = 14'b0000001000110111; // vC=  567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011000; // iC=  856 
vC = 14'b0000001001110010; // vC=  626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010001; // iC=  785 
vC = 14'b0000001000100011; // vC=  547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001101; // iC=  845 
vC = 14'b0000001010000000; // vC=  640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110000; // iC=  752 
vC = 14'b0000001000001101; // vC=  525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010000; // iC=  848 
vC = 14'b0000001000000001; // vC=  513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100111; // iC=  743 
vC = 14'b0000001001011101; // vC=  605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001001; // iC=  841 
vC = 14'b0000001000010000; // vC=  528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100111; // iC=  807 
vC = 14'b0000001010000110; // vC=  646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010010; // iC=  722 
vC = 14'b0000001010011010; // vC=  666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000110; // iC=  838 
vC = 14'b0000001001001111; // vC=  591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010110; // iC=  726 
vC = 14'b0000001001101010; // vC=  618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001011; // iC=  843 
vC = 14'b0000001010100010; // vC=  674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010110; // iC=  726 
vC = 14'b0000001000011100; // vC=  540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101010; // iC=  810 
vC = 14'b0000001010010011; // vC=  659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111110; // iC=  766 
vC = 14'b0000001000011011; // vC=  539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100101; // iC=  741 
vC = 14'b0000001001001101; // vC=  589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010111; // iC=  727 
vC = 14'b0000001010111001; // vC=  697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110000; // iC=  688 
vC = 14'b0000001001111100; // vC=  636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111111; // iC=  703 
vC = 14'b0000001010011110; // vC=  670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101100; // iC=  748 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101010; // iC=  810 
vC = 14'b0000001000101011; // vC=  555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011110; // iC=  670 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100011; // iC=  803 
vC = 14'b0000001000100111; // vC=  551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101000; // iC=  680 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111001; // iC=  761 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010000; // iC=  720 
vC = 14'b0000001011010000; // vC=  720 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001101; // iC=  653 
vC = 14'b0000001010011000; // vC=  664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010000; // iC=  720 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011010; // iC=  794 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101001; // iC=  745 
vC = 14'b0000001010111111; // vC=  703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110111; // iC=  759 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101100; // iC=  684 
vC = 14'b0000001011011010; // vC=  730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111001; // iC=  761 
vC = 14'b0000001000111111; // vC=  575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111101; // iC=  765 
vC = 14'b0000001011000110; // vC=  710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000111; // iC=  647 
vC = 14'b0000001001111001; // vC=  633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001110; // iC=  718 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101001; // iC=  681 
vC = 14'b0000001001011011; // vC=  603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000011; // iC=  707 
vC = 14'b0000001001111110; // vC=  638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100000; // iC=  736 
vC = 14'b0000001010110000; // vC=  688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001110; // iC=  654 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b0000001010111101; // vC=  701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011101; // iC=  605 
vC = 14'b0000001011100111; // vC=  743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010011; // iC=  595 
vC = 14'b0000001010010011; // vC=  659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001010; // iC=  714 
vC = 14'b0000001010010000; // vC=  656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100000; // iC=  608 
vC = 14'b0000001001110010; // vC=  626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100101; // iC=  677 
vC = 14'b0000001011100100; // vC=  740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011010; // iC=  666 
vC = 14'b0000001011001101; // vC=  717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001001; // iC=  585 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100000; // iC=  608 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000001; // iC=  641 
vC = 14'b0000001011100001; // vC=  737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000101; // iC=  581 
vC = 14'b0000001010101011; // vC=  683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011110; // iC=  606 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110100; // iC=  564 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011011; // iC=  539 
vC = 14'b0000001010111101; // vC=  701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011111; // iC=  607 
vC = 14'b0000001011001010; // vC=  714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011001; // iC=  537 
vC = 14'b0000001001101011; // vC=  619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101001; // iC=  553 
vC = 14'b0000001010001010; // vC=  650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001000; // iC=  520 
vC = 14'b0000001001110011; // vC=  627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011001; // iC=  601 
vC = 14'b0000001011010100; // vC=  724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000011; // iC=  579 
vC = 14'b0000001100001100; // vC=  780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111110; // iC=  574 
vC = 14'b0000001010110010; // vC=  690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000110; // iC=  582 
vC = 14'b0000001100001111; // vC=  783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110001; // iC=  625 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000010; // iC=  578 
vC = 14'b0000001011001011; // vC=  715 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110100; // iC=  564 
vC = 14'b0000001001111101; // vC=  637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000000; // iC=  576 
vC = 14'b0000001011111011; // vC=  763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011010; // iC=  538 
vC = 14'b0000001100001111; // vC=  783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100000; // iC=  544 
vC = 14'b0000001010101111; // vC=  687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111111; // iC=  511 
vC = 14'b0000001011111110; // vC=  766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001101; // iC=  525 
vC = 14'b0000001010010011; // vC=  659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001001; // iC=  585 
vC = 14'b0000001011101000; // vC=  744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100011; // iC=  547 
vC = 14'b0000001010110010; // vC=  690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011110; // iC=  606 
vC = 14'b0000001010001111; // vC=  655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011101; // iC=  541 
vC = 14'b0000001010101101; // vC=  685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110000; // iC=  496 
vC = 14'b0000001100010111; // vC=  791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000101; // iC=  517 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101100; // iC=  556 
vC = 14'b0000001010101110; // vC=  686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100011; // iC=  547 
vC = 14'b0000001010110101; // vC=  693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001101; // iC=  525 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011100; // iC=  476 
vC = 14'b0000001011110101; // vC=  757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001011; // iC=  459 
vC = 14'b0000001010010101; // vC=  661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010110; // iC=  470 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100110; // iC=  486 
vC = 14'b0000001011000001; // vC=  705 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000100; // iC=  516 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010000; // iC=  400 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010001; // iC=  465 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011101; // iC=  413 
vC = 14'b0000001010010110; // vC=  662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111110; // iC=  446 
vC = 14'b0000001100010000; // vC=  784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011111; // iC=  415 
vC = 14'b0000001100001010; // vC=  778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011001; // iC=  409 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111101; // iC=  381 
vC = 14'b0000001011010100; // vC=  724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001100; // iC=  524 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111011; // iC=  443 
vC = 14'b0000001011010100; // vC=  724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101000; // iC=  424 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000100; // iC=  516 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101100; // iC=  364 
vC = 14'b0000001011011110; // vC=  734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101001; // iC=  361 
vC = 14'b0000001011110011; // vC=  755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100101; // iC=  421 
vC = 14'b0000001100010101; // vC=  789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100110; // iC=  358 
vC = 14'b0000001010101110; // vC=  686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101010; // iC=  362 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100111; // iC=  423 
vC = 14'b0000001010110001; // vC=  689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100001; // iC=  353 
vC = 14'b0000001100011101; // vC=  797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101100; // iC=  364 
vC = 14'b0000001100110001; // vC=  817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001000; // iC=  328 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000111; // iC=  327 
vC = 14'b0000001011100100; // vC=  740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010010; // iC=  402 
vC = 14'b0000001100101000; // vC=  808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000001; // iC=  385 
vC = 14'b0000001100100010; // vC=  802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101010; // iC=  426 
vC = 14'b0000001011111111; // vC=  767 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111010; // iC=  442 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111001; // iC=  377 
vC = 14'b0000001010111110; // vC=  702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011101; // iC=  349 
vC = 14'b0000001100011110; // vC=  798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100111; // iC=  295 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110000; // iC=  368 
vC = 14'b0000001010111110; // vC=  702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110011; // iC=  371 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011101; // iC=  413 
vC = 14'b0000001010110101; // vC=  693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110101; // iC=  309 
vC = 14'b0000001101001000; // vC=  840 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011010; // iC=  346 
vC = 14'b0000001100011110; // vC=  798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100101; // iC=  357 
vC = 14'b0000001100000010; // vC=  770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100110; // iC=  358 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011010; // iC=  282 
vC = 14'b0000001011011010; // vC=  730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011110; // iC=  350 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111000; // iC=  376 
vC = 14'b0000001011010100; // vC=  724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011001; // iC=  345 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111101; // iC=  381 
vC = 14'b0000001100100101; // vC=  805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111100; // iC=  380 
vC = 14'b0000001011100100; // vC=  740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101001; // iC=  297 
vC = 14'b0000001100111000; // vC=  824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100100; // iC=  228 
vC = 14'b0000001011100111; // vC=  743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100110; // iC=  358 
vC = 14'b0000001100101100; // vC=  812 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101001; // iC=  361 
vC = 14'b0000001101010010; // vC=  850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001001; // iC=  329 
vC = 14'b0000001101001110; // vC=  846 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000010; // iC=  322 
vC = 14'b0000001011101001; // vC=  745 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000110; // iC=  326 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000111; // iC=  263 
vC = 14'b0000001101010111; // vC=  855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101000; // iC=  296 
vC = 14'b0000001011001100; // vC=  716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111111; // iC=  191 
vC = 14'b0000001011010100; // vC=  724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111111; // iC=  191 
vC = 14'b0000001100100111; // vC=  807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010111; // iC=  279 
vC = 14'b0000001011011001; // vC=  729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011010; // iC=  282 
vC = 14'b0000001011011101; // vC=  733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111100; // iC=  316 
vC = 14'b0000001100000100; // vC=  772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011010; // iC=  218 
vC = 14'b0000001100001000; // vC=  776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010110; // iC=  278 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000101; // iC=  261 
vC = 14'b0000001011011111; // vC=  735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101000; // iC=  168 
vC = 14'b0000001011101010; // vC=  746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100001; // iC=  225 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011001; // iC=  281 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001110; // iC=  142 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101000; // iC=  232 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011011; // iC=  283 
vC = 14'b0000001101000101; // vC=  837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010001; // iC=  145 
vC = 14'b0000001100010000; // vC=  784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010110; // iC=  150 
vC = 14'b0000001100110010; // vC=  818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001111; // iC=  143 
vC = 14'b0000001101101001; // vC=  873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101100; // iC=  108 
vC = 14'b0000001100001011; // vC=  779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011011; // iC=  219 
vC = 14'b0000001100111011; // vC=  827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100111; // iC=  167 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010000; // iC=  144 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010101; // iC=  149 
vC = 14'b0000001100110010; // vC=  818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000101; // iC=   69 
vC = 14'b0000001100000101; // vC=  773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111100; // iC=  124 
vC = 14'b0000001101000011; // vC=  835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101000; // iC=  104 
vC = 14'b0000001101001111; // vC=  847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011100; // iC=   28 
vC = 14'b0000001100010111; // vC=  791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011011; // iC=   27 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101001; // iC=  -23 
vC = 14'b0000001100001010; // vC=  778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101110; // iC=  -18 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000011; // iC=   67 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100010; // iC=  -30 
vC = 14'b0000001101101000; // vC=  872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110101; // iC=  -11 
vC = 14'b0000001101100100; // vC=  868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101000; // iC=  -88 
vC = 14'b0000001100110110; // vC=  822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010111; // iC=  -41 
vC = 14'b0000001100001110; // vC=  782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000010; // iC= -126 
vC = 14'b0000001011100011; // vC=  739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110100; // iC=  -76 
vC = 14'b0000001101001001; // vC=  841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010100; // iC= -108 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110111; // iC= -137 
vC = 14'b0000001100111100; // vC=  828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110011; // iC= -205 
vC = 14'b0000001101011000; // vC=  856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011110; // iC= -162 
vC = 14'b0000001100100010; // vC=  802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011000; // iC= -168 
vC = 14'b0000001100001101; // vC=  781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001000; // iC= -184 
vC = 14'b0000001011010110; // vC=  726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001100; // iC= -180 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101011; // iC= -213 
vC = 14'b0000001100010001; // vC=  785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110110; // iC= -266 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101001; // iC= -215 
vC = 14'b0000001011110011; // vC=  755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111011; // iC= -261 
vC = 14'b0000001100110000; // vC=  816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100101; // iC= -283 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111101; // iC= -387 
vC = 14'b0000001010111100; // vC=  700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110101; // iC= -331 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101110; // iC= -466 
vC = 14'b0000001100101010; // vC=  810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010100; // iC= -428 
vC = 14'b0000001100000110; // vC=  774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101010; // iC= -470 
vC = 14'b0000001100101100; // vC=  812 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001000; // iC= -504 
vC = 14'b0000001101000001; // vC=  833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101001; // iC= -535 
vC = 14'b0000001010110111; // vC=  695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101110; // iC= -466 
vC = 14'b0000001011000110; // vC=  710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011001; // iC= -487 
vC = 14'b0000001100001111; // vC=  783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111001; // iC= -519 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011111; // iC= -481 
vC = 14'b0000001011000101; // vC=  709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111000; // iC= -520 
vC = 14'b0000001100000100; // vC=  772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101011; // iC= -661 
vC = 14'b0000001100110000; // vC=  816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101011; // iC= -597 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001010; // iC= -630 
vC = 14'b0000001011011100; // vC=  732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011011; // iC= -677 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010011; // iC= -749 
vC = 14'b0000001011010101; // vC=  725 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100010; // iC= -670 
vC = 14'b0000001010100011; // vC=  675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100010; // iC= -670 
vC = 14'b0000001011001101; // vC=  717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000000; // iC= -768 
vC = 14'b0000001100100010; // vC=  802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110010; // iC= -718 
vC = 14'b0000001011000000; // vC=  704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001100; // iC= -756 
vC = 14'b0000001100001011; // vC=  779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100000; // iC= -736 
vC = 14'b0000001010101100; // vC=  684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010101; // iC= -875 
vC = 14'b0000001011100110; // vC=  742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011110; // iC= -802 
vC = 14'b0000001011100000; // vC=  736 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010001; // iC= -943 
vC = 14'b0000001010111100; // vC=  700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001110; // iC= -818 
vC = 14'b0000001011110000; // vC=  752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101000; // iC= -856 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010101; // iC= -939 
vC = 14'b0000001011011110; // vC=  734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011111; // iC= -929 
vC = 14'b0000001011000011; // vC=  707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110111; // iC= -969 
vC = 14'b0000001001111101; // vC=  637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b0000001001110011; // vC=  627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100101; // iC= -987 
vC = 14'b0000001011100001; // vC=  737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110111; // iC= -969 
vC = 14'b0000001011100010; // vC=  738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101010; // iC=-1046 
vC = 14'b0000001001010011; // vC=  595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010101; // iC=-1003 
vC = 14'b0000001010000100; // vC=  644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011101; // iC= -995 
vC = 14'b0000001001001000; // vC=  584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111011; // iC=-1157 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100110; // iC=-1178 
vC = 14'b0000001001111111; // vC=  639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010100; // iC=-1068 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101001; // iC=-1111 
vC = 14'b0000001001110011; // vC=  627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010011; // iC=-1133 
vC = 14'b0000001011010000; // vC=  720 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000100; // iC=-1148 
vC = 14'b0000001000111011; // vC=  571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101000; // iC=-1240 
vC = 14'b0000001000110010; // vC=  562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001000; // iC=-1272 
vC = 14'b0000001001100000; // vC=  608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b0000001010001100; // vC=  652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010111; // iC=-1193 
vC = 14'b0000001001010101; // vC=  597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100001; // iC=-1311 
vC = 14'b0000001001100100; // vC=  612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101011; // iC=-1301 
vC = 14'b0000001010011010; // vC=  666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110100; // iC=-1292 
vC = 14'b0000001001100100; // vC=  612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110000; // iC=-1232 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100100; // iC=-1244 
vC = 14'b0000001001000100; // vC=  580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101111; // iC=-1297 
vC = 14'b0000001010001010; // vC=  650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b0000001010000100; // vC=  644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000010; // iC=-1278 
vC = 14'b0000001000011010; // vC=  538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b0000000111110000; // vC=  496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010000; // iC=-1328 
vC = 14'b0000001001101010; // vC=  618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010000; // iC=-1328 
vC = 14'b0000001000110100; // vC=  564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010000; // iC=-1328 
vC = 14'b0000001001011000; // vC=  600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000010; // iC=-1470 
vC = 14'b0000000111111101; // vC=  509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001111; // iC=-1393 
vC = 14'b0000001000000101; // vC=  517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b0000000111001001; // vC=  457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000011; // iC=-1405 
vC = 14'b0000000111110110; // vC=  502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011111; // iC=-1377 
vC = 14'b0000001000011110; // vC=  542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b0000000111000100; // vC=  452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000001001001100; // vC=  588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000000111011011; // vC=  475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011110; // iC=-1442 
vC = 14'b0000001000011101; // vC=  541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101011; // iC=-1493 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b0000001000111111; // vC=  575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010000; // iC=-1456 
vC = 14'b0000000110110000; // vC=  432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b0000001000000001; // vC=  513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000011; // iC=-1533 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111101; // iC=-1475 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000001; // iC=-1599 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011101; // iC=-1507 
vC = 14'b0000001000000101; // vC=  517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010100; // iC=-1516 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000000110001101; // vC=  397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000000110010011; // vC=  403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b0000000111101110; // vC=  494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b0000000111011001; // vC=  473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b0000000101111011; // vC=  379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b0000000110100111; // vC=  423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b0000000101010111; // vC=  343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b0000000101111110; // vC=  382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000000101110100; // vC=  372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b0000000110101000; // vC=  424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b0000000111000011; // vC=  451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b0000000110011001; // vC=  409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b0000000110001010; // vC=  394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b0000000110101000; // vC=  424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b0000000100000101; // vC=  261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b0000000100001110; // vC=  270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b0000000011111011; // vC=  251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b0000000101000101; // vC=  325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b0000000100011010; // vC=  282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010011; // iC=-1581 
vC = 14'b0000000100010000; // vC=  272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b0000000011101001; // vC=  233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b0000000101000110; // vC=  326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b0000000011100110; // vC=  230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000101; // iC=-1595 
vC = 14'b0000000011010011; // vC=  211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b0000000011110010; // vC=  242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011111; // iC=-1633 
vC = 14'b0000000101010110; // vC=  342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b0000000101010010; // vC=  338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000101; // iC=-1595 
vC = 14'b0000000100101001; // vC=  297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b0000000100000101; // vC=  261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b0000000100100100; // vC=  292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b0000000011000011; // vC=  195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b0000000100010010; // vC=  274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101010; // iC=-1686 
vC = 14'b0000000010111110; // vC=  190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b0000000010011000; // vC=  152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b0000000010000011; // vC=  131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b0000000100000100; // vC=  260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110100; // iC=-1612 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100100; // iC=-1564 
vC = 14'b0000000011111010; // vC=  250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b0000000001110010; // vC=  114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110110; // iC=-1674 
vC = 14'b0000000001101001; // vC=  105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b0000000011001111; // vC=  207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000000010001110; // vC=  142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001100; // iC=-1588 
vC = 14'b0000000011000110; // vC=  198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010011; // iC=-1581 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101011; // iC=-1557 
vC = 14'b0000000011001100; // vC=  204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b0000000011001011; // vC=  203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b0000000000100101; // vC=   37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011111; // iC=-1633 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001010; // iC=-1654 
vC = 14'b0000000010100010; // vC=  162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001100; // iC=-1588 
vC = 14'b0000000000001111; // vC=   15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b0000000000001111; // vC=   15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b0000000001011011; // vC=   91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110111; // iC=-1609 
vC = 14'b0000000010001110; // vC=  142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010010; // iC=-1518 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b1111111111111101; // vC=   -3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100011; // iC=-1629 
vC = 14'b1111111111010011; // vC=  -45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100010; // iC=-1502 
vC = 14'b0000000000100101; // vC=   37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111111; // iC=-1473 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100011; // iC=-1501 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100100; // iC=-1628 
vC = 14'b1111111111101101; // vC=  -19 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b0000000001001110; // vC=   78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000000000011011; // vC=   27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101101; // iC=-1491 
vC = 14'b1111111111111001; // vC=   -7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100100; // iC=-1500 
vC = 14'b0000000000100000; // vC=   32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b1111111110101110; // vC=  -82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b1111111110111011; // vC=  -69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b1111111111110001; // vC=  -15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100100; // iC=-1564 
vC = 14'b1111111110010010; // vC= -110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010011; // iC=-1581 
vC = 14'b1111111111011011; // vC=  -37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100101; // iC=-1435 
vC = 14'b1111111110111001; // vC=  -71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b1111111111101100; // vC=  -20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b1111111110101101; // vC=  -83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110011; // iC=-1421 
vC = 14'b1111111110001101; // vC= -115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010011; // iC=-1453 
vC = 14'b1111111110011011; // vC= -101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b1111111110101100; // vC=  -84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b1111111110110011; // vC=  -77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b1111111101011110; // vC= -162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b1111111111100101; // vC=  -27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b1111111111000100; // vC=  -60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110001; // iC=-1551 
vC = 14'b1111111110000001; // vC= -127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111111; // iC=-1409 
vC = 14'b1111111101000010; // vC= -190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b1111111110000000; // vC= -128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111100; // iC=-1476 
vC = 14'b1111111110011100; // vC= -100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010111; // iC=-1449 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101101; // iC=-1491 
vC = 14'b1111111110001101; // vC= -115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110010; // iC=-1486 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b1111111110010100; // vC= -108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011001; // iC=-1447 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b1111111100011110; // vC= -226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100110; // iC=-1370 
vC = 14'b1111111101010010; // vC= -174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110100; // iC=-1356 
vC = 14'b1111111101000011; // vC= -189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111001; // iC=-1415 
vC = 14'b1111111101010010; // vC= -174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b1111111100111010; // vC= -198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110100; // iC=-1420 
vC = 14'b1111111101000101; // vC= -187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b1111111100101100; // vC= -212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b1111111100101011; // vC= -213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010010; // iC=-1390 
vC = 14'b1111111011101001; // vC= -279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b1111111100101011; // vC= -213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010010; // iC=-1454 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010101; // iC=-1323 
vC = 14'b1111111100101000; // vC= -216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010100; // iC=-1388 
vC = 14'b1111111011110100; // vC= -268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010010; // iC=-1390 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010111; // iC=-1321 
vC = 14'b1111111101000000; // vC= -192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110001; // iC=-1359 
vC = 14'b1111111100001100; // vC= -244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000111; // iC=-1337 
vC = 14'b1111111100100111; // vC= -217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100111; // iC=-1369 
vC = 14'b1111111011100011; // vC= -285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b1111111100001010; // vC= -246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001101; // iC=-1331 
vC = 14'b1111111010111001; // vC= -327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010010; // iC=-1326 
vC = 14'b1111111100001000; // vC= -248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b1111111011001111; // vC= -305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b1111111011010001; // vC= -303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101101; // iC=-1363 
vC = 14'b1111111011011100; // vC= -292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001011; // iC=-1397 
vC = 14'b1111111011011001; // vC= -295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111110; // iC=-1282 
vC = 14'b1111111100000100; // vC= -252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b1111111011101010; // vC= -278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110111; // iC=-1289 
vC = 14'b1111111010101010; // vC= -342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000001; // iC=-1279 
vC = 14'b1111111010001001; // vC= -375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111010; // iC=-1350 
vC = 14'b1111111010101000; // vC= -344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111111001110000; // vC= -400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011100; // iC=-1316 
vC = 14'b1111111010001110; // vC= -370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001001; // iC=-1271 
vC = 14'b1111111011101111; // vC= -273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011000; // iC=-1384 
vC = 14'b1111111010101101; // vC= -339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111111011110111; // vC= -265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100001; // iC=-1247 
vC = 14'b1111111010111110; // vC= -322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011001; // iC=-1255 
vC = 14'b1111111001011001; // vC= -423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100101; // iC=-1307 
vC = 14'b1111111010000001; // vC= -383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b1111111001011100; // vC= -420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100111; // iC=-1305 
vC = 14'b1111111010101010; // vC= -342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010001; // iC=-1327 
vC = 14'b1111111011000001; // vC= -319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010111; // iC=-1193 
vC = 14'b1111111001010100; // vC= -428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001011; // iC=-1205 
vC = 14'b1111111010101000; // vC= -344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101110; // iC=-1234 
vC = 14'b1111111010110000; // vC= -336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111111001010000; // vC= -432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011010; // iC=-1318 
vC = 14'b1111111010000010; // vC= -382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011100; // iC=-1252 
vC = 14'b1111111001100010; // vC= -414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101101; // iC=-1171 
vC = 14'b1111111010101111; // vC= -337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011000; // iC=-1192 
vC = 14'b1111111001010110; // vC= -426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011010; // iC=-1254 
vC = 14'b1111111001000010; // vC= -446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100111; // iC=-1241 
vC = 14'b1111111000101001; // vC= -471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000000; // iC=-1216 
vC = 14'b1111111001101001; // vC= -407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111011; // iC=-1221 
vC = 14'b1111111010100011; // vC= -349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111110; // iC=-1154 
vC = 14'b1111111000110110; // vC= -458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001011; // iC=-1269 
vC = 14'b1111111001000110; // vC= -442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001010; // iC=-1270 
vC = 14'b1111111001000111; // vC= -441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b1111111000101111; // vC= -465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001000; // iC=-1144 
vC = 14'b1111111010010011; // vC= -365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b1111111001010010; // vC= -430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b1111111001001010; // vC= -438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010100; // iC=-1132 
vC = 14'b1111110111111001; // vC= -519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011100; // iC=-1188 
vC = 14'b1111111010000011; // vC= -381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100001; // iC=-1183 
vC = 14'b1111111000010010; // vC= -494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101011; // iC=-1173 
vC = 14'b1111111000010100; // vC= -492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001110; // iC=-1202 
vC = 14'b1111111000010101; // vC= -491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000000; // iC=-1216 
vC = 14'b1111110111100010; // vC= -542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011011; // iC=-1189 
vC = 14'b1111111001100001; // vC= -415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001101; // iC=-1139 
vC = 14'b1111111000001111; // vC= -497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001010; // iC=-1078 
vC = 14'b1111111001010000; // vC= -432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111001; // iC=-1223 
vC = 14'b1111111000001000; // vC= -504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001110; // iC=-1074 
vC = 14'b1111111001011001; // vC= -423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011111; // iC=-1057 
vC = 14'b1111111000001000; // vC= -504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100000; // iC=-1120 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011000; // iC=-1064 
vC = 14'b1111110111101010; // vC= -534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001011; // iC=-1141 
vC = 14'b1111110111101011; // vC= -533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110110; // iC=-1162 
vC = 14'b1111110110111111; // vC= -577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000101; // iC=-1083 
vC = 14'b1111110111111110; // vC= -514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001101; // iC=-1139 
vC = 14'b1111111000101011; // vC= -469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001111; // iC=-1073 
vC = 14'b1111110110110101; // vC= -587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110001; // iC=-1103 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100101; // iC=-1051 
vC = 14'b1111110110111000; // vC= -584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011010; // iC=-1062 
vC = 14'b1111110110010101; // vC= -619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000100; // iC=-1148 
vC = 14'b1111110111101010; // vC= -534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101001; // iC=-1111 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111101; // iC=-1091 
vC = 14'b1111110110001010; // vC= -630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011011; // iC=-1125 
vC = 14'b1111110111011100; // vC= -548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111101; // iC=-1027 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110111; // iC=-1033 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001111; // iC=-1009 
vC = 14'b1111110110101111; // vC= -593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b1111110111001101; // vC= -563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111010; // iC=-1030 
vC = 14'b1111110110111010; // vC= -582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000011; // iC=-1021 
vC = 14'b1111110111100000; // vC= -544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100000; // iC=-1056 
vC = 14'b1111110111000110; // vC= -570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011011; // iC= -997 
vC = 14'b1111110111110101; // vC= -523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010101; // iC=-1067 
vC = 14'b1111110111110010; // vC= -526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010011; // iC=-1005 
vC = 14'b1111110101101010; // vC= -662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000010; // iC=-1022 
vC = 14'b1111110111001000; // vC= -568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101010; // iC=-1046 
vC = 14'b1111110110010000; // vC= -624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001001; // iC= -951 
vC = 14'b1111110110010110; // vC= -618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001010; // iC= -950 
vC = 14'b1111110110101001; // vC= -599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001011; // iC= -949 
vC = 14'b1111110111001111; // vC= -561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011000; // iC= -936 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101011; // iC=-1045 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011111; // iC=-1057 
vC = 14'b1111110101110000; // vC= -656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110011; // iC=-1037 
vC = 14'b1111110101011011; // vC= -677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101101; // iC= -979 
vC = 14'b1111110101111000; // vC= -648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000000; // iC= -960 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101110; // iC= -978 
vC = 14'b1111110110011011; // vC= -613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b1111110100101101; // vC= -723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100100; // iC= -924 
vC = 14'b1111110101010000; // vC= -688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101110; // iC= -978 
vC = 14'b1111110101001011; // vC= -693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001010; // iC= -886 
vC = 14'b1111110100111111; // vC= -705 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100011; // iC= -861 
vC = 14'b1111110100110100; // vC= -716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011010; // iC= -934 
vC = 14'b1111110110100110; // vC= -602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101101; // iC= -851 
vC = 14'b1111110110100101; // vC= -603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100010; // iC= -862 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100011; // iC= -925 
vC = 14'b1111110110001100; // vC= -628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110100; // iC= -908 
vC = 14'b1111110110001010; // vC= -630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001100; // iC= -948 
vC = 14'b1111110101101100; // vC= -660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111000; // iC= -904 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011110; // iC= -930 
vC = 14'b1111110100010100; // vC= -748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111000; // iC= -968 
vC = 14'b1111110100010001; // vC= -751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011110; // iC= -930 
vC = 14'b1111110101011001; // vC= -679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000011; // iC= -829 
vC = 14'b1111110101100110; // vC= -666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001011; // iC= -885 
vC = 14'b1111110110001101; // vC= -627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011010; // iC= -934 
vC = 14'b1111110011111101; // vC= -771 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100010; // iC= -798 
vC = 14'b1111110100000111; // vC= -761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100001; // iC= -863 
vC = 14'b1111110011110111; // vC= -777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101101; // iC= -851 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011101; // iC= -803 
vC = 14'b1111110100110010; // vC= -718 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001100; // iC= -884 
vC = 14'b1111110100000101; // vC= -763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111001; // iC= -839 
vC = 14'b1111110100111111; // vC= -705 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010111; // iC= -873 
vC = 14'b1111110101001100; // vC= -692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101100; // iC= -852 
vC = 14'b1111110100111100; // vC= -708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110110; // iC= -778 
vC = 14'b1111110101010010; // vC= -686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111110101011000; // vC= -680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011001; // iC= -871 
vC = 14'b1111110100101001; // vC= -727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010100; // iC= -876 
vC = 14'b1111110100001001; // vC= -759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110101; // iC= -843 
vC = 14'b1111110101100011; // vC= -669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101110; // iC= -850 
vC = 14'b1111110100011001; // vC= -743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010100; // iC= -748 
vC = 14'b1111110011011111; // vC= -801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001000; // iC= -760 
vC = 14'b1111110100110010; // vC= -718 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011100; // iC= -868 
vC = 14'b1111110101001111; // vC= -689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010001; // iC= -751 
vC = 14'b1111110100100100; // vC= -732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000110; // iC= -826 
vC = 14'b1111110101010111; // vC= -681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100110; // iC= -730 
vC = 14'b1111110011110000; // vC= -784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001010; // iC= -694 
vC = 14'b1111110101000011; // vC= -701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111100; // iC= -836 
vC = 14'b1111110100101001; // vC= -727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011111; // iC= -737 
vC = 14'b1111110011111101; // vC= -771 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011011; // iC= -677 
vC = 14'b1111110011001101; // vC= -819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011000; // iC= -808 
vC = 14'b1111110100001011; // vC= -757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111110100101110; // vC= -722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100011; // iC= -797 
vC = 14'b1111110011111100; // vC= -772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011001; // iC= -679 
vC = 14'b1111110011010011; // vC= -813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111110010101001; // vC= -855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011111; // iC= -737 
vC = 14'b1111110011110001; // vC= -783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110001; // iC= -719 
vC = 14'b1111110010101100; // vC= -852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000001; // iC= -639 
vC = 14'b1111110011010111; // vC= -809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110101; // iC= -651 
vC = 14'b1111110010111110; // vC= -834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001011; // iC= -693 
vC = 14'b1111110011110001; // vC= -783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001111; // iC= -625 
vC = 14'b1111110100100001; // vC= -735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000010; // iC= -766 
vC = 14'b1111110010101001; // vC= -855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100101; // iC= -731 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011000; // iC= -616 
vC = 14'b1111110010101011; // vC= -853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111101; // iC= -707 
vC = 14'b1111110010110011; // vC= -845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010011; // iC= -621 
vC = 14'b1111110011010011; // vC= -813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100000; // iC= -672 
vC = 14'b1111110001111010; // vC= -902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111000; // iC= -648 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001110; // iC= -690 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100101; // iC= -667 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010101; // iC= -619 
vC = 14'b1111110100001001; // vC= -759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111000; // iC= -712 
vC = 14'b1111110100001111; // vC= -753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000000; // iC= -576 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010101; // iC= -619 
vC = 14'b1111110011100111; // vC= -793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000100; // iC= -572 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110010; // iC= -654 
vC = 14'b1111110001101101; // vC= -915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000100; // iC= -572 
vC = 14'b1111110100000100; // vC= -764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011110; // iC= -610 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000000; // iC= -640 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111000; // iC= -648 
vC = 14'b1111110010100101; // vC= -859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000000; // iC= -640 
vC = 14'b1111110010001011; // vC= -885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010111; // iC= -617 
vC = 14'b1111110001101000; // vC= -920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100011; // iC= -605 
vC = 14'b1111110001011100; // vC= -932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101000; // iC= -600 
vC = 14'b1111110001011111; // vC= -929 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111000; // iC= -648 
vC = 14'b1111110001011001; // vC= -935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000001; // iC= -639 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111011; // iC= -517 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010101; // iC= -555 
vC = 14'b1111110010000111; // vC= -889 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000100; // iC= -508 
vC = 14'b1111110011011101; // vC= -803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000011; // iC= -509 
vC = 14'b1111110010000000; // vC= -896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000100; // iC= -508 
vC = 14'b1111110001111001; // vC= -903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110000; // iC= -592 
vC = 14'b1111110011001101; // vC= -819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001100; // iC= -500 
vC = 14'b1111110011011111; // vC= -801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001010; // iC= -502 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100001; // iC= -479 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000001; // iC= -447 
vC = 14'b1111110001111011; // vC= -901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010000; // iC= -560 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111001; // iC= -455 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010001; // iC= -495 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100110; // iC= -538 
vC = 14'b1111110011001101; // vC= -819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010011; // iC= -493 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101011; // iC= -469 
vC = 14'b1111110011000011; // vC= -829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100001; // iC= -479 
vC = 14'b1111110011001111; // vC= -817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010000; // iC= -432 
vC = 14'b1111110010101011; // vC= -853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001001; // iC= -503 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110101; // iC= -395 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100110; // iC= -410 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111100; // iC= -516 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110011; // iC= -397 
vC = 14'b1111110001001100; // vC= -948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000111; // iC= -377 
vC = 14'b1111110010010001; // vC= -879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010111; // iC= -425 
vC = 14'b1111110000110111; // vC= -969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011000; // iC= -360 
vC = 14'b1111110010100110; // vC= -858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000010; // iC= -446 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110111; // iC= -329 
vC = 14'b1111110010111110; // vC= -834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000110; // iC= -378 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011101; // iC= -419 
vC = 14'b1111110001000110; // vC= -954 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101110; // iC= -466 
vC = 14'b1111110001000000; // vC= -960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000100; // iC= -316 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010101; // iC= -299 
vC = 14'b1111110010100111; // vC= -857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101011; // iC= -405 
vC = 14'b1111110001111010; // vC= -902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001100; // iC= -308 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011011; // iC= -357 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000010; // iC= -382 
vC = 14'b1111110010001100; // vC= -884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110101; // iC= -395 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110001; // iC= -399 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110100; // iC= -268 
vC = 14'b1111110000001100; // vC=-1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101111; // iC= -273 
vC = 14'b1111110000001110; // vC=-1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111001; // iC= -327 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000001; // iC= -319 
vC = 14'b1111110000100001; // vC= -991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010110; // iC= -362 
vC = 14'b1111110000101111; // vC= -977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001101; // iC= -243 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011010; // iC= -358 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011111; // iC= -353 
vC = 14'b1111110000100111; // vC= -985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111011; // iC= -261 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110000; // iC= -336 
vC = 14'b1111110000001111; // vC=-1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011000; // iC= -296 
vC = 14'b1111110000100011; // vC= -989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100111; // iC= -345 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101101; // iC= -211 
vC = 14'b1111110001100011; // vC= -925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101000; // iC= -344 
vC = 14'b1111110000010011; // vC=-1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100000; // iC= -224 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010001; // iC= -239 
vC = 14'b1111110000100000; // vC= -992 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001101; // iC= -179 
vC = 14'b1111110001110101; // vC= -907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101011; // iC= -213 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000101; // iC= -187 
vC = 14'b1111110000111001; // vC= -967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101000; // iC= -280 
vC = 14'b1111110000100111; // vC= -985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110010; // iC= -142 
vC = 14'b1111110000011010; // vC= -998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010000; // iC= -240 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000111; // iC= -249 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010100; // iC= -108 
vC = 14'b1111101111110100; // vC=-1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011001; // iC= -167 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100001; // iC= -159 
vC = 14'b1111110001100100; // vC= -924 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101100; // iC= -148 
vC = 14'b1111110000100101; // vC= -987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001000; // iC= -184 
vC = 14'b1111110000100100; // vC= -988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110111; // iC=  -73 
vC = 14'b1111110000111011; // vC= -965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100000; // iC=  -96 
vC = 14'b1111110000101000; // vC= -984 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111011; // iC= -133 
vC = 14'b1111101111111111; // vC=-1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000101; // iC=    5 
vC = 14'b1111101111110110; // vC=-1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011110; // iC=  -34 
vC = 14'b1111110010000100; // vC= -892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000100; // iC=  -60 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011111; // iC=  -33 
vC = 14'b1111110001111010; // vC= -902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000010; // iC=   66 
vC = 14'b1111110010010001; // vC= -879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010010; // iC=   82 
vC = 14'b1111110000100100; // vC= -988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010111; // iC=   23 
vC = 14'b1111110000111001; // vC= -967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110111; // iC=  119 
vC = 14'b1111110000111100; // vC= -964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111111; // iC=   63 
vC = 14'b1111110000010111; // vC=-1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110000; // iC=  112 
vC = 14'b1111110001011001; // vC= -935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110000; // iC=  112 
vC = 14'b1111110000010011; // vC=-1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110100; // iC=  180 
vC = 14'b1111110010001000; // vC= -888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110011; // iC=  179 
vC = 14'b1111110000110011; // vC= -973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110110; // iC=  182 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110100; // iC=  116 
vC = 14'b1111110000010000; // vC=-1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100111; // iC=  231 
vC = 14'b1111101111111111; // vC=-1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011010; // iC=  154 
vC = 14'b1111110000000111; // vC=-1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000000; // iC=  256 
vC = 14'b1111110010000001; // vC= -895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111110; // iC=  190 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111001; // iC=  313 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011001; // iC=  281 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110101; // iC=  373 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110000; // iC=  432 
vC = 14'b1111110010001011; // vC= -885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010101; // iC=  405 
vC = 14'b1111101111111100; // vC=-1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011010; // iC=  474 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111001; // iC=  505 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111011; // iC=  507 
vC = 14'b1111110010010001; // vC= -879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001111; // iC=  463 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000011; // iC=  515 
vC = 14'b1111110000111100; // vC= -964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111001; // iC=  441 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000011; // iC=  515 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101011; // iC=  491 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011110; // iC=  542 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011111; // iC=  671 
vC = 14'b1111110001001110; // vC= -946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010101; // iC=  597 
vC = 14'b1111110000010111; // vC=-1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110010; // iC=  690 
vC = 14'b1111110000111100; // vC= -964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b1111110000010101; // vC=-1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001010; // iC=  778 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110011; // iC=  755 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100011; // iC=  675 
vC = 14'b1111110000111000; // vC= -968 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101111; // iC=  751 
vC = 14'b1111110010110010; // vC= -846 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001110; // iC=  846 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011111; // iC=  799 
vC = 14'b1111110010110101; // vC= -843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001101; // iC=  781 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011100; // iC=  924 
vC = 14'b1111110000111001; // vC= -967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010100; // iC=  916 
vC = 14'b1111110010101000; // vC= -856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010101; // iC=  917 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101100; // iC=  876 
vC = 14'b1111110010100111; // vC= -857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111110; // iC=  894 
vC = 14'b1111110011001011; // vC= -821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010001; // iC=  977 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011111; // iC=  991 
vC = 14'b1111110001010111; // vC= -937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110101; // iC= 1077 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000000; // iC=  960 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101110; // iC= 1070 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010101; // iC=  981 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111100; // iC= 1084 
vC = 14'b1111110011010010; // vC= -814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110011; // iC= 1075 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101110; // iC= 1070 
vC = 14'b1111110010000100; // vC= -892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b1111110011001000; // vC= -824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000111; // iC= 1223 
vC = 14'b1111110010111100; // vC= -836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101100; // iC= 1132 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000010; // iC= 1154 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111110; // iC= 1150 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111111; // iC= 1215 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010000; // iC= 1168 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000000; // iC= 1344 
vC = 14'b1111110010110101; // vC= -843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011011; // iC= 1243 
vC = 14'b1111110011101000; // vC= -792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010010; // iC= 1362 
vC = 14'b1111110100001111; // vC= -753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010011; // iC= 1235 
vC = 14'b1111110010010101; // vC= -875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110000; // iC= 1328 
vC = 14'b1111110100100011; // vC= -733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000010; // iC= 1346 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110001; // iC= 1329 
vC = 14'b1111110100100100; // vC= -732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010100; // iC= 1428 
vC = 14'b1111110100111001; // vC= -711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010010; // iC= 1362 
vC = 14'b1111110100101101; // vC= -723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000001; // iC= 1409 
vC = 14'b1111110010101100; // vC= -852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011001; // iC= 1433 
vC = 14'b1111110100100100; // vC= -732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000010; // iC= 1410 
vC = 14'b1111110011000111; // vC= -825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101000; // iC= 1384 
vC = 14'b1111110011010011; // vC= -813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111001; // iC= 1529 
vC = 14'b1111110100111101; // vC= -707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100000; // iC= 1440 
vC = 14'b1111110101001111; // vC= -689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110000; // iC= 1456 
vC = 14'b1111110100001011; // vC= -757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100111; // iC= 1511 
vC = 14'b1111110011011100; // vC= -804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110000; // iC= 1456 
vC = 14'b1111110011110001; // vC= -783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010100; // iC= 1492 
vC = 14'b1111110101100101; // vC= -667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001100; // iC= 1484 
vC = 14'b1111110100000000; // vC= -768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000100; // iC= 1540 
vC = 14'b1111110100011111; // vC= -737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111110; // iC= 1534 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001001; // iC= 1609 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010010; // iC= 1554 
vC = 14'b1111110011111110; // vC= -770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101101; // iC= 1645 
vC = 14'b1111110110000100; // vC= -636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110101; // iC= 1653 
vC = 14'b1111110100010100; // vC= -748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100101; // iC= 1573 
vC = 14'b1111110100110100; // vC= -716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010000; // iC= 1616 
vC = 14'b1111110110011000; // vC= -616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b1111110101100001; // vC= -671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111010; // iC= 1594 
vC = 14'b1111110110010101; // vC= -619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b1111110101010101; // vC= -683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b1111110110101110; // vC= -594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b1111110101010010; // vC= -686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111110; // iC= 1726 
vC = 14'b1111110111001011; // vC= -565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b1111110110001010; // vC= -630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111110101100001; // vC= -671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011011; // iC= 1755 
vC = 14'b1111110101100011; // vC= -669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b1111110111011110; // vC= -546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b1111110110101001; // vC= -599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b1111110110000011; // vC= -637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011011; // iC= 1755 
vC = 14'b1111110111001100; // vC= -564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110101; // iC= 1845 
vC = 14'b1111110110100011; // vC= -605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b1111110111100010; // vC= -542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111110111101011; // vC= -533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b1111110110001000; // vC= -632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b1111110110101001; // vC= -599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001000; // iC= 1864 
vC = 14'b1111110110010001; // vC= -623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000100; // iC= 1732 
vC = 14'b1111110111011100; // vC= -548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b1111111000010100; // vC= -492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100100; // iC= 1764 
vC = 14'b1111110111101100; // vC= -532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011001; // iC= 1881 
vC = 14'b1111111000000101; // vC= -507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001010; // iC= 1738 
vC = 14'b1111111000001001; // vC= -503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b1111110111100101; // vC= -539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b1111110110101011; // vC= -597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b1111111000100010; // vC= -478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b1111111001001101; // vC= -435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111011; // iC= 1851 
vC = 14'b1111110111110011; // vC= -525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011011; // iC= 1819 
vC = 14'b1111110111011000; // vC= -552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010010; // iC= 1874 
vC = 14'b1111110111111010; // vC= -518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b1111111000101001; // vC= -471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010011; // iC= 1747 
vC = 14'b1111111001011110; // vC= -418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111111001011001; // vC= -423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b1111110111100110; // vC= -538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b1111110111111011; // vC= -517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b1111111001010110; // vC= -426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b1111111010010001; // vC= -367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b1111111000101010; // vC= -470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110101; // iC= 1781 
vC = 14'b1111111000010111; // vC= -489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010111; // iC= 1751 
vC = 14'b1111111001001110; // vC= -434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000010; // iC= 1858 
vC = 14'b1111111001111110; // vC= -386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011011; // iC= 1755 
vC = 14'b1111111000011101; // vC= -483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001101; // iC= 1869 
vC = 14'b1111111001000001; // vC= -447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b1111111010100110; // vC= -346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b1111111011001011; // vC= -309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b1111111011001111; // vC= -305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b1111111000111101; // vC= -451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111111; // iC= 1791 
vC = 14'b1111111001100110; // vC= -410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110110; // iC= 1846 
vC = 14'b1111111001010110; // vC= -426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000101; // iC= 1797 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b1111111010011110; // vC= -354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b1111111010110110; // vC= -330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b1111111010111100; // vC= -324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b1111111001110011; // vC= -397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b1111111010101000; // vC= -344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b1111111010100010; // vC= -350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b1111111010111000; // vC= -328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b1111111100001110; // vC= -242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111111100000110; // vC= -250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000101; // iC= 1797 
vC = 14'b1111111011001010; // vC= -310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b1111111011101110; // vC= -274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b1111111100100110; // vC= -218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011011; // iC= 1819 
vC = 14'b1111111100001111; // vC= -241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b1111111101010010; // vC= -174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b1111111011001100; // vC= -308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001001; // iC= 1737 
vC = 14'b1111111011000010; // vC= -318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b1111111101010001; // vC= -175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100000; // iC= 1824 
vC = 14'b1111111101010101; // vC= -171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001101; // iC= 1869 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b1111111101001001; // vC= -183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110001; // iC= 1777 
vC = 14'b1111111101010010; // vC= -174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111111101011010; // vC= -166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110101; // iC= 1845 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001100; // iC= 1804 
vC = 14'b1111111100001000; // vC= -248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b1111111110000101; // vC= -123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b1111111110001111; // vC= -113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b1111111101110001; // vC= -143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110000; // iC= 1840 
vC = 14'b1111111110000001; // vC= -127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b1111111100101110; // vC= -210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110100; // iC= 1780 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111100; // iC= 1788 
vC = 14'b1111111110100010; // vC=  -94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b1111111101101001; // vC= -151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000111; // iC= 1799 
vC = 14'b1111111111010111; // vC=  -41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110111; // iC= 1783 
vC = 14'b1111111110111110; // vC=  -66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b1111111111001001; // vC=  -55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010110; // iC= 1686 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b1111111110011011; // vC= -101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b1111111101101110; // vC= -146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b1111111101100011; // vC= -157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000110; // iC= 1734 
vC = 14'b1111111111100110; // vC=  -26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111110; // iC= 1790 
vC = 14'b1111111110011101; // vC=  -99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111111101101101; // vC= -147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b1111111110010010; // vC= -110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b1111111110011110; // vC=  -98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111111111100000; // vC=  -32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000000000010110; // vC=   22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b1111111111010010; // vC=  -46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b1111111111110000; // vC=  -16 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000000000111000; // vC=   56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111101; // iC= 1789 
vC = 14'b0000000000100010; // vC=   34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100110; // iC= 1702 
vC = 14'b1111111111011001; // vC=  -39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b0000000000101001; // vC=   41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100100; // iC= 1764 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b0000000000110000; // vC=   48 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101110; // iC= 1646 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b1111111111010110; // vC=  -42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b0000000001011011; // vC=   91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000000000010101; // vC=   21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000100; // iC= 1668 
vC = 14'b1111111111110001; // vC=  -15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b0000000000100101; // vC=   37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b1111111111110111; // vC=   -9 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011100; // iC= 1628 
vC = 14'b1111111111101010; // vC=  -22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111110; // iC= 1726 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010011; // iC= 1619 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000100; // iC= 1732 
vC = 14'b0000000010000100; // vC=  132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100010; // iC= 1762 
vC = 14'b0000000010000001; // vC=  129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100000; // iC= 1632 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b0000000010011000; // vC=  152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110100; // iC= 1652 
vC = 14'b0000000001011110; // vC=   94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b0000000000011010; // vC=   26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b0000000010101100; // vC=  172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010111; // iC= 1751 
vC = 14'b0000000010111110; // vC=  190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b0000000010100100; // vC=  164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100101; // iC= 1637 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010101; // iC= 1685 
vC = 14'b0000000001011110; // vC=   94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100111; // iC= 1639 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b0000000001101011; // vC=  107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111111; // iC= 1663 
vC = 14'b0000000011101100; // vC=  236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b0000000010011110; // vC=  158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100001; // iC= 1633 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b0000000011110110; // vC=  246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b0000000011010100; // vC=  212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110000; // iC= 1648 
vC = 14'b0000000010100011; // vC=  163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011011; // iC= 1627 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b0000000011000101; // vC=  197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100001; // iC= 1633 
vC = 14'b0000000011110101; // vC=  245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100110; // iC= 1574 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b0000000011010110; // vC=  214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b0000000010110010; // vC=  178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b0000000010111001; // vC=  185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b0000000100000111; // vC=  263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b0000000010111101; // vC=  189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b0000000100101011; // vC=  299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000101; // iC= 1669 
vC = 14'b0000000101001100; // vC=  332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001100; // iC= 1676 
vC = 14'b0000000011011101; // vC=  221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b0000000100100111; // vC=  295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010110; // iC= 1558 
vC = 14'b0000000011100001; // vC=  225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111001; // iC= 1593 
vC = 14'b0000000100000000; // vC=  256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010001; // iC= 1553 
vC = 14'b0000000100001001; // vC=  265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110111; // iC= 1527 
vC = 14'b0000000101011101; // vC=  349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b0000000100000111; // vC=  263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000001; // iC= 1601 
vC = 14'b0000000100000001; // vC=  257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011110; // iC= 1630 
vC = 14'b0000000101011111; // vC=  351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101100; // iC= 1644 
vC = 14'b0000000100001111; // vC=  271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011110; // iC= 1630 
vC = 14'b0000000101010010; // vC=  338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110000; // iC= 1520 
vC = 14'b0000000100100011; // vC=  291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110000; // iC= 1584 
vC = 14'b0000000011110100; // vC=  244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000010; // iC= 1538 
vC = 14'b0000000100001010; // vC=  266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101000; // iC= 1576 
vC = 14'b0000000100010101; // vC=  277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101010; // iC= 1514 
vC = 14'b0000000101100110; // vC=  358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010010; // iC= 1618 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101101; // iC= 1581 
vC = 14'b0000000110100001; // vC=  417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000100; // iC= 1604 
vC = 14'b0000000100111100; // vC=  316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000111; // iC= 1543 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011111; // iC= 1567 
vC = 14'b0000000101011011; // vC=  347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111000; // iC= 1464 
vC = 14'b0000000101001010; // vC=  330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001101; // iC= 1549 
vC = 14'b0000000111000001; // vC=  449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011111; // iC= 1567 
vC = 14'b0000000110001010; // vC=  394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010011; // iC= 1555 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011110; // iC= 1502 
vC = 14'b0000000110011011; // vC=  411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110101; // iC= 1525 
vC = 14'b0000000101000000; // vC=  320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110101; // iC= 1461 
vC = 14'b0000000101111010; // vC=  378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101100; // iC= 1580 
vC = 14'b0000000110011100; // vC=  412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011001; // iC= 1561 
vC = 14'b0000000101101111; // vC=  367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100100; // iC= 1444 
vC = 14'b0000000101111010; // vC=  378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010101; // iC= 1429 
vC = 14'b0000000101100011; // vC=  355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b0000000110101100; // vC=  428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101000; // iC= 1512 
vC = 14'b0000000101100110; // vC=  358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111101; // iC= 1533 
vC = 14'b0000000111100101; // vC=  485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110101; // iC= 1461 
vC = 14'b0000000110101011; // vC=  427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010110; // iC= 1430 
vC = 14'b0000000111110111; // vC=  503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001011; // iC= 1483 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011000; // iC= 1496 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011111; // iC= 1439 
vC = 14'b0000001000001011; // vC=  523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011101; // iC= 1437 
vC = 14'b0000000110110011; // vC=  435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101001; // iC= 1449 
vC = 14'b0000000110001111; // vC=  399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101100; // iC= 1388 
vC = 14'b0000000110101100; // vC=  428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100011; // iC= 1507 
vC = 14'b0000000111100101; // vC=  485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000001; // iC= 1473 
vC = 14'b0000001000010000; // vC=  528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101001; // iC= 1385 
vC = 14'b0000001000010001; // vC=  529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000110; // iC= 1478 
vC = 14'b0000001000000011; // vC=  515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101110; // iC= 1454 
vC = 14'b0000000111111111; // vC=  511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011001; // iC= 1433 
vC = 14'b0000000111101000; // vC=  488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011010; // iC= 1370 
vC = 14'b0000001000001100; // vC=  524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100000; // iC= 1504 
vC = 14'b0000000111001011; // vC=  459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111101; // iC= 1405 
vC = 14'b0000001001010111; // vC=  599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010000; // iC= 1360 
vC = 14'b0000001000111111; // vC=  575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101000; // iC= 1384 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000111; // iC= 1415 
vC = 14'b0000001000001111; // vC=  527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100110; // iC= 1446 
vC = 14'b0000001001001111; // vC=  591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000001; // iC= 1473 
vC = 14'b0000001000001100; // vC=  524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111101; // iC= 1405 
vC = 14'b0000001001100100; // vC=  612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011110; // iC= 1438 
vC = 14'b0000001001111001; // vC=  633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001010; // iC= 1354 
vC = 14'b0000000111110100; // vC=  500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010001; // iC= 1425 
vC = 14'b0000001000001010; // vC=  522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100000; // iC= 1440 
vC = 14'b0000000111101010; // vC=  490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100101; // iC= 1317 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001000; // iC= 1352 
vC = 14'b0000001001111011; // vC=  635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110111; // iC= 1463 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110101; // iC= 1461 
vC = 14'b0000001001011000; // vC=  600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101011; // iC= 1323 
vC = 14'b0000001000100101; // vC=  549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000110; // iC= 1350 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b0000001000001011; // vC=  523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101001; // iC= 1321 
vC = 14'b0000001000001110; // vC=  526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110100; // iC= 1332 
vC = 14'b0000001001111001; // vC=  633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001100; // iC= 1356 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001001; // iC= 1353 
vC = 14'b0000001001000011; // vC=  579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101011; // iC= 1387 
vC = 14'b0000001001000000; // vC=  576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110111; // iC= 1271 
vC = 14'b0000001010111100; // vC=  700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010111; // iC= 1367 
vC = 14'b0000001000110000; // vC=  560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000000; // iC= 1344 
vC = 14'b0000001001000100; // vC=  580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111011; // iC= 1339 
vC = 14'b0000001010011011; // vC=  667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010010; // iC= 1298 
vC = 14'b0000001000111010; // vC=  570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001001; // iC= 1353 
vC = 14'b0000001010111000; // vC=  696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100101; // iC= 1253 
vC = 14'b0000001001010011; // vC=  595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011010; // iC= 1242 
vC = 14'b0000001001011000; // vC=  600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101001; // iC= 1385 
vC = 14'b0000001001111001; // vC=  633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101011; // iC= 1259 
vC = 14'b0000001001100110; // vC=  614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111000; // iC= 1336 
vC = 14'b0000001010000110; // vC=  646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001100; // iC= 1292 
vC = 14'b0000001010001001; // vC=  649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001010; // iC= 1226 
vC = 14'b0000001011110100; // vC=  756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111001; // iC= 1273 
vC = 14'b0000001011011011; // vC=  731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111111; // iC= 1343 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010001; // iC= 1297 
vC = 14'b0000001011101101; // vC=  749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001000; // iC= 1352 
vC = 14'b0000001010001000; // vC=  648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110001; // iC= 1329 
vC = 14'b0000001011011011; // vC=  731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000111; // iC= 1287 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101100; // iC= 1324 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011111; // iC= 1247 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000001010110101; // vC=  693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011010; // iC= 1306 
vC = 14'b0000001100011111; // vC=  799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010000; // iC= 1296 
vC = 14'b0000001011011001; // vC=  729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011101; // iC= 1181 
vC = 14'b0000001010010011; // vC=  659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010101; // iC= 1301 
vC = 14'b0000001100100011; // vC=  803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101100; // iC= 1260 
vC = 14'b0000001100001111; // vC=  783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101110; // iC= 1262 
vC = 14'b0000001010110000; // vC=  688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001111; // iC= 1167 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000000; // iC= 1216 
vC = 14'b0000001011011111; // vC=  735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001100; // iC= 1164 
vC = 14'b0000001100000010; // vC=  770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000001; // iC= 1217 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011001; // iC= 1241 
vC = 14'b0000001011000101; // vC=  709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000001100100101; // vC=  805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001100; // iC= 1228 
vC = 14'b0000001101000000; // vC=  832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010101; // iC= 1173 
vC = 14'b0000001100011010; // vC=  794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111110; // iC= 1150 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010111; // iC= 1175 
vC = 14'b0000001101001001; // vC=  841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101000; // iC= 1256 
vC = 14'b0000001100101111; // vC=  815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011110; // iC= 1246 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111001; // iC= 1209 
vC = 14'b0000001011100011; // vC=  739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010111; // iC= 1239 
vC = 14'b0000001011100110; // vC=  742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001111; // iC= 1231 
vC = 14'b0000001011100001; // vC=  737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000000; // iC= 1216 
vC = 14'b0000001100111111; // vC=  831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100101; // iC= 1189 
vC = 14'b0000001100110101; // vC=  821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100101; // iC= 1125 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000101; // iC= 1221 
vC = 14'b0000001011110011; // vC=  755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101000; // iC= 1128 
vC = 14'b0000001101111100; // vC=  892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000110; // iC= 1158 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001011; // iC= 1163 
vC = 14'b0000001100001011; // vC=  779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101000; // iC= 1128 
vC = 14'b0000001100011000; // vC=  792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111100; // iC= 1212 
vC = 14'b0000001101000111; // vC=  839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b0000001101100110; // vC=  870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101010; // iC= 1130 
vC = 14'b0000001100010001; // vC=  785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110001; // iC= 1137 
vC = 14'b0000001100100101; // vC=  805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100110; // iC= 1062 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000100; // iC= 1156 
vC = 14'b0000001101010101; // vC=  853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011110; // iC= 1182 
vC = 14'b0000001100010000; // vC=  784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111101; // iC= 1085 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010101; // iC= 1173 
vC = 14'b0000001101100101; // vC=  869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100110; // iC= 1062 
vC = 14'b0000001100010110; // vC=  790 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111101; // iC= 1085 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001101; // iC= 1101 
vC = 14'b0000001101000011; // vC=  835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011110; // iC= 1118 
vC = 14'b0000001100111010; // vC=  826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000110; // iC= 1030 
vC = 14'b0000001100101110; // vC=  814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010001; // iC= 1041 
vC = 14'b0000001110010010; // vC=  914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100011; // iC= 1123 
vC = 14'b0000001110001000; // vC=  904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100001; // iC=  993 
vC = 14'b0000001101101011; // vC=  875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111100; // iC= 1084 
vC = 14'b0000001101000111; // vC=  839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000111; // iC= 1031 
vC = 14'b0000001101110111; // vC=  887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011111; // iC= 1119 
vC = 14'b0000001100111110; // vC=  830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100110; // iC= 1126 
vC = 14'b0000001101101001; // vC=  873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100001; // iC= 1057 
vC = 14'b0000001110011001; // vC=  921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011011; // iC=  987 
vC = 14'b0000001110001110; // vC=  910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100001; // iC= 1057 
vC = 14'b0000001101001001; // vC=  841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011110; // iC= 1054 
vC = 14'b0000001101010101; // vC=  853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111010; // iC= 1082 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001100; // iC= 1100 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111000; // iC=  952 
vC = 14'b0000001101111111; // vC=  895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100101; // iC=  933 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110000; // iC= 1072 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110010; // iC= 1074 
vC = 14'b0000001110100011; // vC=  931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001011; // iC= 1035 
vC = 14'b0000001101110111; // vC=  887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101010; // iC= 1002 
vC = 14'b0000001101111100; // vC=  892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010011; // iC= 1043 
vC = 14'b0000001101111001; // vC=  889 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010001; // iC=  913 
vC = 14'b0000001110000101; // vC=  901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100101; // iC=  933 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000001; // iC= 1025 
vC = 14'b0000001101110101; // vC=  885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110101; // iC=  885 
vC = 14'b0000001110000000; // vC=  896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010000; // iC=  976 
vC = 14'b0000001111101101; // vC= 1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111001; // iC= 1017 
vC = 14'b0000001110000111; // vC=  903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111100; // iC=  956 
vC = 14'b0000001110001100; // vC=  908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101101; // iC=  941 
vC = 14'b0000001111101100; // vC= 1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110010; // iC=  882 
vC = 14'b0000001110010110; // vC=  918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001100; // iC=  908 
vC = 14'b0000001110101111; // vC=  943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010010; // iC=  978 
vC = 14'b0000001111010010; // vC=  978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011101; // iC=  861 
vC = 14'b0000001111110101; // vC= 1013 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b0000010000100010; // vC= 1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101011; // iC=  939 
vC = 14'b0000001111000000; // vC=  960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010011; // iC=  851 
vC = 14'b0000001110011011; // vC=  923 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101000; // iC=  936 
vC = 14'b0000010000000110; // vC= 1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001111; // iC=  911 
vC = 14'b0000001111111000; // vC= 1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001011; // iC=  971 
vC = 14'b0000010000101011; // vC= 1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010011; // iC=  851 
vC = 14'b0000010000101010; // vC= 1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010011; // iC=  851 
vC = 14'b0000001111101000; // vC= 1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101111; // iC=  943 
vC = 14'b0000010000010111; // vC= 1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101000; // iC=  808 
vC = 14'b0000001110111011; // vC=  955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001010; // iC=  906 
vC = 14'b0000001111100100; // vC=  996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100000; // iC=  800 
vC = 14'b0000001111001001; // vC=  969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011100; // iC=  860 
vC = 14'b0000010001000101; // vC= 1093 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110011; // iC=  819 
vC = 14'b0000001111111100; // vC= 1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011101; // iC=  925 
vC = 14'b0000010000010110; // vC= 1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100001; // iC=  929 
vC = 14'b0000001111110101; // vC= 1013 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011011; // iC=  923 
vC = 14'b0000001111111001; // vC= 1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011101; // iC=  797 
vC = 14'b0000010000010111; // vC= 1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111100; // iC=  764 
vC = 14'b0000010000011100; // vC= 1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110110; // iC=  758 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100111; // iC=  871 
vC = 14'b0000010001011100; // vC= 1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b0000010000101010; // vC= 1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111001; // iC=  825 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101010; // iC=  810 
vC = 14'b0000010001011001; // vC= 1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001001; // iC=  841 
vC = 14'b0000010001010110; // vC= 1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011000; // iC=  792 
vC = 14'b0000010001100000; // vC= 1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001100; // iC=  780 
vC = 14'b0000001111101100; // vC= 1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110101; // iC=  821 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011110; // iC=  798 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101011; // iC=  811 
vC = 14'b0000010000101000; // vC= 1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011101; // iC=  733 
vC = 14'b0000010000100000; // vC= 1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111101; // iC=  765 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100011; // iC=  739 
vC = 14'b0000010001000000; // vC= 1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000011; // iC=  707 
vC = 14'b0000001111101101; // vC= 1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b0000010000100110; // vC= 1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101010; // iC=  810 
vC = 14'b0000010000110000; // vC= 1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000100; // iC=  772 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110100; // iC=  692 
vC = 14'b0000001111110111; // vC= 1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111100; // iC=  700 
vC = 14'b0000010000110101; // vC= 1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111101; // iC=  765 
vC = 14'b0000010001010100; // vC= 1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001000; // iC=  648 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110011; // iC=  691 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001001; // iC=  713 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000001; // iC=  769 
vC = 14'b0000010000001101; // vC= 1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000001; // iC=  705 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111100; // iC=  636 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101010; // iC=  746 
vC = 14'b0000010010000101; // vC= 1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101101; // iC=  749 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000101; // iC=  645 
vC = 14'b0000010000010101; // vC= 1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100100; // iC=  676 
vC = 14'b0000010000110001; // vC= 1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111101; // iC=  637 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011101; // iC=  733 
vC = 14'b0000001111111111; // vC= 1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100101; // iC=  613 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001100; // iC=  652 
vC = 14'b0000010001110000; // vC= 1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001110; // iC=  590 
vC = 14'b0000010000000100; // vC= 1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011010; // iC=  730 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100110; // iC=  614 
vC = 14'b0000010000001100; // vC= 1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011111; // iC=  607 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001110; // iC=  718 
vC = 14'b0000010000100001; // vC= 1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100100; // iC=  676 
vC = 14'b0000010001111001; // vC= 1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110111; // iC=  695 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011111; // iC=  543 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100000; // iC=  608 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010010; // iC=  594 
vC = 14'b0000010001001110; // vC= 1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011100; // iC=  604 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000111; // iC=  647 
vC = 14'b0000010010010101; // vC= 1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000001; // iC=  577 
vC = 14'b0000010010010111; // vC= 1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010100; // iC=  596 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011001; // iC=  665 
vC = 14'b0000010000100111; // vC= 1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101001; // iC=  617 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100111; // iC=  615 
vC = 14'b0000010010101101; // vC= 1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001000; // iC=  520 
vC = 14'b0000010000101110; // vC= 1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001111; // iC=  591 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011011; // iC=  603 
vC = 14'b0000010001110110; // vC= 1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000101; // iC=  517 
vC = 14'b0000010011000011; // vC= 1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111110; // iC=  574 
vC = 14'b0000010010010101; // vC= 1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100111; // iC=  615 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001101; // iC=  589 
vC = 14'b0000010000110001; // vC= 1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110100; // iC=  500 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010011; // iC=  531 
vC = 14'b0000010001101001; // vC= 1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111110; // iC=  446 
vC = 14'b0000010011001011; // vC= 1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010001; // iC=  529 
vC = 14'b0000010001000000; // vC= 1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010011; // iC=  467 
vC = 14'b0000010001010110; // vC= 1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100000; // iC=  544 
vC = 14'b0000010010001011; // vC= 1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000001; // iC=  513 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001101; // iC=  461 
vC = 14'b0000010001101110; // vC= 1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110101; // iC=  565 
vC = 14'b0000010010011110; // vC= 1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010100; // iC=  468 
vC = 14'b0000010001000001; // vC= 1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000101; // iC=  453 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101100; // iC=  556 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101011; // iC=  491 
vC = 14'b0000010011000110; // vC= 1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001010; // iC=  394 
vC = 14'b0000010010100111; // vC= 1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010110; // iC=  406 
vC = 14'b0000010010001100; // vC= 1164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111010; // iC=  506 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110011; // iC=  435 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011101; // iC=  413 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111010; // iC=  378 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111011; // iC=  443 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110010; // iC=  434 
vC = 14'b0000010010011101; // vC= 1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100111; // iC=  423 
vC = 14'b0000010001100000; // vC= 1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011111; // iC=  415 
vC = 14'b0000010001100011; // vC= 1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111001; // iC=  441 
vC = 14'b0000010001111111; // vC= 1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011011; // iC=  347 
vC = 14'b0000010010110001; // vC= 1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011101; // iC=  477 
vC = 14'b0000010001111101; // vC= 1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111110; // iC=  382 
vC = 14'b0000010011001011; // vC= 1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010111; // iC=  343 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110100; // iC=  436 
vC = 14'b0000010001111111; // vC= 1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100110; // iC=  422 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010011; // iC=  403 
vC = 14'b0000010001110010; // vC= 1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000001; // iC=  321 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001111; // iC=  335 
vC = 14'b0000010011010101; // vC= 1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101000; // iC=  360 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100010; // iC=  290 
vC = 14'b0000010011101111; // vC= 1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100000; // iC=  416 
vC = 14'b0000010011010111; // vC= 1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101001; // iC=  297 
vC = 14'b0000010010101011; // vC= 1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101001; // iC=  361 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010001; // iC=  337 
vC = 14'b0000010011101110; // vC= 1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101111; // iC=  239 
vC = 14'b0000010001011001; // vC= 1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111111; // iC=  319 
vC = 14'b0000010010100100; // vC= 1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110101; // iC=  309 
vC = 14'b0000010010010111; // vC= 1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111111; // iC=  191 
vC = 14'b0000010011000010; // vC= 1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010100; // iC=  276 
vC = 14'b0000010011010000; // vC= 1232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110100; // iC=  244 
vC = 14'b0000010001111100; // vC= 1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110110; // iC=  246 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010110; // iC=  214 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010111; // iC=  279 
vC = 14'b0000010001101111; // vC= 1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000100; // iC=  132 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000110; // iC=  198 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010111; // iC=  151 
vC = 14'b0000010011101100; // vC= 1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101110; // iC=  110 
vC = 14'b0000010010010110; // vC= 1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111001; // iC=  121 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111011; // iC=  123 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001110; // iC=   78 
vC = 14'b0000010001011111; // vC= 1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010110; // iC=   86 
vC = 14'b0000010001101111; // vC= 1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010110; // iC=  150 
vC = 14'b0000010001100011; // vC= 1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001111; // iC=   79 
vC = 14'b0000010010010110; // vC= 1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101100; // iC=   44 
vC = 14'b0000010001101011; // vC= 1131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100101; // iC=  -27 
vC = 14'b0000010010110011; // vC= 1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010010; // iC=   18 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110010; // iC=  -14 
vC = 14'b0000010010001101; // vC= 1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101011; // iC=   43 
vC = 14'b0000010010000010; // vC= 1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011110; // iC=  -34 
vC = 14'b0000010011011000; // vC= 1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011111; // iC=  -97 
vC = 14'b0000010011011010; // vC= 1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111000; // iC=   -8 
vC = 14'b0000010010100011; // vC= 1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101010; // iC= -150 
vC = 14'b0000010011001111; // vC= 1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100010; // iC=  -94 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101011; // iC= -149 
vC = 14'b0000010010010100; // vC= 1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101100; // iC= -212 
vC = 14'b0000010001110111; // vC= 1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010101; // iC= -235 
vC = 14'b0000010001011001; // vC= 1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000111; // iC= -185 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010011; // iC= -173 
vC = 14'b0000010010100001; // vC= 1185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011010; // iC= -230 
vC = 14'b0000010011000001; // vC= 1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011110; // iC= -290 
vC = 14'b0000010010100101; // vC= 1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111100; // iC= -196 
vC = 14'b0000010001111101; // vC= 1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011100; // iC= -228 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000011; // iC= -253 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100011; // iC= -413 
vC = 14'b0000010001101000; // vC= 1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111110; // iC= -386 
vC = 14'b0000010010000011; // vC= 1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111011; // iC= -453 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101101; // iC= -403 
vC = 14'b0000010011000110; // vC= 1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010110; // iC= -426 
vC = 14'b0000010010101110; // vC= 1198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010101; // iC= -427 
vC = 14'b0000010001000000; // vC= 1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100010; // iC= -478 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111001; // iC= -519 
vC = 14'b0000010001100011; // vC= 1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111011; // iC= -581 
vC = 14'b0000010010000001; // vC= 1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000010; // iC= -510 
vC = 14'b0000010010100001; // vC= 1185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101101; // iC= -467 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001001; // iC= -631 
vC = 14'b0000010001000010; // vC= 1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101011; // iC= -661 
vC = 14'b0000010001000001; // vC= 1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111100; // iC= -580 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110010; // iC= -590 
vC = 14'b0000010010111111; // vC= 1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001101; // iC= -691 
vC = 14'b0000010001101110; // vC= 1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111001; // iC= -711 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100000; // iC= -672 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101110; // iC= -722 
vC = 14'b0000010001100101; // vC= 1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001010; // iC= -694 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001010; // iC= -694 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001100; // iC= -756 
vC = 14'b0000010000011100; // vC= 1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100010; // iC= -862 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111111; // iC= -769 
vC = 14'b0000010000111001; // vC= 1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000110; // iC= -890 
vC = 14'b0000010000011101; // vC= 1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110001; // iC= -847 
vC = 14'b0000010000110000; // vC= 1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001101; // iC= -883 
vC = 14'b0000010000000100; // vC= 1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100010; // iC= -798 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001111; // iC= -817 
vC = 14'b0000010000101100; // vC= 1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000111; // iC= -953 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000100; // iC= -892 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111110; // iC= -962 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000010; // iC=-1022 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011000; // iC= -936 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101011; // iC= -981 
vC = 14'b0000010001101001; // vC= 1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000000; // iC= -960 
vC = 14'b0000010001000110; // vC= 1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100001; // iC=-1119 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000010; // iC=-1022 
vC = 14'b0000010000101000; // vC= 1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111001; // iC=-1031 
vC = 14'b0000001111011000; // vC=  984 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101100; // iC=-1044 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101011; // iC=-1109 
vC = 14'b0000001111011111; // vC=  991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000011; // iC=-1149 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000011; // iC=-1213 
vC = 14'b0000001111000011; // vC=  963 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010111; // iC=-1193 
vC = 14'b0000010000100100; // vC= 1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110000; // iC=-1232 
vC = 14'b0000001111110010; // vC= 1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110000; // iC=-1232 
vC = 14'b0000010000000000; // vC= 1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001000; // iC=-1208 
vC = 14'b0000010000111010; // vC= 1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010111; // iC=-1193 
vC = 14'b0000001110100100; // vC=  932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110011; // iC=-1229 
vC = 14'b0000010000010001; // vC= 1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001001; // iC=-1271 
vC = 14'b0000001111011010; // vC=  986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001011; // iC=-1269 
vC = 14'b0000010000000100; // vC= 1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000100; // iC=-1276 
vC = 14'b0000001110010110; // vC=  918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010101; // iC=-1323 
vC = 14'b0000001111111010; // vC= 1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100001; // iC=-1375 
vC = 14'b0000001111010011; // vC=  979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001110; // iC=-1266 
vC = 14'b0000001110111100; // vC=  956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110100; // iC=-1356 
vC = 14'b0000001111001100; // vC=  972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101110; // iC=-1362 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011111; // iC=-1313 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010100; // iC=-1324 
vC = 14'b0000001101100100; // vC=  868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010110; // iC=-1322 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b0000001101110010; // vC=  882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b0000001101001001; // vC=  841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011101; // iC=-1443 
vC = 14'b0000001111001110; // vC=  974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b0000001110010001; // vC=  913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100110; // iC=-1434 
vC = 14'b0000001100111100; // vC=  828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010001; // iC=-1455 
vC = 14'b0000001111000011; // vC=  963 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010001; // iC=-1391 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111101; // iC=-1475 
vC = 14'b0000001100011010; // vC=  794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010101; // iC=-1451 
vC = 14'b0000001100110010; // vC=  818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b0000001101001111; // vC=  847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010111; // iC=-1449 
vC = 14'b0000001101100000; // vC=  864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b0000001101111011; // vC=  891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100100; // iC=-1500 
vC = 14'b0000001110000100; // vC=  900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011110; // iC=-1442 
vC = 14'b0000001110010010; // vC=  914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011000; // iC=-1512 
vC = 14'b0000001011111100; // vC=  764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000111; // iC=-1465 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b0000001101011111; // vC=  863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010111; // iC=-1449 
vC = 14'b0000001011100001; // vC=  737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b0000001011011101; // vC=  733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100100; // iC=-1436 
vC = 14'b0000001100011101; // vC=  797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b0000001011101000; // vC=  744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111110; // iC=-1538 
vC = 14'b0000001011000100; // vC=  708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110001; // iC=-1487 
vC = 14'b0000001011101010; // vC=  746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011011; // iC=-1445 
vC = 14'b0000001101001100; // vC=  844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b0000001101001110; // vC=  846 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b0000001010101010; // vC=  682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b0000001100111010; // vC=  826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000011; // iC=-1469 
vC = 14'b0000001010110011; // vC=  691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b0000001100011010; // vC=  794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010001; // iC=-1455 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100100; // iC=-1564 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010010; // iC=-1518 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b0000001011101011; // vC=  747 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100111; // iC=-1497 
vC = 14'b0000001010110101; // vC=  693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b0000001010001101; // vC=  653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b0000001001111000; // vC=  632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001101; // iC=-1459 
vC = 14'b0000001010010101; // vC=  661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b0000001010100101; // vC=  677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b0000001001100010; // vC=  610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b0000001001010111; // vC=  599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b0000001011010111; // vC=  727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000100; // iC=-1468 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111101; // iC=-1539 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b0000001011000111; // vC=  711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010111; // iC=-1513 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000001001110100; // vC=  628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111010; // iC=-1478 
vC = 14'b0000001000111100; // vC=  572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100111; // iC=-1497 
vC = 14'b0000001001100111; // vC=  615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001111; // iC=-1457 
vC = 14'b0000001000100100; // vC=  548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b0000001001101010; // vC=  618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100100; // iC=-1564 
vC = 14'b0000001001110101; // vC=  629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000001001001111; // vC=  591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111111; // iC=-1537 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b0000001001001000; // vC=  584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000001001001111; // vC=  591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b0000001001101100; // vC=  620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b0000001000110111; // vC=  567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000111; // iC=-1465 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b0000001001001111; // vC=  591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b0000000111011000; // vC=  472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b0000001000011010; // vC=  538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b0000000111101001; // vC=  489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001101; // iC=-1459 
vC = 14'b0000001000110010; // vC=  562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000001000111101; // vC=  573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b0000001000100010; // vC=  546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000000111101110; // vC=  494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b0000000110100010; // vC=  418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b0000000110010011; // vC=  403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b0000000110110101; // vC=  437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100111; // iC=-1497 
vC = 14'b0000001000011101; // vC=  541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110010; // iC=-1486 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b0000000111010100; // vC=  468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b0000000111101111; // vC=  495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010111; // iC=-1513 
vC = 14'b0000000110110100; // vC=  436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b0000000110101101; // vC=  429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b0000000101110011; // vC=  371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b0000000111001011; // vC=  459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111001; // iC=-1479 
vC = 14'b0000000101110000; // vC=  368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011011; // iC=-1445 
vC = 14'b0000000101011000; // vC=  344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111100; // iC=-1540 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100111; // iC=-1497 
vC = 14'b0000000110100011; // vC=  419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b0000000100111101; // vC=  317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b0000000101101101; // vC=  365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b0000000110010100; // vC=  404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111011; // iC=-1541 
vC = 14'b0000000100110000; // vC=  304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000000101100010; // vC=  354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000000101101110; // vC=  366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b0000000101011101; // vC=  349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000110; // iC=-1402 
vC = 14'b0000000101111000; // vC=  376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000000100010100; // vC=  276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b0000000101111110; // vC=  382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b0000000101111101; // vC=  381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b0000000101001110; // vC=  334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000000101001111; // vC=  335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000111; // iC=-1529 
vC = 14'b0000000011111000; // vC=  248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010010; // iC=-1518 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011000; // iC=-1448 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b0000000101010110; // vC=  342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b0000000100001011; // vC=  267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000000100101010; // vC=  298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b0000000100110101; // vC=  309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b0000000011000010; // vC=  194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100100; // iC=-1436 
vC = 14'b0000000011011001; // vC=  217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b0000000100100101; // vC=  293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100101; // iC=-1435 
vC = 14'b0000000100010001; // vC=  273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b0000000100100100; // vC=  292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110001; // iC=-1487 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001110; // iC=-1458 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b0000000100010100; // vC=  276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b0000000010110010; // vC=  178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101010; // iC=-1430 
vC = 14'b0000000011101110; // vC=  238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b0000000010110010; // vC=  178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100100; // iC=-1372 
vC = 14'b0000000011111011; // vC=  251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011111; // iC=-1505 
vC = 14'b0000000011111100; // vC=  252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110011; // iC=-1357 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010110; // iC=-1386 
vC = 14'b0000000011110010; // vC=  242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011011; // iC=-1381 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111001; // iC=-1415 
vC = 14'b0000000100000110; // vC=  262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b0000000010010011; // vC=  147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100110; // iC=-1370 
vC = 14'b0000000011000000; // vC=  192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101011; // iC=-1365 
vC = 14'b0000000010011011; // vC=  155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010000; // iC=-1456 
vC = 14'b0000000011100111; // vC=  231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101110; // iC=-1362 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010001; // iC=-1391 
vC = 14'b0000000010000000; // vC=  128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011111; // iC=-1441 
vC = 14'b0000000011010111; // vC=  215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b0000000001000100; // vC=   68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110010; // iC=-1422 
vC = 14'b0000000010000110; // vC=  134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000011; // iC=-1341 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101100; // iC=-1428 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010011; // iC=-1325 
vC = 14'b0000000001110010; // vC=  114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111100; // iC=-1412 
vC = 14'b0000000001011101; // vC=   93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110011; // iC=-1421 
vC = 14'b0000000000100100; // vC=   36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001110; // iC=-1458 
vC = 14'b0000000001111000; // vC=  120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b0000000000100101; // vC=   37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b0000000000011011; // vC=   27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100111; // iC=-1305 
vC = 14'b0000000000011100; // vC=   28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b0000000000010110; // vC=   22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101101; // iC=-1363 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101101; // iC=-1363 
vC = 14'b0000000001111111; // vC=  127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011100; // iC=-1444 
vC = 14'b0000000000000100; // vC=    4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b1111111111110001; // vC=  -15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110101; // iC=-1419 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100011; // iC=-1309 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110000; // iC=-1360 
vC = 14'b1111111111100011; // vC=  -29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010101; // iC=-1387 
vC = 14'b1111111111111110; // vC=   -2 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011011; // iC=-1381 
vC = 14'b0000000001100000; // vC=   96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101001; // iC=-1367 
vC = 14'b0000000000111111; // vC=   63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110101; // iC=-1419 
vC = 14'b1111111111110001; // vC=  -15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111111111001000; // vC=  -56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110000; // iC=-1360 
vC = 14'b0000000000111110; // vC=   62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b0000000000101110; // vC=   46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b1111111111001001; // vC=  -55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111000; // iC=-1416 
vC = 14'b1111111111011010; // vC=  -38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111111; // iC=-1409 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011000; // iC=-1320 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010001; // iC=-1391 
vC = 14'b1111111111010010; // vC=  -46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001001; // iC=-1399 
vC = 14'b1111111110111111; // vC=  -65 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111000; // iC=-1352 
vC = 14'b0000000000001101; // vC=   13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010010; // iC=-1262 
vC = 14'b1111111111001011; // vC=  -53 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110101; // iC=-1355 
vC = 14'b1111111111110100; // vC=  -12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001010; // iC=-1334 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000000; // iC=-1280 
vC = 14'b1111111110000000; // vC= -128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111100; // iC=-1348 
vC = 14'b1111111110111011; // vC=  -69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111111; // iC=-1281 
vC = 14'b0000000000001101; // vC=   13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100011; // iC=-1373 
vC = 14'b0000000000000111; // vC=    7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010001; // iC=-1327 
vC = 14'b1111111110100110; // vC=  -90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111110; // iC=-1282 
vC = 14'b1111111101111011; // vC= -133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b1111111111100111; // vC=  -25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b1111111110111001; // vC=  -71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110000; // iC=-1360 
vC = 14'b1111111101011000; // vC= -168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110100; // iC=-1292 
vC = 14'b1111111111001100; // vC=  -52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110101; // iC=-1227 
vC = 14'b1111111111100011; // vC=  -29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111010; // iC=-1350 
vC = 14'b1111111101010100; // vC= -172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101010; // iC=-1302 
vC = 14'b1111111110011100; // vC= -100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100111; // iC=-1241 
vC = 14'b1111111110011011; // vC= -101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001000; // iC=-1208 
vC = 14'b1111111110001000; // vC= -120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101100; // iC=-1236 
vC = 14'b1111111110111101; // vC=  -67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111111; // iC=-1281 
vC = 14'b1111111110010000; // vC= -112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000101; // iC=-1211 
vC = 14'b1111111101010111; // vC= -169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000011; // iC=-1341 
vC = 14'b1111111110100001; // vC=  -95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100100; // iC=-1308 
vC = 14'b1111111101111111; // vC= -129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001111; // iC=-1265 
vC = 14'b1111111100101000; // vC= -216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000111; // iC=-1273 
vC = 14'b1111111100101111; // vC= -209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101011; // iC=-1237 
vC = 14'b1111111110101010; // vC=  -86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010111; // iC=-1257 
vC = 14'b1111111110100011; // vC=  -93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001010; // iC=-1270 
vC = 14'b1111111110000011; // vC= -125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000001; // iC=-1215 
vC = 14'b1111111100000110; // vC= -250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111010; // iC=-1286 
vC = 14'b1111111100101111; // vC= -209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b1111111101000110; // vC= -186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110111; // iC=-1289 
vC = 14'b1111111100010101; // vC= -235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b1111111110010010; // vC= -110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000101; // iC=-1211 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000010; // iC=-1278 
vC = 14'b1111111100010100; // vC= -236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110011; // iC=-1229 
vC = 14'b1111111100110111; // vC= -201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100001; // iC=-1247 
vC = 14'b1111111011111110; // vC= -258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000110; // iC=-1210 
vC = 14'b1111111101000101; // vC= -187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001001; // iC=-1271 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110101; // iC=-1163 
vC = 14'b1111111101010010; // vC= -174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101101; // iC=-1235 
vC = 14'b1111111101010101; // vC= -171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001100; // iC=-1140 
vC = 14'b1111111011101101; // vC= -275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101010; // iC=-1174 
vC = 14'b1111111100111011; // vC= -197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000111; // iC=-1209 
vC = 14'b1111111101011011; // vC= -165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100001; // iC=-1183 
vC = 14'b1111111011001000; // vC= -312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001000; // iC=-1272 
vC = 14'b1111111011100100; // vC= -284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110010; // iC=-1230 
vC = 14'b1111111100101000; // vC= -216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111010; // iC=-1222 
vC = 14'b1111111011110010; // vC= -270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111101; // iC=-1155 
vC = 14'b1111111100000000; // vC= -256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000000; // iC=-1216 
vC = 14'b1111111011100001; // vC= -287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101111; // iC=-1169 
vC = 14'b1111111011011001; // vC= -295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b1111111010111100; // vC= -324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100101; // iC=-1115 
vC = 14'b1111111011110101; // vC= -267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110110; // iC=-1226 
vC = 14'b1111111011001100; // vC= -308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011010; // iC=-1126 
vC = 14'b1111111011110011; // vC= -269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001100; // iC=-1204 
vC = 14'b1111111011100111; // vC= -281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100111; // iC=-1177 
vC = 14'b1111111011011100; // vC= -292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100100; // iC=-1116 
vC = 14'b1111111010001000; // vC= -376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101000; // iC=-1176 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110011; // iC=-1229 
vC = 14'b1111111011001111; // vC= -305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001100; // iC=-1076 
vC = 14'b1111111011011100; // vC= -292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011101; // iC=-1059 
vC = 14'b1111111011101100; // vC= -276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100100; // iC=-1180 
vC = 14'b1111111011001011; // vC= -309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100111; // iC=-1113 
vC = 14'b1111111100000010; // vC= -254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011001; // iC=-1191 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100000; // iC=-1120 
vC = 14'b1111111010010000; // vC= -368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101001; // iC=-1111 
vC = 14'b1111111001101011; // vC= -405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001010; // iC=-1142 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001000; // iC=-1080 
vC = 14'b1111111001110100; // vC= -396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011010; // iC=-1126 
vC = 14'b1111111001011100; // vC= -420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011000; // iC=-1128 
vC = 14'b1111111011000011; // vC= -317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100000; // iC=-1184 
vC = 14'b1111111011011001; // vC= -295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011001; // iC=-1063 
vC = 14'b1111111001011110; // vC= -418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110010; // iC=-1102 
vC = 14'b1111111010110100; // vC= -332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100111; // iC=-1113 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011111; // iC=-1121 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100111; // iC=-1049 
vC = 14'b1111111001011100; // vC= -420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111110; // iC=-1090 
vC = 14'b1111111000111010; // vC= -454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111111; // iC=-1025 
vC = 14'b1111111000101111; // vC= -465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110100; // iC=-1036 
vC = 14'b1111111010100011; // vC= -349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001110; // iC=-1138 
vC = 14'b1111111011000011; // vC= -317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001010; // iC=-1078 
vC = 14'b1111111001011001; // vC= -423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010111; // iC=-1129 
vC = 14'b1111111000011011; // vC= -485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111001; // iC=-1095 
vC = 14'b1111111010000011; // vC= -381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111111; // iC=-1025 
vC = 14'b1111111010101010; // vC= -342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101110; // iC=-1042 
vC = 14'b1111111000011111; // vC= -481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110000; // iC=-1040 
vC = 14'b1111111010011001; // vC= -359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110111; // iC= -969 
vC = 14'b1111111001001010; // vC= -438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011000; // iC=-1128 
vC = 14'b1111111000001101; // vC= -499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001001; // iC=-1079 
vC = 14'b1111111000001101; // vC= -499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001111; // iC=-1009 
vC = 14'b1111111010010000; // vC= -368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110101; // iC=-1099 
vC = 14'b1111111010000101; // vC= -379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010001; // iC=-1007 
vC = 14'b1111111001111011; // vC= -389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110010; // iC=-1038 
vC = 14'b1111111000101011; // vC= -469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001111; // iC=-1009 
vC = 14'b1111111010001101; // vC= -371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111011; // iC= -965 
vC = 14'b1111111001110110; // vC= -394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011001; // iC=-1063 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000011; // iC=-1021 
vC = 14'b1111111001001100; // vC= -436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000110; // iC=-1082 
vC = 14'b1111111001011011; // vC= -421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101011; // iC=-1045 
vC = 14'b1111110111101011; // vC= -533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001110; // iC=-1074 
vC = 14'b1111111001000010; // vC= -446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110001; // iC=-1039 
vC = 14'b1111111000111111; // vC= -449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100100; // iC=-1052 
vC = 14'b1111111001100101; // vC= -411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101000; // iC=-1048 
vC = 14'b1111111001011001; // vC= -423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010011; // iC= -941 
vC = 14'b1111110111001101; // vC= -563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011110; // iC= -994 
vC = 14'b1111111000011011; // vC= -485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011000; // iC= -936 
vC = 14'b1111110111000010; // vC= -574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101100; // iC= -916 
vC = 14'b1111111001010100; // vC= -428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010100; // iC=-1004 
vC = 14'b1111110111000010; // vC= -574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010010; // iC= -942 
vC = 14'b1111111000111010; // vC= -454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000111; // iC=-1017 
vC = 14'b1111111000010000; // vC= -496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000101; // iC=-1019 
vC = 14'b1111110110111011; // vC= -581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110110; // iC=-1034 
vC = 14'b1111111000111101; // vC= -451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010101; // iC= -939 
vC = 14'b1111110111011101; // vC= -547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111000; // iC= -968 
vC = 14'b1111110111010100; // vC= -556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000100; // iC= -956 
vC = 14'b1111111000101101; // vC= -467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011010; // iC= -934 
vC = 14'b1111111000001101; // vC= -499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011100; // iC= -932 
vC = 14'b1111110111111111; // vC= -513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010101; // iC= -875 
vC = 14'b1111111000010110; // vC= -490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010000; // iC= -880 
vC = 14'b1111111000001011; // vC= -501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000101; // iC= -891 
vC = 14'b1111110110011010; // vC= -614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100001; // iC= -991 
vC = 14'b1111110111011011; // vC= -549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101010; // iC= -854 
vC = 14'b1111111000001101; // vC= -499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111110; // iC= -834 
vC = 14'b1111110110100011; // vC= -605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111011; // iC= -965 
vC = 14'b1111111000000100; // vC= -508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110000; // iC= -848 
vC = 14'b1111110110111010; // vC= -582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110001; // iC= -911 
vC = 14'b1111110110010011; // vC= -621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110100; // iC= -844 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101111; // iC= -849 
vC = 14'b1111110110010111; // vC= -617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010010; // iC= -814 
vC = 14'b1111110111001010; // vC= -566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100110; // iC= -922 
vC = 14'b1111111000001001; // vC= -503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111101; // iC= -899 
vC = 14'b1111110111001111; // vC= -561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000110; // iC= -954 
vC = 14'b1111110101111011; // vC= -645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001100; // iC= -948 
vC = 14'b1111110110111001; // vC= -583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001010; // iC= -886 
vC = 14'b1111110110110000; // vC= -592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111000; // iC= -840 
vC = 14'b1111110101100101; // vC= -667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100110; // iC= -858 
vC = 14'b1111110101111000; // vC= -648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101101; // iC= -851 
vC = 14'b1111110110111011; // vC= -581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110010; // iC= -910 
vC = 14'b1111110101011100; // vC= -676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000000; // iC= -768 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011100; // iC= -804 
vC = 14'b1111110110010100; // vC= -620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010111; // iC= -873 
vC = 14'b1111110110011010; // vC= -614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000010; // iC= -766 
vC = 14'b1111110101110010; // vC= -654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101111; // iC= -849 
vC = 14'b1111110101001000; // vC= -696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111001; // iC= -839 
vC = 14'b1111110110100001; // vC= -607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001101; // iC= -883 
vC = 14'b1111110101000001; // vC= -703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000101; // iC= -763 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100100; // iC= -796 
vC = 14'b1111110111010100; // vC= -556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111000; // iC= -776 
vC = 14'b1111110111001000; // vC= -568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011110; // iC= -738 
vC = 14'b1111110101011001; // vC= -679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100110; // iC= -858 
vC = 14'b1111110101000010; // vC= -702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001111; // iC= -753 
vC = 14'b1111110110101011; // vC= -597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010100; // iC= -876 
vC = 14'b1111110101111000; // vC= -648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100110; // iC= -730 
vC = 14'b1111110110001010; // vC= -630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111100; // iC= -836 
vC = 14'b1111110100111001; // vC= -711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011101; // iC= -739 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000101; // iC= -763 
vC = 14'b1111110110110101; // vC= -587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001100; // iC= -820 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111101; // iC= -707 
vC = 14'b1111110101100011; // vC= -669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100111; // iC= -729 
vC = 14'b1111110110110000; // vC= -592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101010; // iC= -790 
vC = 14'b1111110110011000; // vC= -616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011111; // iC= -801 
vC = 14'b1111110101010100; // vC= -684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000011; // iC= -765 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011011; // iC= -805 
vC = 14'b1111110100100001; // vC= -735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001000; // iC= -696 
vC = 14'b1111110100001100; // vC= -756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110110; // iC= -778 
vC = 14'b1111110101000010; // vC= -702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000101; // iC= -699 
vC = 14'b1111110100011000; // vC= -744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010010; // iC= -750 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111010; // iC= -774 
vC = 14'b1111110100011100; // vC= -740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000111; // iC= -697 
vC = 14'b1111110100011001; // vC= -743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011011; // iC= -677 
vC = 14'b1111110100011110; // vC= -738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101110; // iC= -786 
vC = 14'b1111110101010001; // vC= -687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110111; // iC= -777 
vC = 14'b1111110101011001; // vC= -679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110011; // iC= -653 
vC = 14'b1111110100101110; // vC= -722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100100; // iC= -668 
vC = 14'b1111110100001100; // vC= -756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010001; // iC= -687 
vC = 14'b1111110011111100; // vC= -772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101001; // iC= -727 
vC = 14'b1111110011101100; // vC= -788 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000010; // iC= -766 
vC = 14'b1111110100111010; // vC= -710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100100; // iC= -732 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100000; // iC= -608 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100010; // iC= -670 
vC = 14'b1111110101001010; // vC= -694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100011; // iC= -605 
vC = 14'b1111110011101001; // vC= -791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011111; // iC= -737 
vC = 14'b1111110101010101; // vC= -683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011001; // iC= -743 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011110; // iC= -610 
vC = 14'b1111110100110111; // vC= -713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011001; // iC= -615 
vC = 14'b1111110101100001; // vC= -671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101000; // iC= -728 
vC = 14'b1111110100010111; // vC= -745 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b1111110101001010; // vC= -694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000111; // iC= -569 
vC = 14'b1111110011100111; // vC= -793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111110; // iC= -578 
vC = 14'b1111110101100011; // vC= -669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010001; // iC= -559 
vC = 14'b1111110101011010; // vC= -678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010100; // iC= -620 
vC = 14'b1111110100101101; // vC= -723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001111; // iC= -625 
vC = 14'b1111110101011001; // vC= -679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111101; // iC= -643 
vC = 14'b1111110100011100; // vC= -740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001000; // iC= -632 
vC = 14'b1111110100100111; // vC= -729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001110; // iC= -562 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111111; // iC= -641 
vC = 14'b1111110100000100; // vC= -764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001001; // iC= -567 
vC = 14'b1111110100111000; // vC= -712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100111; // iC= -537 
vC = 14'b1111110011111010; // vC= -774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101001; // iC= -535 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000001; // iC= -639 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111110; // iC= -642 
vC = 14'b1111110011110100; // vC= -780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010100; // iC= -556 
vC = 14'b1111110011100010; // vC= -798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001010; // iC= -566 
vC = 14'b1111110100111000; // vC= -712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111011; // iC= -517 
vC = 14'b1111110100101011; // vC= -725 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100010; // iC= -606 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100110; // iC= -538 
vC = 14'b1111110010100111; // vC= -857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111101; // iC= -579 
vC = 14'b1111110100011101; // vC= -739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b1111110010101000; // vC= -856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101100; // iC= -468 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001111; // iC= -497 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001101; // iC= -563 
vC = 14'b1111110010011101; // vC= -867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110100; // iC= -588 
vC = 14'b1111110011100100; // vC= -796 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000000; // iC= -576 
vC = 14'b1111110100001001; // vC= -759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011000; // iC= -488 
vC = 14'b1111110010010110; // vC= -874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111100; // iC= -452 
vC = 14'b1111110011111100; // vC= -772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100100; // iC= -540 
vC = 14'b1111110100011001; // vC= -743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110100; // iC= -524 
vC = 14'b1111110011110111; // vC= -777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001000; // iC= -568 
vC = 14'b1111110011010100; // vC= -812 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101110; // iC= -530 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001010; // iC= -566 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100010; // iC= -414 
vC = 14'b1111110011000111; // vC= -825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111110; // iC= -450 
vC = 14'b1111110010010111; // vC= -873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110111; // iC= -457 
vC = 14'b1111110011100110; // vC= -794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011110; // iC= -482 
vC = 14'b1111110100000011; // vC= -765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010100; // iC= -556 
vC = 14'b1111110010010101; // vC= -875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101010; // iC= -406 
vC = 14'b1111110010010000; // vC= -880 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110101; // iC= -523 
vC = 14'b1111110010111110; // vC= -834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110000; // iC= -400 
vC = 14'b1111110010110001; // vC= -847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100011; // iC= -413 
vC = 14'b1111110010100111; // vC= -857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000101; // iC= -507 
vC = 14'b1111110011011100; // vC= -804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000010; // iC= -510 
vC = 14'b1111110011110101; // vC= -779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001000; // iC= -504 
vC = 14'b1111110100001110; // vC= -754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011101; // iC= -419 
vC = 14'b1111110011001111; // vC= -817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111101; // iC= -515 
vC = 14'b1111110011000000; // vC= -832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000011; // iC= -381 
vC = 14'b1111110010001100; // vC= -884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110001; // iC= -463 
vC = 14'b1111110011000011; // vC= -829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110000; // iC= -464 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000111; // iC= -441 
vC = 14'b1111110011101101; // vC= -787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010001; // iC= -431 
vC = 14'b1111110010001110; // vC= -882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011000; // iC= -424 
vC = 14'b1111110001111011; // vC= -901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001001; // iC= -375 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010101; // iC= -363 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100010; // iC= -414 
vC = 14'b1111110010001110; // vC= -882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111110; // iC= -322 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111000; // iC= -392 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000111; // iC= -313 
vC = 14'b1111110011011110; // vC= -802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111011; // iC= -453 
vC = 14'b1111110010010000; // vC= -880 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011010; // iC= -358 
vC = 14'b1111110010000110; // vC= -890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010111; // iC= -361 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100001; // iC= -415 
vC = 14'b1111110011110101; // vC= -779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001010; // iC= -310 
vC = 14'b1111110010010010; // vC= -878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010000; // iC= -304 
vC = 14'b1111110001011001; // vC= -935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000010; // iC= -318 
vC = 14'b1111110001111100; // vC= -900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000100; // iC= -380 
vC = 14'b1111110011011111; // vC= -801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000011; // iC= -317 
vC = 14'b1111110010000100; // vC= -892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101100; // iC= -340 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111001; // iC= -327 
vC = 14'b1111110011101101; // vC= -787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110001; // iC= -271 
vC = 14'b1111110010100011; // vC= -861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110010; // iC= -398 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111000; // iC= -264 
vC = 14'b1111110011000011; // vC= -829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101110; // iC= -338 
vC = 14'b1111110011011101; // vC= -803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001110; // iC= -370 
vC = 14'b1111110001110110; // vC= -906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101111; // iC= -337 
vC = 14'b1111110001101101; // vC= -915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101001; // iC= -343 
vC = 14'b1111110001001010; // vC= -950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000111; // iC= -249 
vC = 14'b1111110011000101; // vC= -827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101110; // iC= -274 
vC = 14'b1111110010010001; // vC= -879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101011; // iC= -213 
vC = 14'b1111110001111110; // vC= -898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000001; // iC= -191 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101111; // iC= -273 
vC = 14'b1111110010101100; // vC= -852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000100; // iC= -188 
vC = 14'b1111110010010001; // vC= -879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011101; // iC= -163 
vC = 14'b1111110010101110; // vC= -850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001100; // iC= -180 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110100; // iC= -140 
vC = 14'b1111110010110001; // vC= -847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101101; // iC= -211 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100111; // iC=  -89 
vC = 14'b1111110010001000; // vC= -888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101111; // iC= -209 
vC = 14'b1111110011010110; // vC= -810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110101; // iC= -203 
vC = 14'b1111110010001111; // vC= -881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101100; // iC=  -84 
vC = 14'b1111110011000010; // vC= -830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011110; // iC=  -34 
vC = 14'b1111110010101101; // vC= -851 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011011; // iC= -101 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000000; // iC= -128 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100000; // iC=  -96 
vC = 14'b1111110011010001; // vC= -815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110100; // iC= -140 
vC = 14'b1111110010100001; // vC= -863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000100; // iC=  -60 
vC = 14'b1111110001011001; // vC= -935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100101; // iC=  -91 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000101; // iC=    5 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101110; // iC=  -82 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110110; // iC=  -10 
vC = 14'b1111110000111100; // vC= -964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100000; // iC=   32 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101000; // iC=  -24 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001010; // iC=   10 
vC = 14'b1111110010001000; // vC= -888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001100; // iC=   12 
vC = 14'b1111110001101111; // vC= -913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100001; // iC=  161 
vC = 14'b1111110010100011; // vC= -861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100001; // iC=   97 
vC = 14'b1111110010100000; // vC= -864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100000; // iC=  160 
vC = 14'b1111110010110101; // vC= -843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101101; // iC=  173 
vC = 14'b1111110010000010; // vC= -894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100011; // iC=   99 
vC = 14'b1111110011000010; // vC= -830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000001; // iC=  129 
vC = 14'b1111110001111100; // vC= -900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001111; // iC=  207 
vC = 14'b1111110010011110; // vC= -866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001011; // iC=  203 
vC = 14'b1111110011000010; // vC= -830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100000; // iC=  160 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110011; // iC=  243 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101011; // iC=  363 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100111; // iC=  231 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001010; // iC=  330 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010110; // iC=  342 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111011; // iC=  443 
vC = 14'b1111110001011100; // vC= -932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010101; // iC=  469 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010000; // iC=  464 
vC = 14'b1111110010000010; // vC= -894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101111; // iC=  367 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001000; // iC=  520 
vC = 14'b1111110010101111; // vC= -849 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011111; // iC=  479 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101101; // iC=  493 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001110; // iC=  590 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010010; // iC=  594 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101010; // iC=  490 
vC = 14'b1111110010111010; // vC= -838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101110; // iC=  622 
vC = 14'b1111110001111101; // vC= -899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100111; // iC=  551 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010011; // iC=  659 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001111; // iC=  719 
vC = 14'b1111110011011101; // vC= -803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011011; // iC=  667 
vC = 14'b1111110001101111; // vC= -913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010101; // iC=  725 
vC = 14'b1111110010100011; // vC= -861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111111; // iC=  767 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100001; // iC=  801 
vC = 14'b1111110010000110; // vC= -890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100101; // iC=  677 
vC = 14'b1111110011000101; // vC= -827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001100; // iC=  780 
vC = 14'b1111110010010010; // vC= -878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001011; // iC=  779 
vC = 14'b1111110010000101; // vC= -891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101100; // iC=  876 
vC = 14'b1111110100000111; // vC= -761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010000; // iC=  848 
vC = 14'b1111110011001111; // vC= -817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110000; // iC=  816 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101001; // iC=  809 
vC = 14'b1111110011001110; // vC= -818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000000; // iC=  832 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b1111110010010110; // vC= -874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100011; // iC=  931 
vC = 14'b1111110011000111; // vC= -825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001000; // iC=  968 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010101; // iC= 1045 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011111; // iC= 1055 
vC = 14'b1111110010110001; // vC= -847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010100; // iC=  980 
vC = 14'b1111110011000010; // vC= -830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011100; // iC=  988 
vC = 14'b1111110100010111; // vC= -745 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001100; // iC=  972 
vC = 14'b1111110011001011; // vC= -821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100101; // iC=  997 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110010; // iC= 1138 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000001; // iC= 1089 
vC = 14'b1111110100101101; // vC= -723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111011; // iC= 1147 
vC = 14'b1111110100011101; // vC= -739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110101; // iC= 1205 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010010; // iC= 1106 
vC = 14'b1111110100000100; // vC= -764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b1111110101001101; // vC= -691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111111; // iC= 1151 
vC = 14'b1111110011101001; // vC= -791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100001; // iC= 1249 
vC = 14'b1111110100101001; // vC= -727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100000; // iC= 1312 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011001; // iC= 1177 
vC = 14'b1111110101011010; // vC= -678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000001; // iC= 1345 
vC = 14'b1111110011101000; // vC= -792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000110; // iC= 1286 
vC = 14'b1111110100001111; // vC= -753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101110; // iC= 1326 
vC = 14'b1111110011101110; // vC= -786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101111; // iC= 1263 
vC = 14'b1111110101011111; // vC= -673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010100; // iC= 1364 
vC = 14'b1111110011111100; // vC= -772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011001; // iC= 1369 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000001; // iC= 1409 
vC = 14'b1111110100100100; // vC= -732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100010; // iC= 1314 
vC = 14'b1111110101110111; // vC= -649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110111; // iC= 1335 
vC = 14'b1111110101110000; // vC= -656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010000; // iC= 1424 
vC = 14'b1111110100100010; // vC= -734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000110; // iC= 1414 
vC = 14'b1111110100001111; // vC= -753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011001; // iC= 1433 
vC = 14'b1111110101010100; // vC= -684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011001; // iC= 1497 
vC = 14'b1111110101110111; // vC= -649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110111; // iC= 1463 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101111; // iC= 1455 
vC = 14'b1111110100101110; // vC= -722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010010; // iC= 1426 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b1111110110001101; // vC= -627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b1111110100111010; // vC= -710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101100; // iC= 1452 
vC = 14'b1111110101001000; // vC= -696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010010; // iC= 1490 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001001; // iC= 1481 
vC = 14'b1111110110011111; // vC= -609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100100; // iC= 1572 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111111; // iC= 1599 
vC = 14'b1111110110001100; // vC= -628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100011; // iC= 1571 
vC = 14'b1111110101010001; // vC= -687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001101; // iC= 1549 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010010; // iC= 1618 
vC = 14'b1111110110111110; // vC= -578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110010; // iC= 1522 
vC = 14'b1111110111001110; // vC= -562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110010; // iC= 1522 
vC = 14'b1111110101011010; // vC= -678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b1111110111001110; // vC= -562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010000; // iC= 1552 
vC = 14'b1111110101110101; // vC= -651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111000; // iC= 1592 
vC = 14'b1111110111111110; // vC= -514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010010; // iC= 1554 
vC = 14'b1111110111100010; // vC= -542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b1111110110000111; // vC= -633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110000; // iC= 1584 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001111; // iC= 1679 
vC = 14'b1111110111010110; // vC= -554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b1111110111110011; // vC= -525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010111; // iC= 1623 
vC = 14'b1111111000001110; // vC= -498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b1111110110010101; // vC= -619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010001; // iC= 1745 
vC = 14'b1111110110110100; // vC= -588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b1111111000110010; // vC= -462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100000; // iC= 1632 
vC = 14'b1111111000000100; // vC= -508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011110; // iC= 1630 
vC = 14'b1111110110110110; // vC= -586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011000; // iC= 1688 
vC = 14'b1111110111111000; // vC= -520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100110; // iC= 1638 
vC = 14'b1111111000110000; // vC= -464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b1111110111010001; // vC= -559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111110; // iC= 1662 
vC = 14'b1111110111000011; // vC= -573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011101; // iC= 1693 
vC = 14'b1111111000010010; // vC= -494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b1111110111010100; // vC= -556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b1111111000001111; // vC= -497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b1111111001100110; // vC= -410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100111; // iC= 1639 
vC = 14'b1111110111110100; // vC= -524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110110; // iC= 1654 
vC = 14'b1111111001100111; // vC= -409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000010; // iC= 1794 
vC = 14'b1111111001110110; // vC= -394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100101; // iC= 1637 
vC = 14'b1111111001111001; // vC= -391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b1111111000101101; // vC= -467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111111001110001; // vC= -399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111111001101100; // vC= -404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b1111111001100100; // vC= -412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111111010100010; // vC= -350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101011; // iC= 1643 
vC = 14'b1111111001011011; // vC= -421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000010; // iC= 1794 
vC = 14'b1111111001110111; // vC= -393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b1111111001001010; // vC= -438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b1111111010001100; // vC= -372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101011; // iC= 1643 
vC = 14'b1111111001001000; // vC= -440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000000; // iC= 1792 
vC = 14'b1111111010001011; // vC= -373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b1111111001010000; // vC= -432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000100; // iC= 1668 
vC = 14'b1111111010101111; // vC= -337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001011; // iC= 1739 
vC = 14'b1111111010000111; // vC= -377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b1111111010010001; // vC= -367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b1111111011111101; // vC= -259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101001; // iC= 1705 
vC = 14'b1111111011000011; // vC= -317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100110; // iC= 1638 
vC = 14'b1111111010000100; // vC= -380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001011; // iC= 1739 
vC = 14'b1111111011010111; // vC= -297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110011; // iC= 1651 
vC = 14'b1111111100010011; // vC= -237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001101; // iC= 1677 
vC = 14'b1111111100001101; // vC= -243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000110; // iC= 1734 
vC = 14'b1111111011100100; // vC= -284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b1111111010100111; // vC= -345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010011; // iC= 1747 
vC = 14'b1111111011101100; // vC= -276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b1111111100010001; // vC= -239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010100; // iC= 1748 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111110; // iC= 1726 
vC = 14'b1111111100111101; // vC= -195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011000; // iC= 1624 
vC = 14'b1111111101001000; // vC= -184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110000; // iC= 1648 
vC = 14'b1111111100101000; // vC= -216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011100; // iC= 1628 
vC = 14'b1111111100111010; // vC= -198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b1111111100011101; // vC= -227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110111; // iC= 1655 
vC = 14'b1111111100001111; // vC= -241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110010; // iC= 1650 
vC = 14'b1111111100010100; // vC= -236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100100; // iC= 1636 
vC = 14'b1111111101011011; // vC= -165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100010; // iC= 1698 
vC = 14'b1111111100010100; // vC= -236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110010; // iC= 1650 
vC = 14'b1111111100101100; // vC= -212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b1111111100110001; // vC= -207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b1111111100101001; // vC= -215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101001; // iC= 1641 
vC = 14'b1111111100111100; // vC= -196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101001; // iC= 1641 
vC = 14'b1111111110011001; // vC= -103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b1111111101100011; // vC= -157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000001; // iC= 1665 
vC = 14'b1111111110000001; // vC= -127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011111; // iC= 1695 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110000; // iC= 1648 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111010; // iC= 1594 
vC = 14'b1111111101000101; // vC= -187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110010; // iC= 1650 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b1111111110011111; // vC=  -97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b1111111101111110; // vC= -130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111111; // iC= 1663 
vC = 14'b1111111110110110; // vC=  -74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111111; // iC= 1599 
vC = 14'b1111111110101101; // vC=  -83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011101; // iC= 1629 
vC = 14'b1111111101001110; // vC= -178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b1111111111101001; // vC=  -23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001000; // iC= 1672 
vC = 14'b1111111101101111; // vC= -145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001010; // iC= 1610 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010110; // iC= 1686 
vC = 14'b1111111111100011; // vC=  -29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b1111111110001100; // vC= -116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b1111111111010110; // vC=  -42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001001; // iC= 1609 
vC = 14'b1111111110100101; // vC=  -91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b1111111111111001; // vC=   -7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000000; // iC= 1600 
vC = 14'b1111111111011100; // vC=  -36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b1111111110100000; // vC=  -96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b1111111110111100; // vC=  -68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100111; // iC= 1639 
vC = 14'b1111111111011000; // vC=  -40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001100; // iC= 1612 
vC = 14'b0000000000110001; // vC=   49 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100101; // iC= 1573 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000000; // iC= 1664 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010110; // iC= 1558 
vC = 14'b1111111111100001; // vC=  -31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110101; // iC= 1589 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b0000000000010101; // vC=   21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b1111111111001110; // vC=  -50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b0000000000011001; // vC=   25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b0000000000001101; // vC=   13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b0000000001010011; // vC=   83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b1111111111111100; // vC=   -4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b0000000000011101; // vC=   29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010101; // iC= 1685 
vC = 14'b0000000000101000; // vC=   40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b0000000001100111; // vC=  103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000000; // iC= 1664 
vC = 14'b0000000000101100; // vC=   44 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110101; // iC= 1525 
vC = 14'b0000000000111001; // vC=   57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100100; // iC= 1636 
vC = 14'b0000000000010111; // vC=   23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b0000000001011100; // vC=   92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110011; // iC= 1523 
vC = 14'b0000000001101000; // vC=  104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001001; // iC= 1609 
vC = 14'b0000000010001010; // vC=  138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110000; // iC= 1520 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110111; // iC= 1591 
vC = 14'b0000000000011010; // vC=   26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100101; // iC= 1573 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000010; // iC= 1538 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b0000000000101100; // vC=   44 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101111; // iC= 1647 
vC = 14'b0000000001111101; // vC=  125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100100; // iC= 1572 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101011; // iC= 1579 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010011; // iC= 1491 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010001; // iC= 1553 
vC = 14'b0000000010100110; // vC=  166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100100; // iC= 1572 
vC = 14'b0000000010111011; // vC=  187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b0000000010101100; // vC=  172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011001; // iC= 1625 
vC = 14'b0000000001111011; // vC=  123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010111; // iC= 1495 
vC = 14'b0000000010111100; // vC=  188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010100; // iC= 1556 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101001; // iC= 1513 
vC = 14'b0000000011010111; // vC=  215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110010; // iC= 1522 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110110; // iC= 1590 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010001; // iC= 1489 
vC = 14'b0000000011111010; // vC=  250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000110; // iC= 1478 
vC = 14'b0000000001111011; // vC=  123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110101; // iC= 1589 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000000100001101; // vC=  269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110111; // iC= 1463 
vC = 14'b0000000010001100; // vC=  140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b0000000100010100; // vC=  276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111001; // iC= 1593 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110011; // iC= 1459 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101011; // iC= 1451 
vC = 14'b0000000010001001; // vC=  137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011110; // iC= 1502 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110010; // iC= 1522 
vC = 14'b0000000010010110; // vC=  150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110101; // iC= 1525 
vC = 14'b0000000011100001; // vC=  225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010000; // iC= 1488 
vC = 14'b0000000100110000; // vC=  304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100000; // iC= 1504 
vC = 14'b0000000101000101; // vC=  325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010110; // iC= 1430 
vC = 14'b0000000100111110; // vC=  318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101001; // iC= 1513 
vC = 14'b0000000100010111; // vC=  279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001110; // iC= 1550 
vC = 14'b0000000101000001; // vC=  321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000011; // iC= 1475 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100110; // iC= 1510 
vC = 14'b0000000100111010; // vC=  314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000010; // iC= 1538 
vC = 14'b0000000100000100; // vC=  260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111111; // iC= 1407 
vC = 14'b0000000101100101; // vC=  357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110110; // iC= 1462 
vC = 14'b0000000100100110; // vC=  294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011010; // iC= 1562 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111000; // iC= 1400 
vC = 14'b0000000101000111; // vC=  327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011101; // iC= 1501 
vC = 14'b0000000011101110; // vC=  238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011101; // iC= 1437 
vC = 14'b0000000100101010; // vC=  298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101111; // iC= 1391 
vC = 14'b0000000100001110; // vC=  270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110000; // iC= 1520 
vC = 14'b0000000100101101; // vC=  301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111111; // iC= 1471 
vC = 14'b0000000100111111; // vC=  319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100100; // iC= 1380 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101110; // iC= 1518 
vC = 14'b0000000100100000; // vC=  288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b0000000110001011; // vC=  395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010110; // iC= 1430 
vC = 14'b0000000101010110; // vC=  342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111001; // iC= 1465 
vC = 14'b0000000110000010; // vC=  386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110110; // iC= 1398 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000010; // iC= 1474 
vC = 14'b0000000101001111; // vC=  335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110011; // iC= 1459 
vC = 14'b0000000100110001; // vC=  305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110111; // iC= 1463 
vC = 14'b0000000100101011; // vC=  299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010111; // iC= 1367 
vC = 14'b0000000110010111; // vC=  407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001110; // iC= 1486 
vC = 14'b0000000101100111; // vC=  359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001111; // iC= 1359 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100111; // iC= 1447 
vC = 14'b0000000110001110; // vC=  398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001010; // iC= 1418 
vC = 14'b0000000101000101; // vC=  325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010101; // iC= 1493 
vC = 14'b0000000110000010; // vC=  386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100000; // iC= 1376 
vC = 14'b0000000111010001; // vC=  465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111101; // iC= 1405 
vC = 14'b0000000110001001; // vC=  393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110110; // iC= 1398 
vC = 14'b0000000111000001; // vC=  449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100100; // iC= 1380 
vC = 14'b0000000111001100; // vC=  460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000011; // iC= 1475 
vC = 14'b0000000110011100; // vC=  412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010010; // iC= 1362 
vC = 14'b0000000101110110; // vC=  374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011101; // iC= 1437 
vC = 14'b0000000110000001; // vC=  385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110000; // iC= 1328 
vC = 14'b0000000110010000; // vC=  400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100010; // iC= 1442 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110001; // iC= 1457 
vC = 14'b0000000110010011; // vC=  403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111001; // iC= 1337 
vC = 14'b0000000111110101; // vC=  501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110111; // iC= 1335 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101101; // iC= 1389 
vC = 14'b0000000111011101; // vC=  477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101100; // iC= 1324 
vC = 14'b0000001000010100; // vC=  532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001000; // iC= 1416 
vC = 14'b0000000110011111; // vC=  415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011000; // iC= 1432 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011001; // iC= 1433 
vC = 14'b0000000110101000; // vC=  424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001010; // iC= 1354 
vC = 14'b0000000110100110; // vC=  422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000001000100100; // vC=  548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011000; // iC= 1368 
vC = 14'b0000001000100111; // vC=  551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111001; // iC= 1273 
vC = 14'b0000001000000111; // vC=  519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110010; // iC= 1330 
vC = 14'b0000000111010011; // vC=  467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010001; // iC= 1361 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001000; // iC= 1416 
vC = 14'b0000001000101111; // vC=  559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010100; // iC= 1364 
vC = 14'b0000001000011000; // vC=  536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001011; // iC= 1291 
vC = 14'b0000001000011010; // vC=  538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100101; // iC= 1317 
vC = 14'b0000001000001110; // vC=  526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000111; // iC= 1287 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000001; // iC= 1345 
vC = 14'b0000000110111010; // vC=  442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011000; // iC= 1240 
vC = 14'b0000001000101010; // vC=  554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000011; // iC= 1283 
vC = 14'b0000001001001110; // vC=  590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000111; // iC= 1287 
vC = 14'b0000001000100100; // vC=  548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101100; // iC= 1260 
vC = 14'b0000001001100100; // vC=  612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011001; // iC= 1305 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011101; // iC= 1309 
vC = 14'b0000001000100111; // vC=  551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100111; // iC= 1255 
vC = 14'b0000001001000001; // vC=  577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010000; // iC= 1296 
vC = 14'b0000001001011101; // vC=  605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110110; // iC= 1334 
vC = 14'b0000001001001101; // vC=  589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001101; // iC= 1229 
vC = 14'b0000001001001111; // vC=  591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000110; // iC= 1350 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100011; // iC= 1251 
vC = 14'b0000001000010100; // vC=  532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000111; // iC= 1223 
vC = 14'b0000001000001000; // vC=  520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000010; // iC= 1346 
vC = 14'b0000000111111010; // vC=  506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010101; // iC= 1301 
vC = 14'b0000000111111011; // vC=  507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010101; // iC= 1301 
vC = 14'b0000001001110010; // vC=  626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110101; // iC= 1205 
vC = 14'b0000001001001001; // vC=  585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101110; // iC= 1198 
vC = 14'b0000001001110110; // vC=  630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100010; // iC= 1314 
vC = 14'b0000001010001110; // vC=  654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001011; // iC= 1291 
vC = 14'b0000001000101110; // vC=  558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111011; // iC= 1211 
vC = 14'b0000001001111001; // vC=  633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101001; // iC= 1257 
vC = 14'b0000001000011011; // vC=  539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011100; // iC= 1180 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100000; // iC= 1248 
vC = 14'b0000001000101011; // vC=  555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001010; // iC= 1226 
vC = 14'b0000001000100101; // vC=  549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011100; // iC= 1180 
vC = 14'b0000001001111010; // vC=  634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101001; // iC= 1257 
vC = 14'b0000001000101110; // vC=  558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111100; // iC= 1148 
vC = 14'b0000001010011010; // vC=  666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011000; // iC= 1240 
vC = 14'b0000001001001111; // vC=  591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000110; // iC= 1222 
vC = 14'b0000001010011110; // vC=  670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110001; // iC= 1201 
vC = 14'b0000001010110111; // vC=  695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011000; // iC= 1176 
vC = 14'b0000001001111111; // vC=  639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110011; // iC= 1203 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001000; // iC= 1224 
vC = 14'b0000001001111001; // vC=  633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100010; // iC= 1186 
vC = 14'b0000001001110000; // vC=  624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111100; // iC= 1148 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100101; // iC= 1125 
vC = 14'b0000001010101100; // vC=  684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101111; // iC= 1135 
vC = 14'b0000001010101110; // vC=  686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010001; // iC= 1105 
vC = 14'b0000001010110010; // vC=  690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100100; // iC= 1188 
vC = 14'b0000001010101011; // vC=  683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001001; // iC= 1161 
vC = 14'b0000001001110110; // vC=  630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111101; // iC= 1149 
vC = 14'b0000001011111001; // vC=  761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011010; // iC= 1178 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111100; // iC= 1084 
vC = 14'b0000001100000110; // vC=  774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111100; // iC= 1212 
vC = 14'b0000001001111111; // vC=  639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111100; // iC= 1148 
vC = 14'b0000001010101011; // vC=  683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111111; // iC= 1215 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101111; // iC= 1199 
vC = 14'b0000001011010010; // vC=  722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100000; // iC= 1056 
vC = 14'b0000001010101111; // vC=  687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b0000001010100010; // vC=  674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100010; // iC= 1058 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011000; // iC= 1176 
vC = 14'b0000001010100101; // vC=  677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101001; // iC= 1065 
vC = 14'b0000001011001110; // vC=  718 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111011; // iC= 1083 
vC = 14'b0000001011001101; // vC=  717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101100; // iC= 1068 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111010; // iC= 1146 
vC = 14'b0000001100011010; // vC=  794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000110; // iC= 1094 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000001; // iC= 1025 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000101; // iC= 1093 
vC = 14'b0000001010111000; // vC=  696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111001; // iC= 1017 
vC = 14'b0000001100011010; // vC=  794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001101; // iC= 1101 
vC = 14'b0000001100101100; // vC=  812 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000000; // iC= 1088 
vC = 14'b0000001011101001; // vC=  745 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110101; // iC= 1141 
vC = 14'b0000001011111110; // vC=  766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000000; // iC= 1088 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110111; // iC= 1015 
vC = 14'b0000001100000010; // vC=  770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110011; // iC= 1075 
vC = 14'b0000001010111000; // vC=  696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110010; // iC= 1074 
vC = 14'b0000001011110010; // vC=  754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110010; // iC= 1074 
vC = 14'b0000001101011001; // vC=  857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001011; // iC= 1099 
vC = 14'b0000001011111100; // vC=  764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100100; // iC= 1124 
vC = 14'b0000001100001001; // vC=  777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111010; // iC= 1082 
vC = 14'b0000001100000001; // vC=  769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001000; // iC= 1096 
vC = 14'b0000001011001110; // vC=  718 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010001; // iC= 1105 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101111; // iC= 1071 
vC = 14'b0000001100111011; // vC=  827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111010; // iC= 1018 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000100; // iC= 1092 
vC = 14'b0000001101011100; // vC=  860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111100; // iC=  956 
vC = 14'b0000001100110010; // vC=  818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101111; // iC= 1071 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111100; // iC= 1020 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011000; // iC=  984 
vC = 14'b0000001100101111; // vC=  815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101011; // iC= 1003 
vC = 14'b0000001101110000; // vC=  880 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001011; // iC=  971 
vC = 14'b0000001101011010; // vC=  858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010000; // iC=  912 
vC = 14'b0000001100101010; // vC=  810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101011; // iC=  939 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100001; // iC= 1057 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010111; // iC=  983 
vC = 14'b0000001100011111; // vC=  799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000011; // iC=  963 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110010; // iC=  946 
vC = 14'b0000001101001111; // vC=  847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011100; // iC=  924 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011110; // iC=  926 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100110; // iC=  998 
vC = 14'b0000001101000000; // vC=  832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000111; // iC=  903 
vC = 14'b0000001100010111; // vC=  791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101100; // iC= 1004 
vC = 14'b0000001101101100; // vC=  876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101000; // iC=  936 
vC = 14'b0000001100011101; // vC=  797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111010; // iC=  954 
vC = 14'b0000001101111000; // vC=  888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001110; // iC=  974 
vC = 14'b0000001100111000; // vC=  824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111111; // iC=  959 
vC = 14'b0000001101101000; // vC=  872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001011; // iC=  907 
vC = 14'b0000001101000001; // vC=  833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010101; // iC=  981 
vC = 14'b0000001101010001; // vC=  849 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110101; // iC=  885 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001100; // iC=  908 
vC = 14'b0000001100100111; // vC=  807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001110; // iC=  846 
vC = 14'b0000001101010000; // vC=  848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111001; // iC=  825 
vC = 14'b0000001101101000; // vC=  872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110010; // iC=  946 
vC = 14'b0000001101111110; // vC=  894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000011; // iC=  899 
vC = 14'b0000001101010111; // vC=  855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100011; // iC=  931 
vC = 14'b0000001100110101; // vC=  821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101010; // iC=  938 
vC = 14'b0000001101110011; // vC=  883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000010; // iC=  834 
vC = 14'b0000001101111110; // vC=  894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001011; // iC=  907 
vC = 14'b0000001110011111; // vC=  927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100001; // iC=  801 
vC = 14'b0000001101101110; // vC=  878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000011; // iC=  835 
vC = 14'b0000001110000110; // vC=  902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001110; // iC=  910 
vC = 14'b0000001110101101; // vC=  941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001110; // iC=  782 
vC = 14'b0000001110000101; // vC=  901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100011; // iC=  803 
vC = 14'b0000001111011110; // vC=  990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000000; // iC=  896 
vC = 14'b0000001110110100; // vC=  948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000011; // iC=  835 
vC = 14'b0000001110101101; // vC=  941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111000; // iC=  824 
vC = 14'b0000001111001111; // vC=  975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001101; // iC=  845 
vC = 14'b0000001110010011; // vC=  915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111000; // iC=  824 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111110; // iC=  766 
vC = 14'b0000001110100011; // vC=  931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000001; // iC=  897 
vC = 14'b0000001110001011; // vC=  907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111001; // iC=  889 
vC = 14'b0000001101101011; // vC=  875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001110; // iC=  782 
vC = 14'b0000001110011101; // vC=  925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111000; // iC=  760 
vC = 14'b0000001110111111; // vC=  959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100101; // iC=  741 
vC = 14'b0000001111110010; // vC= 1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011100; // iC=  860 
vC = 14'b0000001110000010; // vC=  898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010111; // iC=  791 
vC = 14'b0000001110100000; // vC=  928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111101; // iC=  829 
vC = 14'b0000001111000010; // vC=  962 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001010; // iC=  714 
vC = 14'b0000001111111010; // vC= 1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001011; // iC=  715 
vC = 14'b0000001110011010; // vC=  922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110011; // iC=  755 
vC = 14'b0000001111110100; // vC= 1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110001; // iC=  817 
vC = 14'b0000001110010111; // vC=  919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010011; // iC=  787 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010111; // iC=  791 
vC = 14'b0000001110110100; // vC=  948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101111; // iC=  687 
vC = 14'b0000001110011000; // vC=  920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000100; // iC=  772 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001011; // iC=  715 
vC = 14'b0000001110010001; // vC=  913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110001; // iC=  689 
vC = 14'b0000001111101001; // vC= 1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100100; // iC=  740 
vC = 14'b0000001111000110; // vC=  966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111101; // iC=  701 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111010; // iC=  762 
vC = 14'b0000001110000010; // vC=  898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001100; // iC=  780 
vC = 14'b0000001110010001; // vC=  913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110011; // iC=  691 
vC = 14'b0000001110001011; // vC=  907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101111; // iC=  751 
vC = 14'b0000001111011101; // vC=  989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110110; // iC=  758 
vC = 14'b0000001110010110; // vC=  918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011001; // iC=  729 
vC = 14'b0000001111001000; // vC=  968 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000000; // iC=  640 
vC = 14'b0000001110101010; // vC=  938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b0000010000100111; // vC= 1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000011; // iC=  707 
vC = 14'b0000001111010101; // vC=  981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100101; // iC=  613 
vC = 14'b0000001111111101; // vC= 1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101100; // iC=  748 
vC = 14'b0000001110101101; // vC=  941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101101; // iC=  749 
vC = 14'b0000010000110011; // vC= 1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010110; // iC=  726 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101000; // iC=  616 
vC = 14'b0000001111101100; // vC= 1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011111; // iC=  607 
vC = 14'b0000001111000001; // vC=  961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000110; // iC=  646 
vC = 14'b0000001111101101; // vC= 1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110111; // iC=  695 
vC = 14'b0000001110101100; // vC=  940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001101; // iC=  717 
vC = 14'b0000001111111011; // vC= 1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001101; // iC=  589 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110001; // iC=  625 
vC = 14'b0000001110110110; // vC=  950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100110; // iC=  678 
vC = 14'b0000010000010000; // vC= 1040 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100010; // iC=  610 
vC = 14'b0000001111010011; // vC=  979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001010; // iC=  586 
vC = 14'b0000010000000110; // vC= 1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100100; // iC=  676 
vC = 14'b0000010001000000; // vC= 1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000100; // iC=  580 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001100; // iC=  652 
vC = 14'b0000001111001111; // vC=  975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111011; // iC=  635 
vC = 14'b0000001111011010; // vC=  986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010110; // iC=  662 
vC = 14'b0000010000000100; // vC= 1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000001; // iC=  577 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001010; // iC=  522 
vC = 14'b0000010001010101; // vC= 1109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111000; // iC=  568 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101001; // iC=  617 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000101; // iC=  645 
vC = 14'b0000001111111000; // vC= 1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101001; // iC=  617 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000101; // iC=  581 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111101; // iC=  509 
vC = 14'b0000010001100000; // vC= 1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011110; // iC=  542 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110000; // iC=  560 
vC = 14'b0000010000011100; // vC= 1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101000; // iC=  616 
vC = 14'b0000010000011100; // vC= 1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001000; // iC=  584 
vC = 14'b0000001111110101; // vC= 1013 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000110; // iC=  582 
vC = 14'b0000010000101100; // vC= 1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001110; // iC=  590 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010011; // iC=  531 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111101; // iC=  573 
vC = 14'b0000010000111000; // vC= 1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111000; // iC=  504 
vC = 14'b0000001111101011; // vC= 1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111010; // iC=  442 
vC = 14'b0000010000010100; // vC= 1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100010; // iC=  482 
vC = 14'b0000001111001111; // vC=  975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011111; // iC=  479 
vC = 14'b0000001111011110; // vC=  990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111000; // iC=  568 
vC = 14'b0000010001000111; // vC= 1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000001; // iC=  513 
vC = 14'b0000010000101011; // vC= 1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001100; // iC=  460 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000111; // iC=  519 
vC = 14'b0000010000100011; // vC= 1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100001; // iC=  417 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100101; // iC=  549 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101001; // iC=  489 
vC = 14'b0000001111101100; // vC= 1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110011; // iC=  499 
vC = 14'b0000010001100101; // vC= 1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001100; // iC=  396 
vC = 14'b0000010001000000; // vC= 1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000111; // iC=  391 
vC = 14'b0000010000100000; // vC= 1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010101; // iC=  533 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010000; // iC=  400 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101110; // iC=  494 
vC = 14'b0000001111100110; // vC=  998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101101; // iC=  429 
vC = 14'b0000010000110111; // vC= 1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000001; // iC=  513 
vC = 14'b0000010000010101; // vC= 1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110001; // iC=  369 
vC = 14'b0000010000000010; // vC= 1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111100; // iC=  380 
vC = 14'b0000010001000001; // vC= 1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000110; // iC=  390 
vC = 14'b0000010000100011; // vC= 1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011100; // iC=  412 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010001; // iC=  337 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000001; // iC=  385 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000100; // iC=  452 
vC = 14'b0000001111110111; // vC= 1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001001; // iC=  329 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111110; // iC=  382 
vC = 14'b0000001111110100; // vC= 1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010001; // iC=  465 
vC = 14'b0000010001001000; // vC= 1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100011; // iC=  355 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110010; // iC=  434 
vC = 14'b0000010001000001; // vC= 1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001100; // iC=  332 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110100; // iC=  308 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001100; // iC=  396 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010111; // iC=  407 
vC = 14'b0000010001011110; // vC= 1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100010; // iC=  354 
vC = 14'b0000010010000010; // vC= 1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111010; // iC=  378 
vC = 14'b0000010000110011; // vC= 1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100101; // iC=  357 
vC = 14'b0000010001000001; // vC= 1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100100; // iC=  292 
vC = 14'b0000010001000111; // vC= 1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011000; // iC=  280 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000101; // iC=  325 
vC = 14'b0000010000000110; // vC= 1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110101; // iC=  309 
vC = 14'b0000010001101000; // vC= 1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111110; // iC=  318 
vC = 14'b0000010001110010; // vC= 1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011010; // iC=  282 
vC = 14'b0000010000010100; // vC= 1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100100; // iC=  356 
vC = 14'b0000010000100001; // vC= 1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010100; // iC=  212 
vC = 14'b0000010001110010; // vC= 1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000001; // iC=  321 
vC = 14'b0000010000101011; // vC= 1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001100; // iC=  332 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111100; // iC=  252 
vC = 14'b0000010001001110; // vC= 1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110001; // iC=  305 
vC = 14'b0000010000101010; // vC= 1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110100; // iC=  180 
vC = 14'b0000010001100101; // vC= 1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100101; // iC=  229 
vC = 14'b0000010001101001; // vC= 1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000001; // iC=  193 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010000; // iC=  208 
vC = 14'b0000010001010110; // vC= 1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010110; // iC=  150 
vC = 14'b0000010001110110; // vC= 1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000000; // iC=  192 
vC = 14'b0000010010000101; // vC= 1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101110; // iC=  174 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011101; // iC=  157 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111001; // iC=  185 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000111; // iC=  199 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000101; // iC=  197 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000110; // iC=   70 
vC = 14'b0000010010001011; // vC= 1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010111; // iC=  151 
vC = 14'b0000010001101110; // vC= 1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010011; // iC=   83 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000000; // iC=  128 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111001; // iC=   -7 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110111; // iC=   55 
vC = 14'b0000010010011011; // vC= 1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000101; // iC=    5 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011000; // iC=   88 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110100; // iC=  -76 
vC = 14'b0000010000110001; // vC= 1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000101; // iC=  -59 
vC = 14'b0000010001100011; // vC= 1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101001; // iC=   41 
vC = 14'b0000010000011001; // vC= 1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111110; // iC=  -66 
vC = 14'b0000010000001001; // vC= 1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100110; // iC=  -26 
vC = 14'b0000010001110110; // vC= 1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000110; // iC= -122 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001111; // iC= -113 
vC = 14'b0000010001111100; // vC= 1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110011; // iC= -141 
vC = 14'b0000010001110011; // vC= 1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001100; // iC= -180 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011001; // iC= -103 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101011; // iC= -213 
vC = 14'b0000010000011001; // vC= 1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101000; // iC= -280 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110110; // iC= -266 
vC = 14'b0000010000100100; // vC= 1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001000; // iC= -184 
vC = 14'b0000010001111111; // vC= 1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010101; // iC= -299 
vC = 14'b0000010001111001; // vC= 1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000000; // iC= -256 
vC = 14'b0000010000111010; // vC= 1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011101; // iC= -291 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001000; // iC= -376 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111011; // iC= -325 
vC = 14'b0000010000011001; // vC= 1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111110; // iC= -386 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000010; // iC= -382 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101101; // iC= -467 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000001; // iC= -383 
vC = 14'b0000010000000101; // vC= 1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110110; // iC= -394 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101110; // iC= -530 
vC = 14'b0000010000100001; // vC= 1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010101; // iC= -555 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111010; // iC= -518 
vC = 14'b0000010000101110; // vC= 1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001010; // iC= -566 
vC = 14'b0000001111100010; // vC=  994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000000; // iC= -512 
vC = 14'b0000001111001111; // vC=  975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100010; // iC= -542 
vC = 14'b0000001111111111; // vC= 1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110100; // iC= -588 
vC = 14'b0000010000000001; // vC= 1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000101; // iC= -635 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001010; // iC= -630 
vC = 14'b0000010000101111; // vC= 1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011101; // iC= -675 
vC = 14'b0000010000001000; // vC= 1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001001; // iC= -631 
vC = 14'b0000010000110101; // vC= 1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111111; // iC= -705 
vC = 14'b0000001110111110; // vC=  958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110101; // iC= -715 
vC = 14'b0000010001010011; // vC= 1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000111; // iC= -825 
vC = 14'b0000001110110101; // vC=  949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001100; // iC= -756 
vC = 14'b0000001111000110; // vC=  966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011011; // iC= -741 
vC = 14'b0000001110111001; // vC=  953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001110; // iC= -818 
vC = 14'b0000001111001111; // vC=  975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010011; // iC= -813 
vC = 14'b0000001110110000; // vC=  944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001100; // iC= -884 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101111; // iC= -849 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101010; // iC= -854 
vC = 14'b0000001111010111; // vC=  983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001000; // iC= -888 
vC = 14'b0000010000001101; // vC= 1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110110; // iC= -906 
vC = 14'b0000001110010110; // vC=  918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111101; // iC= -899 
vC = 14'b0000001111000000; // vC=  960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111001; // iC=-1031 
vC = 14'b0000001110001100; // vC=  908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100000; // iC= -992 
vC = 14'b0000010000000000; // vC= 1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101011; // iC=-1045 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111101; // iC=-1027 
vC = 14'b0000001101111101; // vC=  893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110001; // iC=-1103 
vC = 14'b0000010000000000; // vC= 1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000001; // iC=-1087 
vC = 14'b0000001111001110; // vC=  974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101100; // iC= -980 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001111; // iC=-1137 
vC = 14'b0000001101101101; // vC=  877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011110; // iC=-1122 
vC = 14'b0000001110101110; // vC=  942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011000; // iC=-1064 
vC = 14'b0000001101111001; // vC=  889 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100101; // iC=-1051 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010101; // iC=-1131 
vC = 14'b0000001110001000; // vC=  904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111111; // iC=-1089 
vC = 14'b0000001110011101; // vC=  925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110010; // iC=-1102 
vC = 14'b0000001111011010; // vC=  986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110101; // iC=-1099 
vC = 14'b0000001110101010; // vC=  938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100110; // iC=-1178 
vC = 14'b0000001110101111; // vC=  943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010100; // iC=-1196 
vC = 14'b0000001110011000; // vC=  920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b0000001101011101; // vC=  861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111001; // iC=-1287 
vC = 14'b0000001110000010; // vC=  898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111000; // iC=-1224 
vC = 14'b0000001110101000; // vC=  936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001011; // iC=-1205 
vC = 14'b0000001110100100; // vC=  932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110000; // iC=-1296 
vC = 14'b0000001111001110; // vC=  974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000100; // iC=-1340 
vC = 14'b0000001110001010; // vC=  906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111101; // iC=-1347 
vC = 14'b0000001100101010; // vC=  810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101011; // iC=-1301 
vC = 14'b0000001101011010; // vC=  858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010111; // iC=-1257 
vC = 14'b0000001110110001; // vC=  945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111010; // iC=-1286 
vC = 14'b0000001110011001; // vC=  921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100010; // iC=-1310 
vC = 14'b0000001100110101; // vC=  821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100110; // iC=-1370 
vC = 14'b0000001100110110; // vC=  822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101011; // iC=-1429 
vC = 14'b0000001100110010; // vC=  818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011110; // iC=-1378 
vC = 14'b0000001100000110; // vC=  774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001011; // iC=-1397 
vC = 14'b0000001101110100; // vC=  884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110011; // iC=-1421 
vC = 14'b0000001011110111; // vC=  759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b0000001100001011; // vC=  779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b0000001101110001; // vC=  881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b0000001101000000; // vC=  832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010010; // iC=-1390 
vC = 14'b0000001011100010; // vC=  738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b0000001101101100; // vC=  876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101110; // iC=-1362 
vC = 14'b0000001101010010; // vC=  850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010011; // iC=-1517 
vC = 14'b0000001100011101; // vC=  797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001010; // iC=-1526 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111101; // iC=-1411 
vC = 14'b0000001101011010; // vC=  858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b0000001011001111; // vC=  719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b0000001011000111; // vC=  711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111111; // iC=-1409 
vC = 14'b0000001100010101; // vC=  789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010101; // iC=-1451 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b0000001100001011; // vC=  779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100110; // iC=-1434 
vC = 14'b0000001100011101; // vC=  797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b0000001010010101; // vC=  661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000001010011110; // vC=  670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b0000001010011010; // vC=  666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b0000001011111001; // vC=  761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011001; // iC=-1447 
vC = 14'b0000001010100111; // vC=  679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000011; // iC=-1469 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b0000001010001000; // vC=  648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011000; // iC=-1512 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b0000001011000110; // vC=  710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b0000001011001001; // vC=  713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b0000001001101101; // vC=  621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b0000001001001100; // vC=  588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b0000001001100101; // vC=  613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b0000001010011011; // vC=  667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111010; // iC=-1478 
vC = 14'b0000001001101110; // vC=  622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101101; // iC=-1555 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b0000001001100110; // vC=  614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001000; // iC=-1464 
vC = 14'b0000001001000000; // vC=  576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b0000001000100011; // vC=  547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b0000001010001110; // vC=  654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110111; // iC=-1609 
vC = 14'b0000001010000101; // vC=  645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b0000001001111101; // vC=  637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b0000001000111011; // vC=  571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b0000001001011010; // vC=  602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b0000001001011001; // vC=  601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100111; // iC=-1497 
vC = 14'b0000001000111111; // vC=  575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b0000001000010101; // vC=  533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010100; // iC=-1580 
vC = 14'b0000001000000100; // vC=  516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010000; // iC=-1456 
vC = 14'b0000001001010001; // vC=  593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111001; // iC=-1479 
vC = 14'b0000001001111010; // vC=  634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000001000111001; // vC=  569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000010; // iC=-1470 
vC = 14'b0000000111110101; // vC=  501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101100; // iC=-1556 
vC = 14'b0000001001101110; // vC=  622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b0000000111100110; // vC=  486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000001001010101; // vC=  597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b0000001000100001; // vC=  545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100111; // iC=-1497 
vC = 14'b0000001000100010; // vC=  546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b0000001001010010; // vC=  594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001111; // iC=-1457 
vC = 14'b0000001000000110; // vC=  518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b0000000111010010; // vC=  466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b0000001000101100; // vC=  556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101100; // iC=-1556 
vC = 14'b0000000110101001; // vC=  425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b0000000110010110; // vC=  406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000001000001111; // vC=  527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b0000000110110000; // vC=  432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110111; // iC=-1545 
vC = 14'b0000001000000011; // vC=  515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110000; // iC=-1552 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b0000001000000110; // vC=  518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b0000000101110010; // vC=  370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000000110111011; // vC=  443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b0000000101100111; // vC=  359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000011; // iC=-1469 
vC = 14'b0000000111100010; // vC=  482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b0000000101001011; // vC=  331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000000101100101; // vC=  357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b0000000111010101; // vC=  469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011110; // iC=-1442 
vC = 14'b0000000111010001; // vC=  465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001100; // iC=-1588 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b0000000101010110; // vC=  342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b0000000101000110; // vC=  326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b0000000101111110; // vC=  382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000000110100100; // vC=  420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b0000000100111110; // vC=  318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000000100101001; // vC=  297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b0000000101001111; // vC=  335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b0000000100010011; // vC=  275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b0000000101101010; // vC=  362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110101; // iC=-1483 
vC = 14'b0000000011111111; // vC=  255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b0000000101000110; // vC=  326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b0000000101011110; // vC=  350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b0000000101000011; // vC=  323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111111; // iC=-1537 
vC = 14'b0000000011100011; // vC=  227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010100; // iC=-1580 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b0000000011100010; // vC=  226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b0000000011111100; // vC=  252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b0000000101001000; // vC=  328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b0000000101000001; // vC=  321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b0000000010111001; // vC=  185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000000101010000; // vC=  336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101111; // iC=-1553 
vC = 14'b0000000011000101; // vC=  197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100011; // iC=-1501 
vC = 14'b0000000011100100; // vC=  228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b0000000011100000; // vC=  224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b0000000011100100; // vC=  228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101011; // iC=-1557 
vC = 14'b0000000100000100; // vC=  260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000011; // iC=-1405 
vC = 14'b0000000011000110; // vC=  198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001000; // iC=-1464 
vC = 14'b0000000011110001; // vC=  241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001100; // iC=-1524 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110000; // iC=-1488 
vC = 14'b0000000100001101; // vC=  269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b0000000010000001; // vC=  129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001111; // iC=-1457 
vC = 14'b0000000001110100; // vC=  116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111111; // iC=-1537 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b0000000001101000; // vC=  104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b0000000001101001; // vC=  105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110101; // iC=-1483 
vC = 14'b0000000011011011; // vC=  219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b0000000010100101; // vC=  165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111011; // iC=-1413 
vC = 14'b0000000011001001; // vC=  201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000010; // iC=-1470 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001011; // iC=-1397 
vC = 14'b0000000001101010; // vC=  106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000011; // iC=-1405 
vC = 14'b0000000010011011; // vC=  155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110100; // iC=-1420 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b0000000010011100; // vC=  156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b0000000010001010; // vC=  138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000000001010111; // vC=   87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001100; // iC=-1396 
vC = 14'b0000000000110001; // vC=   49 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b0000000001100101; // vC=  101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b0000000010000101; // vC=  133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110101; // iC=-1483 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100010; // iC=-1502 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111001; // iC=-1351 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110000; // iC=-1488 
vC = 14'b0000000001110111; // vC=  119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b0000000001000111; // vC=   71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100011; // iC=-1373 
vC = 14'b1111111111011010; // vC=  -38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b0000000000100100; // vC=   36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b1111111111110010; // vC=  -14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b0000000001011101; // vC=   93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000100; // iC=-1404 
vC = 14'b1111111111001101; // vC=  -51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001011; // iC=-1333 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010010; // iC=-1454 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110011; // iC=-1357 
vC = 14'b1111111111011001; // vC=  -39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110011; // iC=-1357 
vC = 14'b1111111111110100; // vC=  -12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000110; // iC=-1402 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000110; // iC=-1402 
vC = 14'b1111111110101010; // vC=  -86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b1111111111001010; // vC=  -54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001101; // iC=-1331 
vC = 14'b1111111111011101; // vC=  -35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111111; // iC=-1409 
vC = 14'b1111111111000111; // vC=  -57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b1111111110010110; // vC= -106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011101; // iC=-1443 
vC = 14'b1111111110111110; // vC=  -66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b1111111110001010; // vC= -118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111111110100000; // vC=  -96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011110; // iC=-1378 
vC = 14'b1111111111010010; // vC=  -46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000001; // iC=-1407 
vC = 14'b0000000000001000; // vC=    8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011011; // iC=-1317 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010111; // iC=-1321 
vC = 14'b1111111110011010; // vC= -102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010000; // iC=-1328 
vC = 14'b0000000000000011; // vC=    3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010100; // iC=-1388 
vC = 14'b1111111110000011; // vC= -125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100101; // iC=-1371 
vC = 14'b1111111111110110; // vC=  -10 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011111; // iC=-1313 
vC = 14'b1111111101101100; // vC= -148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111111111011001; // vC=  -39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101010; // iC=-1366 
vC = 14'b1111111110101001; // vC=  -87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b1111111110111011; // vC=  -69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011000; // iC=-1320 
vC = 14'b1111111101111101; // vC= -131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101001; // iC=-1303 
vC = 14'b1111111110001011; // vC= -117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b1111111101000011; // vC= -189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111101; // iC=-1411 
vC = 14'b1111111100111111; // vC= -193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111000; // iC=-1352 
vC = 14'b1111111110001000; // vC= -120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000000; // iC=-1280 
vC = 14'b1111111110110110; // vC=  -74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010110; // iC=-1386 
vC = 14'b1111111101000010; // vC= -190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111010; // iC=-1286 
vC = 14'b1111111110111100; // vC=  -68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001101; // iC=-1267 
vC = 14'b1111111110001000; // vC= -120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000110; // iC=-1402 
vC = 14'b1111111101010100; // vC= -172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011000; // iC=-1384 
vC = 14'b1111111100110000; // vC= -208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001001; // iC=-1399 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111000; // iC=-1352 
vC = 14'b1111111101011110; // vC= -162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010110; // iC=-1386 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b1111111101011011; // vC= -165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110110; // iC=-1290 
vC = 14'b1111111100110101; // vC= -203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010111; // iC=-1257 
vC = 14'b1111111101001100; // vC= -180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111100; // iC=-1348 
vC = 14'b1111111110001100; // vC= -116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010111; // iC=-1257 
vC = 14'b1111111101000000; // vC= -192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011100; // iC=-1252 
vC = 14'b1111111100010100; // vC= -236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100010; // iC=-1246 
vC = 14'b1111111011110011; // vC= -269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110100; // iC=-1356 
vC = 14'b1111111101110001; // vC= -143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011011; // iC=-1253 
vC = 14'b1111111100011110; // vC= -226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010011; // iC=-1325 
vC = 14'b1111111100100000; // vC= -224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101011; // iC=-1365 
vC = 14'b1111111100010110; // vC= -234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000001; // iC=-1215 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011001; // iC=-1255 
vC = 14'b1111111011010101; // vC= -299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101011; // iC=-1301 
vC = 14'b1111111100101100; // vC= -212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100111; // iC=-1241 
vC = 14'b1111111010110111; // vC= -329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111111; // iC=-1281 
vC = 14'b1111111011101010; // vC= -278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010100; // iC=-1324 
vC = 14'b1111111100101000; // vC= -216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010110; // iC=-1258 
vC = 14'b1111111100011100; // vC= -228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011011; // iC=-1317 
vC = 14'b1111111011001101; // vC= -307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101011; // iC=-1237 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b1111111010100000; // vC= -352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010101; // iC=-1259 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b1111111011010101; // vC= -299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011001; // iC=-1319 
vC = 14'b1111111100011111; // vC= -225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b1111111100001100; // vC= -244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111000; // iC=-1224 
vC = 14'b1111111010010001; // vC= -367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110100; // iC=-1228 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101011; // iC=-1237 
vC = 14'b1111111011110011; // vC= -269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101001; // iC=-1239 
vC = 14'b1111111100000111; // vC= -249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011101; // iC=-1251 
vC = 14'b1111111011010010; // vC= -302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011011; // iC=-1253 
vC = 14'b1111111001101111; // vC= -401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110000; // iC=-1168 
vC = 14'b1111111011001100; // vC= -308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b1111111010100111; // vC= -345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100100; // iC=-1244 
vC = 14'b1111111001101011; // vC= -405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101111; // iC=-1233 
vC = 14'b1111111001101101; // vC= -403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001110; // iC=-1202 
vC = 14'b1111111010101000; // vC= -344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b1111111010000011; // vC= -381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110010; // iC=-1166 
vC = 14'b1111111011001110; // vC= -306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100110; // iC=-1242 
vC = 14'b1111111010111100; // vC= -324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011011; // iC=-1253 
vC = 14'b1111111011100000; // vC= -288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110111; // iC=-1161 
vC = 14'b1111111001111101; // vC= -387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111010; // iC=-1286 
vC = 14'b1111111001011101; // vC= -419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000101; // iC=-1147 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101110; // iC=-1170 
vC = 14'b1111111001010001; // vC= -431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001010; // iC=-1270 
vC = 14'b1111111010010100; // vC= -364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101111; // iC=-1233 
vC = 14'b1111111001011010; // vC= -422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001001; // iC=-1207 
vC = 14'b1111111010011001; // vC= -359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101100; // iC=-1108 
vC = 14'b1111111001011001; // vC= -423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001011; // iC=-1141 
vC = 14'b1111111000110101; // vC= -459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010110; // iC=-1258 
vC = 14'b1111111010011111; // vC= -353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000001; // iC=-1215 
vC = 14'b1111111001100100; // vC= -412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011100; // iC=-1188 
vC = 14'b1111111010011011; // vC= -357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110111; // iC=-1161 
vC = 14'b1111111010010111; // vC= -361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111111; // iC=-1089 
vC = 14'b1111111001110110; // vC= -394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011111; // iC=-1185 
vC = 14'b1111111010011001; // vC= -359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010010; // iC=-1198 
vC = 14'b1111111000110011; // vC= -461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001110; // iC=-1138 
vC = 14'b1111111010010101; // vC= -363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011011; // iC=-1125 
vC = 14'b1111111001100101; // vC= -411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001001; // iC=-1079 
vC = 14'b1111111000011000; // vC= -488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b1111111001111110; // vC= -386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010100; // iC=-1132 
vC = 14'b1111110111111100; // vC= -516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001110; // iC=-1074 
vC = 14'b1111110111100011; // vC= -541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100010; // iC=-1118 
vC = 14'b1111110111101111; // vC= -529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011101; // iC=-1059 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011101; // iC=-1123 
vC = 14'b1111111001001000; // vC= -440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111100; // iC=-1092 
vC = 14'b1111111001000011; // vC= -445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110110; // iC=-1098 
vC = 14'b1111110111101111; // vC= -529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110101; // iC=-1099 
vC = 14'b1111110111011001; // vC= -551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101010; // iC=-1174 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010110; // iC=-1066 
vC = 14'b1111110111000111; // vC= -569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110101; // iC=-1035 
vC = 14'b1111110111100011; // vC= -541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100101; // iC=-1115 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110011; // iC=-1101 
vC = 14'b1111111001000101; // vC= -443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010000; // iC=-1072 
vC = 14'b1111111000010011; // vC= -493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000111; // iC=-1081 
vC = 14'b1111110111101110; // vC= -530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101001; // iC=-1111 
vC = 14'b1111111000000000; // vC= -512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110000; // iC=-1104 
vC = 14'b1111110111100100; // vC= -540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000001; // iC=-1023 
vC = 14'b1111111000010101; // vC= -491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101100; // iC=-1108 
vC = 14'b1111110110100100; // vC= -604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011000; // iC=-1128 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010000; // iC=-1136 
vC = 14'b1111110111110000; // vC= -528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011011; // iC=-1061 
vC = 14'b1111110110110011; // vC= -589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111111; // iC=-1089 
vC = 14'b1111110111100011; // vC= -541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010011; // iC=-1005 
vC = 14'b1111110111010010; // vC= -558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001110; // iC=-1010 
vC = 14'b1111110111111010; // vC= -518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100101; // iC=-1115 
vC = 14'b1111111000010000; // vC= -496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001000; // iC=-1016 
vC = 14'b1111110110011111; // vC= -609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111101; // iC=-1027 
vC = 14'b1111110111100100; // vC= -540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011111; // iC= -993 
vC = 14'b1111111000001000; // vC= -504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100010; // iC=-1054 
vC = 14'b1111110110001001; // vC= -631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110100; // iC=-1036 
vC = 14'b1111110111010001; // vC= -559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110011; // iC=-1037 
vC = 14'b1111110110111111; // vC= -577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110101; // iC=-1035 
vC = 14'b1111110111010110; // vC= -554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110011; // iC= -973 
vC = 14'b1111110110000010; // vC= -638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001000; // iC=-1016 
vC = 14'b1111110110010011; // vC= -621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010010; // iC= -942 
vC = 14'b1111110110110101; // vC= -587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101100; // iC=-1044 
vC = 14'b1111110110011100; // vC= -612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101111; // iC= -977 
vC = 14'b1111110101100010; // vC= -670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011000; // iC=-1064 
vC = 14'b1111110110000011; // vC= -637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011000; // iC= -936 
vC = 14'b1111110111000110; // vC= -570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111011; // iC=-1029 
vC = 14'b1111110110001011; // vC= -629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100101; // iC=-1051 
vC = 14'b1111110110100110; // vC= -602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101011; // iC= -981 
vC = 14'b1111110110010101; // vC= -619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001101; // iC= -947 
vC = 14'b1111110101100010; // vC= -670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100111; // iC=-1049 
vC = 14'b1111110101011110; // vC= -674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101110; // iC=-1042 
vC = 14'b1111110100111010; // vC= -710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011001; // iC= -935 
vC = 14'b1111110101101111; // vC= -657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010111; // iC=-1001 
vC = 14'b1111110101100001; // vC= -671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101101; // iC= -915 
vC = 14'b1111110100101111; // vC= -721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111010; // iC=-1030 
vC = 14'b1111110100111010; // vC= -710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101110; // iC= -914 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100011; // iC= -925 
vC = 14'b1111110100110100; // vC= -716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010100; // iC= -940 
vC = 14'b1111110110111000; // vC= -584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001111; // iC=-1009 
vC = 14'b1111110110110010; // vC= -590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101111; // iC= -977 
vC = 14'b1111110101001110; // vC= -690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001011; // iC= -949 
vC = 14'b1111110110011001; // vC= -615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110110; // iC= -906 
vC = 14'b1111110110010000; // vC= -624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111101; // iC= -963 
vC = 14'b1111110101010101; // vC= -683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101010; // iC= -854 
vC = 14'b1111110100101111; // vC= -721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011001; // iC= -871 
vC = 14'b1111110110011000; // vC= -616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111000; // iC= -904 
vC = 14'b1111110100110011; // vC= -717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100100; // iC= -924 
vC = 14'b1111110100000011; // vC= -765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010101; // iC= -939 
vC = 14'b1111110101001101; // vC= -691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110101; // iC= -907 
vC = 14'b1111110101010101; // vC= -683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111000; // iC= -968 
vC = 14'b1111110110000000; // vC= -640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110011; // iC= -845 
vC = 14'b1111110100100000; // vC= -736 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011110; // iC= -866 
vC = 14'b1111110101001000; // vC= -696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010111; // iC= -809 
vC = 14'b1111110011110101; // vC= -779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100011; // iC= -861 
vC = 14'b1111110100001001; // vC= -759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101000; // iC= -920 
vC = 14'b1111110100001000; // vC= -760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010011; // iC= -941 
vC = 14'b1111110100100010; // vC= -734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111111; // iC= -833 
vC = 14'b1111110101111001; // vC= -647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011001; // iC= -871 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001011; // iC= -885 
vC = 14'b1111110100101000; // vC= -728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011111; // iC= -929 
vC = 14'b1111110101101110; // vC= -658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011001; // iC= -807 
vC = 14'b1111110101001111; // vC= -689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000011; // iC= -829 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100110; // iC= -858 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110001; // iC= -911 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110000; // iC= -912 
vC = 14'b1111110100001011; // vC= -757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101010; // iC= -854 
vC = 14'b1111110100011011; // vC= -741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111010; // iC= -838 
vC = 14'b1111110100011101; // vC= -739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110110; // iC= -778 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110111; // iC= -841 
vC = 14'b1111110100001001; // vC= -759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100101; // iC= -859 
vC = 14'b1111110101001100; // vC= -692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110110; // iC= -778 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010101; // iC= -747 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100100; // iC= -796 
vC = 14'b1111110010111100; // vC= -836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101111; // iC= -849 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011101; // iC= -803 
vC = 14'b1111110100010000; // vC= -752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101110; // iC= -850 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011111; // iC= -737 
vC = 14'b1111110100010100; // vC= -748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101101; // iC= -787 
vC = 14'b1111110010011111; // vC= -865 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000000; // iC= -832 
vC = 14'b1111110100011110; // vC= -738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111111; // iC= -769 
vC = 14'b1111110011000101; // vC= -827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011100; // iC= -740 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001001; // iC= -759 
vC = 14'b1111110011000000; // vC= -832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010100; // iC= -684 
vC = 14'b1111110100101000; // vC= -728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010001; // iC= -687 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011111; // iC= -737 
vC = 14'b1111110100100100; // vC= -732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100111; // iC= -729 
vC = 14'b1111110011001101; // vC= -819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011111; // iC= -737 
vC = 14'b1111110011101011; // vC= -789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001010; // iC= -758 
vC = 14'b1111110011101100; // vC= -788 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101010; // iC= -726 
vC = 14'b1111110011010011; // vC= -813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110100; // iC= -780 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111001; // iC= -775 
vC = 14'b1111110010010101; // vC= -875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100011; // iC= -669 
vC = 14'b1111110001110110; // vC= -906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110010; // iC= -654 
vC = 14'b1111110011100110; // vC= -794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010110; // iC= -682 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101010; // iC= -662 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001011; // iC= -629 
vC = 14'b1111110010000001; // vC= -895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011111; // iC= -737 
vC = 14'b1111110001111110; // vC= -898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001010; // iC= -758 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000011; // iC= -701 
vC = 14'b1111110010101001; // vC= -855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000101; // iC= -699 
vC = 14'b1111110010011110; // vC= -866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010111; // iC= -681 
vC = 14'b1111110001111101; // vC= -899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110110; // iC= -650 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010010; // iC= -686 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101001; // iC= -599 
vC = 14'b1111110010110011; // vC= -845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110011; // iC= -653 
vC = 14'b1111110011011100; // vC= -804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000100; // iC= -636 
vC = 14'b1111110001110111; // vC= -905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111010; // iC= -646 
vC = 14'b1111110010010011; // vC= -877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101111; // iC= -721 
vC = 14'b1111110010001011; // vC= -885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000000; // iC= -640 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101001; // iC= -727 
vC = 14'b1111110011011111; // vC= -801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010010; // iC= -686 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000100; // iC= -572 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110100; // iC= -652 
vC = 14'b1111110010111010; // vC= -838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100100; // iC= -668 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110101; // iC= -587 
vC = 14'b1111110010100101; // vC= -859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110111; // iC= -649 
vC = 14'b1111110010110101; // vC= -843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100101; // iC= -539 
vC = 14'b1111110011010011; // vC= -813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100011; // iC= -541 
vC = 14'b1111110001000010; // vC= -958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011011; // iC= -549 
vC = 14'b1111110010110011; // vC= -845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101101; // iC= -595 
vC = 14'b1111110011000101; // vC= -827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011010; // iC= -614 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100001; // iC= -607 
vC = 14'b1111110001100110; // vC= -922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101010; // iC= -662 
vC = 14'b1111110010101000; // vC= -856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101111; // iC= -529 
vC = 14'b1111110010000011; // vC= -893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011100; // iC= -548 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011101; // iC= -547 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111010; // iC= -582 
vC = 14'b1111110001000000; // vC= -960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000011; // iC= -509 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011010; // iC= -486 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011001; // iC= -487 
vC = 14'b1111110010110101; // vC= -843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111001; // iC= -519 
vC = 14'b1111110001001111; // vC= -945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110010; // iC= -526 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010110; // iC= -554 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001010; // iC= -502 
vC = 14'b1111110000110001; // vC= -975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101111; // iC= -529 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011111; // iC= -545 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100111; // iC= -537 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001011; // iC= -501 
vC = 14'b1111110000101010; // vC= -982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001010; // iC= -566 
vC = 14'b1111110000001001; // vC=-1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001001; // iC= -439 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000010; // iC= -446 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010101; // iC= -555 
vC = 14'b1111110000001111; // vC=-1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011011; // iC= -421 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111110010001111; // vC= -881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100000; // iC= -416 
vC = 14'b1111110001110100; // vC= -908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110100; // iC= -524 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011100; // iC= -548 
vC = 14'b1111110000101000; // vC= -984 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101110; // iC= -530 
vC = 14'b1111110010010010; // vC= -878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111011; // iC= -453 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100010; // iC= -414 
vC = 14'b1111110000100010; // vC= -990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100111; // iC= -537 
vC = 14'b1111110010001000; // vC= -888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101011; // iC= -405 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110101; // iC= -395 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010000; // iC= -432 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001011; // iC= -501 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110001; // iC= -463 
vC = 14'b1111110001010001; // vC= -943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100100; // iC= -412 
vC = 14'b1111110000010101; // vC=-1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110000; // iC= -464 
vC = 14'b1111101111110011; // vC=-1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001110; // iC= -434 
vC = 14'b1111110001011001; // vC= -935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110010; // iC= -462 
vC = 14'b1111110001101111; // vC= -913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101001; // iC= -343 
vC = 14'b1111110000100100; // vC= -988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001101; // iC= -371 
vC = 14'b1111110000101001; // vC= -983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000010; // iC= -382 
vC = 14'b1111101111110101; // vC=-1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001100; // iC= -372 
vC = 14'b1111110000100001; // vC= -991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101110; // iC= -466 
vC = 14'b1111110001100001; // vC= -927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101110; // iC= -338 
vC = 14'b1111110001111011; // vC= -901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000000; // iC= -384 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101011; // iC= -341 
vC = 14'b1111110001101000; // vC= -920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111001; // iC= -391 
vC = 14'b1111110001110011; // vC= -909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110101; // iC= -331 
vC = 14'b1111101111100010; // vC=-1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111111; // iC= -321 
vC = 14'b1111101111100011; // vC=-1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100000; // iC= -416 
vC = 14'b1111110000100100; // vC= -988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001010; // iC= -374 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101010; // iC= -406 
vC = 14'b1111101111100001; // vC=-1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001010; // iC= -310 
vC = 14'b1111110001101111; // vC= -913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000101; // iC= -315 
vC = 14'b1111110000100010; // vC= -990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111100; // iC= -388 
vC = 14'b1111110001001110; // vC= -946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011011; // iC= -293 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011100; // iC= -292 
vC = 14'b1111110000000010; // vC=-1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010100; // iC= -364 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001110; // iC= -242 
vC = 14'b1111110000000111; // vC=-1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100000; // iC= -224 
vC = 14'b1111101111001000; // vC=-1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001011; // iC= -309 
vC = 14'b1111101111101110; // vC=-1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001101; // iC= -243 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111000; // iC= -200 
vC = 14'b1111101111001101; // vC=-1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111101; // iC= -195 
vC = 14'b1111110000100101; // vC= -987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000100; // iC= -188 
vC = 14'b1111101111010100; // vC=-1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100100; // iC= -220 
vC = 14'b1111110001001000; // vC= -952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101110; // iC= -210 
vC = 14'b1111110000010011; // vC=-1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110100; // iC= -268 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110000; // iC= -272 
vC = 14'b1111101111011000; // vC=-1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010101; // iC= -171 
vC = 14'b1111101111010111; // vC=-1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011000; // iC= -104 
vC = 14'b1111101111100000; // vC=-1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101011; // iC= -213 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101000; // iC=  -88 
vC = 14'b1111110000110110; // vC= -970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011110; // iC=  -98 
vC = 14'b1111110000010100; // vC=-1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110010; // iC=  -78 
vC = 14'b1111110000010011; // vC=-1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001101; // iC= -179 
vC = 14'b1111101111000010; // vC=-1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011100; // iC=  -36 
vC = 14'b1111110000001101; // vC=-1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001001; // iC=  -55 
vC = 14'b1111101111001000; // vC=-1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100100; // iC=  -28 
vC = 14'b1111101111100001; // vC=-1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111011; // iC=  -69 
vC = 14'b1111101111101111; // vC=-1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011000; // iC=   24 
vC = 14'b1111101111010110; // vC=-1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110101; // iC=  -75 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000111; // iC=  -57 
vC = 14'b1111110000101101; // vC= -979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000010; // iC=  -62 
vC = 14'b1111110000001101; // vC=-1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011001; // iC=  -39 
vC = 14'b1111101111111011; // vC=-1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000001; // iC=   65 
vC = 14'b1111110000110011; // vC= -973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001010; // iC=   10 
vC = 14'b1111101111011001; // vC=-1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100100; // iC=  100 
vC = 14'b1111110000001101; // vC=-1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100000; // iC=   96 
vC = 14'b1111110000000111; // vC=-1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010001; // iC=  145 
vC = 14'b1111110000010100; // vC=-1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100011; // iC=   99 
vC = 14'b1111101111100001; // vC=-1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110111; // iC=  119 
vC = 14'b1111110000100011; // vC= -989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000111; // iC=  199 
vC = 14'b1111110000011000; // vC=-1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010010; // iC=  146 
vC = 14'b1111110000011010; // vC= -998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110000; // iC=  240 
vC = 14'b1111101111110101; // vC=-1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100100; // iC=  228 
vC = 14'b1111110000100111; // vC= -985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001110; // iC=  270 
vC = 14'b1111101111011111; // vC=-1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011000; // iC=  280 
vC = 14'b1111110000101000; // vC= -984 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100001; // iC=  289 
vC = 14'b1111110000100000; // vC= -992 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011111; // iC=  351 
vC = 14'b1111101111000000; // vC=-1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111111; // iC=  383 
vC = 14'b1111101111100001; // vC=-1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010001; // iC=  337 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001001; // iC=  329 
vC = 14'b1111110000010001; // vC=-1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011110; // iC=  350 
vC = 14'b1111110001100110; // vC= -922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010010; // iC=  466 
vC = 14'b1111101111110000; // vC=-1040 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010100; // iC=  404 
vC = 14'b1111101111100100; // vC=-1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000101; // iC=  453 
vC = 14'b1111101111101010; // vC=-1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010110; // iC=  470 
vC = 14'b1111110001101010; // vC= -918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000111; // iC=  519 
vC = 14'b1111101111011000; // vC=-1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011100; // iC=  540 
vC = 14'b1111110000001111; // vC=-1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110010; // iC=  498 
vC = 14'b1111101111111001; // vC=-1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010000; // iC=  528 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100110; // iC=  614 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100000; // iC=  608 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100000; // iC=  672 
vC = 14'b1111110000111111; // vC= -961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010010; // iC=  594 
vC = 14'b1111101111111110; // vC=-1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101101; // iC=  685 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000111; // iC=  711 
vC = 14'b1111110000110110; // vC= -970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001000; // iC=  712 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101101; // iC=  685 
vC = 14'b1111101111100011; // vC=-1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011100; // iC=  668 
vC = 14'b1111110000101010; // vC= -982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111100; // iC=  764 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011001; // iC=  793 
vC = 14'b1111110001110100; // vC= -908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101000; // iC=  744 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101011; // iC=  875 
vC = 14'b1111101111111000; // vC=-1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101111; // iC=  879 
vC = 14'b1111110010000001; // vC= -895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001101; // iC=  909 
vC = 14'b1111101111110110; // vC=-1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111100; // iC=  956 
vC = 14'b1111110000101011; // vC= -981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010011; // iC=  851 
vC = 14'b1111110000110110; // vC= -970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010010; // iC=  978 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100101; // iC=  869 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101111; // iC= 1007 
vC = 14'b1111110001101111; // vC= -913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100001; // iC=  993 
vC = 14'b1111110010010111; // vC= -873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111011; // iC=  955 
vC = 14'b1111110010100000; // vC= -864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101101; // iC= 1005 
vC = 14'b1111110000111001; // vC= -967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100011; // iC= 1123 
vC = 14'b1111110010101011; // vC= -853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001010; // iC= 1034 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101001; // iC= 1129 
vC = 14'b1111110010100001; // vC= -863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110011; // iC= 1139 
vC = 14'b1111110001001110; // vC= -946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000010; // iC= 1154 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000100; // iC= 1092 
vC = 14'b1111110010101001; // vC= -855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101001; // iC= 1193 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101000; // iC= 1128 
vC = 14'b1111110001000101; // vC= -955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111011; // iC= 1211 
vC = 14'b1111110010010010; // vC= -878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100011; // iC= 1187 
vC = 14'b1111110001100000; // vC= -928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011110; // iC= 1246 
vC = 14'b1111110011000111; // vC= -825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010000; // iC= 1232 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000001; // iC= 1217 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100100; // iC= 1316 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111010; // iC= 1274 
vC = 14'b1111110010100011; // vC= -861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010101; // iC= 1365 
vC = 14'b1111110010101001; // vC= -855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010100; // iC= 1364 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101010; // iC= 1322 
vC = 14'b1111110011100010; // vC= -798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111010; // iC= 1274 
vC = 14'b1111110011100100; // vC= -796 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000100; // iC= 1284 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111111; // iC= 1343 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b1111110011101010; // vC= -790 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011100; // iC= 1372 
vC = 14'b1111110011100010; // vC= -798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110010; // iC= 1394 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110011; // iC= 1395 
vC = 14'b1111110011100111; // vC= -793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101111; // iC= 1455 
vC = 14'b1111110100100010; // vC= -734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001000; // iC= 1416 
vC = 14'b1111110010111100; // vC= -836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100110; // iC= 1446 
vC = 14'b1111110100000001; // vC= -767 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111001; // iC= 1529 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111000; // iC= 1528 
vC = 14'b1111110100010101; // vC= -747 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001101; // iC= 1485 
vC = 14'b1111110010100110; // vC= -858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110011; // iC= 1459 
vC = 14'b1111110100010110; // vC= -746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100010; // iC= 1506 
vC = 14'b1111110011000011; // vC= -829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010000; // iC= 1552 
vC = 14'b1111110100111011; // vC= -709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100010; // iC= 1506 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b1111110011000110; // vC= -826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111011; // iC= 1595 
vC = 14'b1111110011100100; // vC= -796 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b1111110011011001; // vC= -807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b1111110100011111; // vC= -737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010000; // iC= 1616 
vC = 14'b1111110100110001; // vC= -719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011001; // iC= 1561 
vC = 14'b1111110100111000; // vC= -712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b1111110101000000; // vC= -704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b1111110100111001; // vC= -711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000101; // iC= 1605 
vC = 14'b1111110100111100; // vC= -708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101111; // iC= 1711 
vC = 14'b1111110110001111; // vC= -625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101111; // iC= 1647 
vC = 14'b1111110100111000; // vC= -712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001011; // iC= 1675 
vC = 14'b1111110100101101; // vC= -723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100000; // iC= 1632 
vC = 14'b1111110110011110; // vC= -610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111101; // iC= 1597 
vC = 14'b1111110100100001; // vC= -735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b1111110100100110; // vC= -730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b1111110110010000; // vC= -624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001111; // iC= 1679 
vC = 14'b1111110110111011; // vC= -581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100010; // iC= 1698 
vC = 14'b1111110100101010; // vC= -726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110100; // iC= 1652 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b1111110100110111; // vC= -713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b1111110101011001; // vC= -679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111011; // iC= 1659 
vC = 14'b1111110101011000; // vC= -680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101010; // iC= 1642 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b1111110110100000; // vC= -608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b1111110101001100; // vC= -692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010110; // iC= 1686 
vC = 14'b1111110111101010; // vC= -534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b1111110101010111; // vC= -681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011011; // iC= 1755 
vC = 14'b1111110110111100; // vC= -580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100011; // iC= 1763 
vC = 14'b1111110111101110; // vC= -530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b1111111000000001; // vC= -511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b1111110110001001; // vC= -631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011111; // iC= 1695 
vC = 14'b1111110110000100; // vC= -636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110101; // iC= 1781 
vC = 14'b1111110111110100; // vC= -524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010010; // iC= 1682 
vC = 14'b1111110111111100; // vC= -516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b1111111000010101; // vC= -491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001010; // iC= 1738 
vC = 14'b1111110111011100; // vC= -548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001110; // iC= 1742 
vC = 14'b1111111000000110; // vC= -506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000100; // iC= 1668 
vC = 14'b1111110111110110; // vC= -522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b1111110111010111; // vC= -553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b1111110111000000; // vC= -576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100110; // iC= 1766 
vC = 14'b1111110111000111; // vC= -569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b1111110111100100; // vC= -540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010101; // iC= 1685 
vC = 14'b1111110111111100; // vC= -516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b1111111000101000; // vC= -472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b1111111000111111; // vC= -449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b1111110111101101; // vC= -531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b1111111000010101; // vC= -491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b1111111001001000; // vC= -440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b1111111001000111; // vC= -441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000111; // iC= 1671 
vC = 14'b1111111001011110; // vC= -418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b1111111000110001; // vC= -463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111001; // iC= 1785 
vC = 14'b1111111000010111; // vC= -489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b1111111000010111; // vC= -489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010010; // iC= 1682 
vC = 14'b1111111001000110; // vC= -442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100010; // iC= 1826 
vC = 14'b1111111000110001; // vC= -463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b1111111001110111; // vC= -393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111110; // iC= 1790 
vC = 14'b1111111001101111; // vC= -401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111111011001000; // vC= -312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000101; // iC= 1797 
vC = 14'b1111111001010011; // vC= -429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b1111111011000001; // vC= -319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110000; // iC= 1776 
vC = 14'b1111111011001110; // vC= -306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100111; // iC= 1703 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000100; // iC= 1796 
vC = 14'b1111111001110001; // vC= -399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b1111111001011101; // vC= -419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000110; // iC= 1734 
vC = 14'b1111111011010111; // vC= -297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111010; // iC= 1658 
vC = 14'b1111111011111101; // vC= -259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111111011111001; // vC= -263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b1111111011000010; // vC= -318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000001; // iC= 1729 
vC = 14'b1111111011101101; // vC= -275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111101; // iC= 1789 
vC = 14'b1111111011001100; // vC= -308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111111; // iC= 1663 
vC = 14'b1111111100001100; // vC= -244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111111011101111; // vC= -273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001011; // iC= 1675 
vC = 14'b1111111011111001; // vC= -263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b1111111011011000; // vC= -296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001001; // iC= 1737 
vC = 14'b1111111100010110; // vC= -234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000000; // iC= 1792 
vC = 14'b1111111011111101; // vC= -259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b1111111100000111; // vC= -249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b1111111100101100; // vC= -212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b1111111101010100; // vC= -172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101000; // iC= 1640 
vC = 14'b1111111101011001; // vC= -167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b1111111100101011; // vC= -213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b1111111011011011; // vC= -293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001110; // iC= 1742 
vC = 14'b1111111100001110; // vC= -242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b1111111100111010; // vC= -198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000100; // iC= 1732 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b1111111011101010; // vC= -278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b1111111100101110; // vC= -210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b1111111101101000; // vC= -152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b1111111100100100; // vC= -220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b1111111100011010; // vC= -230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110100; // iC= 1780 
vC = 14'b1111111101000001; // vC= -191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b1111111101011001; // vC= -167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111111101101011; // vC= -149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010101; // iC= 1749 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b1111111100011010; // vC= -230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b1111111110111001; // vC=  -71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101110; // iC= 1646 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100110; // iC= 1766 
vC = 14'b1111111110011011; // vC= -101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b1111111101011000; // vC= -168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b1111111101111000; // vC= -136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b1111111101100001; // vC= -159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b1111111110010101; // vC= -107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000100; // iC= 1732 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b1111111101001100; // vC= -180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010100; // iC= 1620 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101100; // iC= 1644 
vC = 14'b1111111111011001; // vC=  -39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b1111111111001110; // vC=  -50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b1111111110101010; // vC=  -86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101000; // iC= 1640 
vC = 14'b1111111111010110; // vC=  -42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b1111111111001101; // vC=  -51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010011; // iC= 1619 
vC = 14'b1111111111110011; // vC=  -13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111111; // iC= 1599 
vC = 14'b1111111101111111; // vC= -129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b1111111111100000; // vC=  -32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b0000000000011111; // vC=   31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100010; // iC= 1634 
vC = 14'b0000000000000010; // vC=    2 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b1111111111010011; // vC=  -45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b1111111111010111; // vC=  -41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b1111111110100001; // vC=  -95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b0000000000100000; // vC=   32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010101; // iC= 1685 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000010; // iC= 1730 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001101; // iC= 1677 
vC = 14'b1111111111100000; // vC=  -32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101010; // iC= 1642 
vC = 14'b0000000000101111; // vC=   47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001000; // iC= 1672 
vC = 14'b1111111111010110; // vC=  -42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000110; // iC= 1670 
vC = 14'b0000000001100000; // vC=   96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110011; // iC= 1651 
vC = 14'b0000000000111000; // vC=   56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011110; // iC= 1566 
vC = 14'b1111111111111000; // vC=   -8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011101; // iC= 1693 
vC = 14'b1111111111110100; // vC=  -12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101110; // iC= 1582 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001110; // iC= 1678 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101101; // iC= 1581 
vC = 14'b0000000010101111; // vC=  175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110010; // iC= 1650 
vC = 14'b0000000010110010; // vC=  178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000111; // iC= 1607 
vC = 14'b0000000010111001; // vC=  185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101111; // iC= 1647 
vC = 14'b0000000010111100; // vC=  188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001101; // iC= 1549 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b0000000001110101; // vC=  117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100110; // iC= 1638 
vC = 14'b0000000001101000; // vC=  104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110111; // iC= 1591 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001100; // iC= 1676 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101001; // iC= 1577 
vC = 14'b0000000011001100; // vC=  204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111011; // iC= 1595 
vC = 14'b0000000001101111; // vC=  111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111010; // iC= 1594 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b0000000001111101; // vC=  125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100100; // iC= 1572 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110000; // iC= 1584 
vC = 14'b0000000001101101; // vC=  109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001111; // iC= 1551 
vC = 14'b0000000011101111; // vC=  239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111110; // iC= 1534 
vC = 14'b0000000100000001; // vC=  257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010011; // iC= 1619 
vC = 14'b0000000100000011; // vC=  259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101011; // iC= 1579 
vC = 14'b0000000011100010; // vC=  226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010100; // iC= 1556 
vC = 14'b0000000011100001; // vC=  225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b0000000010100100; // vC=  164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b0000000010111100; // vC=  188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101100; // iC= 1644 
vC = 14'b0000000010001001; // vC=  137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100010; // iC= 1634 
vC = 14'b0000000011000011; // vC=  195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b0000000100101110; // vC=  302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010001; // iC= 1489 
vC = 14'b0000000100101001; // vC=  297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101001; // iC= 1513 
vC = 14'b0000000100101010; // vC=  298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010111; // iC= 1495 
vC = 14'b0000000011100110; // vC=  230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001001; // iC= 1609 
vC = 14'b0000000011110101; // vC=  245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001001; // iC= 1481 
vC = 14'b0000000011111101; // vC=  253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b0000000100010111; // vC=  279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010110; // iC= 1494 
vC = 14'b0000000011010111; // vC=  215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100110; // iC= 1510 
vC = 14'b0000000011110101; // vC=  245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010111; // iC= 1623 
vC = 14'b0000000100110101; // vC=  309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110110; // iC= 1462 
vC = 14'b0000000101001101; // vC=  333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100101; // iC= 1509 
vC = 14'b0000000100011100; // vC=  284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011111; // iC= 1503 
vC = 14'b0000000101011001; // vC=  345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001110; // iC= 1614 
vC = 14'b0000000101101111; // vC=  367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111001; // iC= 1529 
vC = 14'b0000000100001110; // vC=  270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001010; // iC= 1482 
vC = 14'b0000000101101100; // vC=  364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111010; // iC= 1594 
vC = 14'b0000000101010110; // vC=  342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001100; // iC= 1548 
vC = 14'b0000000101001000; // vC=  328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101001; // iC= 1513 
vC = 14'b0000000100100101; // vC=  293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b0000000110001001; // vC=  393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b0000000101110110; // vC=  374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001100; // iC= 1548 
vC = 14'b0000000101111100; // vC=  380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100111; // iC= 1511 
vC = 14'b0000000110000000; // vC=  384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001100; // iC= 1548 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001100; // iC= 1484 
vC = 14'b0000000100011111; // vC=  287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011110; // iC= 1438 
vC = 14'b0000000110011001; // vC=  409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000110; // iC= 1542 
vC = 14'b0000000100011010; // vC=  282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010011; // iC= 1555 
vC = 14'b0000000101100000; // vC=  352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101111; // iC= 1455 
vC = 14'b0000000110111111; // vC=  447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101100; // iC= 1516 
vC = 14'b0000000110100010; // vC=  418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001001; // iC= 1417 
vC = 14'b0000000110011001; // vC=  409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010000; // iC= 1424 
vC = 14'b0000000101110100; // vC=  372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111111; // iC= 1471 
vC = 14'b0000000110000010; // vC=  386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100011; // iC= 1443 
vC = 14'b0000000101100000; // vC=  352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b0000000101100001; // vC=  353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110000; // iC= 1520 
vC = 14'b0000000111000010; // vC=  450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110010; // iC= 1522 
vC = 14'b0000000101101110; // vC=  366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100110; // iC= 1510 
vC = 14'b0000000101111011; // vC=  379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000110; // iC= 1478 
vC = 14'b0000000111001100; // vC=  460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111011; // iC= 1467 
vC = 14'b0000000111011001; // vC=  473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b0000000111001001; // vC=  457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100111; // iC= 1447 
vC = 14'b0000000110101001; // vC=  425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011000; // iC= 1432 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101111; // iC= 1455 
vC = 14'b0000000110100110; // vC=  422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101110; // iC= 1518 
vC = 14'b0000000110110001; // vC=  433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010010; // iC= 1490 
vC = 14'b0000000110101110; // vC=  430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000011; // iC= 1411 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100110; // iC= 1510 
vC = 14'b0000001000000100; // vC=  516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011110; // iC= 1502 
vC = 14'b0000000110101110; // vC=  430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010111; // iC= 1431 
vC = 14'b0000000111110010; // vC=  498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110110; // iC= 1462 
vC = 14'b0000001000001101; // vC=  525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100010; // iC= 1378 
vC = 14'b0000000111101010; // vC=  490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010010; // iC= 1362 
vC = 14'b0000000111100011; // vC=  483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011000; // iC= 1496 
vC = 14'b0000000111000101; // vC=  453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100010; // iC= 1442 
vC = 14'b0000000110111010; // vC=  442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000010; // iC= 1346 
vC = 14'b0000000111100001; // vC=  481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010100; // iC= 1428 
vC = 14'b0000001000100011; // vC=  547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110000; // iC= 1328 
vC = 14'b0000000111110010; // vC=  498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110100; // iC= 1460 
vC = 14'b0000001001000100; // vC=  580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110110; // iC= 1398 
vC = 14'b0000001001001111; // vC=  591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101110; // iC= 1326 
vC = 14'b0000001000100101; // vC=  549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100000; // iC= 1440 
vC = 14'b0000001000000100; // vC=  516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011000; // iC= 1432 
vC = 14'b0000001000100101; // vC=  549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101011; // iC= 1387 
vC = 14'b0000001000001101; // vC=  525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000100; // iC= 1412 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100011; // iC= 1379 
vC = 14'b0000000111011110; // vC=  478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100111; // iC= 1447 
vC = 14'b0000001001101010; // vC=  618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100110; // iC= 1382 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000001000100100; // vC=  548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000001; // iC= 1345 
vC = 14'b0000001001010111; // vC=  599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001010; // iC= 1290 
vC = 14'b0000001000011000; // vC=  536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001100; // iC= 1292 
vC = 14'b0000001000111111; // vC=  575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111100; // iC= 1340 
vC = 14'b0000001010000000; // vC=  640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100010; // iC= 1314 
vC = 14'b0000001000010001; // vC=  529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111110; // iC= 1278 
vC = 14'b0000001001011000; // vC=  600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000100; // iC= 1284 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111111; // iC= 1279 
vC = 14'b0000001000000010; // vC=  514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100011; // iC= 1379 
vC = 14'b0000001001111010; // vC=  634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011100; // iC= 1372 
vC = 14'b0000001000101110; // vC=  558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000010; // iC= 1410 
vC = 14'b0000001010000000; // vC=  640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100010; // iC= 1250 
vC = 14'b0000001001110000; // vC=  624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100111; // iC= 1319 
vC = 14'b0000001010010001; // vC=  657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110011; // iC= 1395 
vC = 14'b0000001001010111; // vC=  599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111010; // iC= 1338 
vC = 14'b0000001000110010; // vC=  562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101011; // iC= 1259 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100001; // iC= 1249 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001111; // iC= 1295 
vC = 14'b0000001001100100; // vC=  612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100011; // iC= 1251 
vC = 14'b0000001001100011; // vC=  611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111000; // iC= 1336 
vC = 14'b0000001000111011; // vC=  571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001000; // iC= 1224 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100011; // iC= 1251 
vC = 14'b0000001001111100; // vC=  636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111111; // iC= 1279 
vC = 14'b0000001010100111; // vC=  679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100011; // iC= 1251 
vC = 14'b0000001001000100; // vC=  580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100010; // iC= 1314 
vC = 14'b0000001010100101; // vC=  677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001100; // iC= 1356 
vC = 14'b0000001010111110; // vC=  702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101111; // iC= 1327 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010000; // iC= 1232 
vC = 14'b0000001001101101; // vC=  621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000101; // iC= 1221 
vC = 14'b0000001010001100; // vC=  652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011111; // iC= 1247 
vC = 14'b0000001001110010; // vC=  626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011110; // iC= 1182 
vC = 14'b0000001001111110; // vC=  638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010110; // iC= 1302 
vC = 14'b0000001011101000; // vC=  744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000100; // iC= 1220 
vC = 14'b0000001001110110; // vC=  630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011100; // iC= 1180 
vC = 14'b0000001011000101; // vC=  709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111111; // iC= 1215 
vC = 14'b0000001001111100; // vC=  636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110011; // iC= 1267 
vC = 14'b0000001010010101; // vC=  661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111011; // iC= 1275 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011111; // iC= 1183 
vC = 14'b0000001100001000; // vC=  776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111111; // iC= 1151 
vC = 14'b0000001011111100; // vC=  764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100001; // iC= 1185 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111110; // iC= 1150 
vC = 14'b0000001100100101; // vC=  805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110111; // iC= 1143 
vC = 14'b0000001100001010; // vC=  778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000100; // iC= 1156 
vC = 14'b0000001100011001; // vC=  793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101100; // iC= 1132 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111110; // iC= 1214 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111110; // iC= 1214 
vC = 14'b0000001011010001; // vC=  721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b0000001100101010; // vC=  810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110101; // iC= 1269 
vC = 14'b0000001010111101; // vC=  701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b0000001011110110; // vC=  758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100101; // iC= 1253 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010110; // iC= 1110 
vC = 14'b0000001011010110; // vC=  726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010111; // iC= 1239 
vC = 14'b0000001100100010; // vC=  802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110000; // iC= 1136 
vC = 14'b0000001011100100; // vC=  740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b0000001011000010; // vC=  706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010100; // iC= 1172 
vC = 14'b0000001101000011; // vC=  835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001010; // iC= 1226 
vC = 14'b0000001011100101; // vC=  741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100000; // iC= 1120 
vC = 14'b0000001011101011; // vC=  747 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011000; // iC= 1112 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110101; // iC= 1077 
vC = 14'b0000001100111100; // vC=  828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111101; // iC= 1085 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110011; // iC= 1203 
vC = 14'b0000001011110101; // vC=  757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110110; // iC= 1078 
vC = 14'b0000001101011101; // vC=  861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110011; // iC= 1075 
vC = 14'b0000001011100000; // vC=  736 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011110; // iC= 1182 
vC = 14'b0000001011110111; // vC=  759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011010; // iC= 1114 
vC = 14'b0000001100100001; // vC=  801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110101; // iC= 1077 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101000; // iC= 1064 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010110; // iC= 1046 
vC = 14'b0000001100111010; // vC=  826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001000; // iC= 1096 
vC = 14'b0000001100100000; // vC=  800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110001; // iC= 1073 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111110; // iC= 1022 
vC = 14'b0000001101111111; // vC=  895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011011; // iC= 1115 
vC = 14'b0000001100001000; // vC=  776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110001; // iC= 1073 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110100; // iC= 1012 
vC = 14'b0000001101000000; // vC=  832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001001; // iC= 1033 
vC = 14'b0000001101011011; // vC=  859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110111; // iC= 1015 
vC = 14'b0000001101100011; // vC=  867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111110; // iC= 1086 
vC = 14'b0000001101110010; // vC=  882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100010; // iC= 1122 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101001; // iC= 1065 
vC = 14'b0000001100010100; // vC=  788 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011000; // iC=  984 
vC = 14'b0000001101101111; // vC=  879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010111; // iC= 1111 
vC = 14'b0000001100100111; // vC=  807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101011; // iC= 1003 
vC = 14'b0000001110101101; // vC=  941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111101; // iC= 1085 
vC = 14'b0000001101101000; // vC=  872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101010; // iC= 1066 
vC = 14'b0000001101000011; // vC=  835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010011; // iC= 1107 
vC = 14'b0000001110000101; // vC=  901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000111; // iC= 1031 
vC = 14'b0000001110101000; // vC=  936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001010; // iC= 1098 
vC = 14'b0000001111001100; // vC=  972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b0000001110101100; // vC=  940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111110; // iC= 1086 
vC = 14'b0000001100111011; // vC=  827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101000; // iC= 1000 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101100; // iC= 1068 
vC = 14'b0000001101101001; // vC=  873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100110; // iC=  934 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100110; // iC=  934 
vC = 14'b0000001110011010; // vC=  922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011111; // iC=  991 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110010; // iC=  946 
vC = 14'b0000001101111010; // vC=  890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001111; // iC=  975 
vC = 14'b0000001101010111; // vC=  855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111101; // iC=  957 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001001; // iC=  905 
vC = 14'b0000001111001001; // vC=  969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011100; // iC= 1052 
vC = 14'b0000001101010000; // vC=  848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111011; // iC= 1019 
vC = 14'b0000001101010011; // vC=  851 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111010; // iC= 1018 
vC = 14'b0000001101101111; // vC=  879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111011; // iC=  891 
vC = 14'b0000001111100000; // vC=  992 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111101; // iC=  893 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111111; // iC= 1023 
vC = 14'b0000001110101010; // vC=  938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101100; // iC= 1004 
vC = 14'b0000001110000000; // vC=  896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101111; // iC=  943 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110001; // iC=  945 
vC = 14'b0000001110100101; // vC=  933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000100; // iC=  964 
vC = 14'b0000001110110001; // vC=  945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011100; // iC=  988 
vC = 14'b0000010000000110; // vC= 1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101001; // iC= 1001 
vC = 14'b0000001110110111; // vC=  951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100010; // iC=  930 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011001; // iC=  985 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001011; // iC=  843 
vC = 14'b0000001110010000; // vC=  912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001100; // iC=  908 
vC = 14'b0000001111011110; // vC=  990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011101; // iC=  925 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010101; // iC=  981 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011001; // iC=  857 
vC = 14'b0000001110111001; // vC=  953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110111; // iC=  951 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001101; // iC=  845 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011001; // iC=  921 
vC = 14'b0000001111101011; // vC= 1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011001; // iC=  857 
vC = 14'b0000001110110110; // vC=  950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100111; // iC=  935 
vC = 14'b0000010000011101; // vC= 1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110110; // iC=  950 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001011; // iC=  843 
vC = 14'b0000001110100101; // vC=  933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001000; // iC=  904 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000011; // iC=  899 
vC = 14'b0000001110100110; // vC=  934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110100; // iC=  820 
vC = 14'b0000001111000000; // vC=  960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110101; // iC=  885 
vC = 14'b0000010001000010; // vC= 1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111000; // iC=  888 
vC = 14'b0000010000011101; // vC= 1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000110; // iC=  774 
vC = 14'b0000010000010101; // vC= 1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010010; // iC=  786 
vC = 14'b0000001110101100; // vC=  940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111000; // iC=  888 
vC = 14'b0000010000111000; // vC= 1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100001; // iC=  801 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101101; // iC=  813 
vC = 14'b0000010000111010; // vC= 1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101111; // iC=  815 
vC = 14'b0000001110110100; // vC=  948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010111; // iC=  791 
vC = 14'b0000001110110011; // vC=  947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001101; // iC=  781 
vC = 14'b0000001110111001; // vC=  953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101010; // iC=  746 
vC = 14'b0000001111000000; // vC=  960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000001; // iC=  833 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000011; // iC=  835 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111000; // iC=  760 
vC = 14'b0000010000100110; // vC= 1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010110; // iC=  726 
vC = 14'b0000001111010101; // vC=  981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100011; // iC=  739 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000110; // iC=  774 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001011; // iC=  779 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110101; // iC=  693 
vC = 14'b0000010000100110; // vC= 1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000110; // iC=  838 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011001; // iC=  793 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000000; // iC=  832 
vC = 14'b0000001111100011; // vC=  995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001001; // iC=  713 
vC = 14'b0000010000001010; // vC= 1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010011; // iC=  787 
vC = 14'b0000010000111100; // vC= 1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000000; // iC=  704 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110100; // iC=  756 
vC = 14'b0000010001001000; // vC= 1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101010; // iC=  810 
vC = 14'b0000010001101111; // vC= 1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001111; // iC=  719 
vC = 14'b0000010000000110; // vC= 1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100100; // iC=  740 
vC = 14'b0000001111101000; // vC= 1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001111; // iC=  655 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010001; // iC=  785 
vC = 14'b0000001111101100; // vC= 1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110101; // iC=  693 
vC = 14'b0000010000110001; // vC= 1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111101; // iC=  701 
vC = 14'b0000010001010011; // vC= 1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111101; // iC=  765 
vC = 14'b0000010000000100; // vC= 1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011011; // iC=  731 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011110; // iC=  670 
vC = 14'b0000010000100100; // vC= 1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111001; // iC=  697 
vC = 14'b0000010001000001; // vC= 1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100001; // iC=  673 
vC = 14'b0000010000010001; // vC= 1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100010; // iC=  610 
vC = 14'b0000010000101111; // vC= 1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010110; // iC=  662 
vC = 14'b0000010000011010; // vC= 1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010101; // iC=  725 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111000; // iC=  632 
vC = 14'b0000010001111011; // vC= 1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000111; // iC=  711 
vC = 14'b0000010010011101; // vC= 1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010100; // iC=  724 
vC = 14'b0000010001111000; // vC= 1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100000; // iC=  672 
vC = 14'b0000010000000111; // vC= 1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011110; // iC=  670 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110100; // iC=  564 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101011; // iC=  683 
vC = 14'b0000010000110110; // vC= 1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000001; // iC=  577 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111011; // iC=  571 
vC = 14'b0000010000011101; // vC= 1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111111; // iC=  639 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110001; // iC=  689 
vC = 14'b0000010000111100; // vC= 1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110011; // iC=  627 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010101; // iC=  597 
vC = 14'b0000010000100111; // vC= 1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110010; // iC=  626 
vC = 14'b0000010001000110; // vC= 1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110100; // iC=  628 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011000; // iC=  536 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101001; // iC=  553 
vC = 14'b0000010001111000; // vC= 1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010100; // iC=  532 
vC = 14'b0000010010001001; // vC= 1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001001; // iC=  521 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100100; // iC=  612 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001101; // iC=  525 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101100; // iC=  620 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110011; // iC=  627 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001110; // iC=  590 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010111; // iC=  599 
vC = 14'b0000010010000001; // vC= 1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111110; // iC=  510 
vC = 14'b0000010010000010; // vC= 1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011010; // iC=  602 
vC = 14'b0000010000110101; // vC= 1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111111; // iC=  511 
vC = 14'b0000010001000111; // vC= 1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100010; // iC=  482 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010101; // iC=  533 
vC = 14'b0000010010001111; // vC= 1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111111; // iC=  575 
vC = 14'b0000010010000100; // vC= 1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011110; // iC=  542 
vC = 14'b0000010011000001; // vC= 1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100011; // iC=  483 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000001; // iC=  449 
vC = 14'b0000010000110110; // vC= 1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101111; // iC=  431 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011001; // iC=  409 
vC = 14'b0000010011001111; // vC= 1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010100; // iC=  468 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010011; // iC=  467 
vC = 14'b0000010011001101; // vC= 1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001111; // iC=  527 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101011; // iC=  427 
vC = 14'b0000010010100011; // vC= 1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011011; // iC=  539 
vC = 14'b0000010000111001; // vC= 1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001110; // iC=  398 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100110; // iC=  486 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010100; // iC=  404 
vC = 14'b0000010001111001; // vC= 1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110101; // iC=  437 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000110; // iC=  518 
vC = 14'b0000010010010111; // vC= 1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101001; // iC=  489 
vC = 14'b0000010010101110; // vC= 1198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101110; // iC=  366 
vC = 14'b0000010001010110; // vC= 1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111100; // iC=  444 
vC = 14'b0000010010110011; // vC= 1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100111; // iC=  359 
vC = 14'b0000010011001110; // vC= 1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010100; // iC=  404 
vC = 14'b0000010001111100; // vC= 1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011001; // iC=  345 
vC = 14'b0000010001111101; // vC= 1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111101; // iC=  381 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010101; // iC=  469 
vC = 14'b0000010010000000; // vC= 1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011000; // iC=  408 
vC = 14'b0000010001110110; // vC= 1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101110; // iC=  366 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000100; // iC=  324 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000110; // iC=  390 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000110; // iC=  390 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001011; // iC=  267 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111100; // iC=  380 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101001; // iC=  361 
vC = 14'b0000010010011001; // vC= 1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111011; // iC=  251 
vC = 14'b0000010011011001; // vC= 1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100101; // iC=  293 
vC = 14'b0000010001100101; // vC= 1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010000; // iC=  336 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010111; // iC=  343 
vC = 14'b0000010011010001; // vC= 1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101000; // iC=  232 
vC = 14'b0000010001011010; // vC= 1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001100; // iC=  332 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111110; // iC=  254 
vC = 14'b0000010001011110; // vC= 1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010000; // iC=  272 
vC = 14'b0000010011011001; // vC= 1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111111; // iC=  191 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111111; // iC=  191 
vC = 14'b0000010001011100; // vC= 1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000110; // iC=  134 
vC = 14'b0000010011010110; // vC= 1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110010; // iC=  242 
vC = 14'b0000010010101000; // vC= 1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110100; // iC=  116 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100000; // iC=  224 
vC = 14'b0000010010011001; // vC= 1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010100; // iC=   84 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111100; // iC=  188 
vC = 14'b0000010011010110; // vC= 1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100010; // iC=   98 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101100; // iC=  108 
vC = 14'b0000010001010010; // vC= 1106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000001; // iC=  129 
vC = 14'b0000010001111000; // vC= 1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111001; // iC=   -7 
vC = 14'b0000010010110010; // vC= 1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110100; // iC=   52 
vC = 14'b0000010001111000; // vC= 1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000011; // iC=    3 
vC = 14'b0000010001111101; // vC= 1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001110; // iC=   14 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111001; // iC=   -7 
vC = 14'b0000010011010111; // vC= 1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000010; // iC=    2 
vC = 14'b0000010011010011; // vC= 1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111110; // iC=  -66 
vC = 14'b0000010011000100; // vC= 1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010011; // iC= -109 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100011; // iC=  -29 
vC = 14'b0000010010010111; // vC= 1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010101; // iC=  -43 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010101; // iC= -107 
vC = 14'b0000010010101001; // vC= 1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101110; // iC=  -82 
vC = 14'b0000010001111011; // vC= 1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110111; // iC=  -73 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011010; // iC= -166 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010100; // iC= -172 
vC = 14'b0000010011000110; // vC= 1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001000; // iC= -120 
vC = 14'b0000010001111101; // vC= 1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110101; // iC= -139 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011000; // iC= -232 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111111; // iC= -321 
vC = 14'b0000010001001000; // vC= 1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101010; // iC= -214 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011101; // iC= -291 
vC = 14'b0000010011011001; // vC= 1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001011; // iC= -245 
vC = 14'b0000010000111111; // vC= 1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000011; // iC= -317 
vC = 14'b0000010001010101; // vC= 1109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000000; // iC= -320 
vC = 14'b0000010001110000; // vC= 1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101100; // iC= -340 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111000; // iC= -392 
vC = 14'b0000010000110001; // vC= 1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111101; // iC= -323 
vC = 14'b0000010000111100; // vC= 1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111110; // iC= -386 
vC = 14'b0000010001110110; // vC= 1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011110; // iC= -482 
vC = 14'b0000010010000011; // vC= 1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110100; // iC= -396 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010100; // iC= -428 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110001; // iC= -527 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100101; // iC= -539 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000001; // iC= -511 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001010; // iC= -630 
vC = 14'b0000010010001101; // vC= 1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000000; // iC= -640 
vC = 14'b0000010010001101; // vC= 1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100110; // iC= -538 
vC = 14'b0000010010100010; // vC= 1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101111; // iC= -593 
vC = 14'b0000010010100101; // vC= 1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001010; // iC= -630 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000101; // iC= -699 
vC = 14'b0000010000010110; // vC= 1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000010; // iC= -766 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100001; // iC= -671 
vC = 14'b0000010001111101; // vC= 1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100011; // iC= -733 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100001; // iC= -671 
vC = 14'b0000010010010100; // vC= 1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111110; // iC= -770 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011000; // iC= -744 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100111; // iC= -729 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001011; // iC= -821 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001000; // iC= -824 
vC = 14'b0000010001110000; // vC= 1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110111; // iC= -841 
vC = 14'b0000010001101101; // vC= 1133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111110; // iC= -834 
vC = 14'b0000010000001001; // vC= 1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001100; // iC= -884 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111011; // iC= -837 
vC = 14'b0000010010000001; // vC= 1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001001; // iC= -951 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b0000010000100000; // vC= 1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101001; // iC= -983 
vC = 14'b0000001111010111; // vC=  983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101000; // iC= -984 
vC = 14'b0000010000111001; // vC= 1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100011; // iC= -925 
vC = 14'b0000010000110100; // vC= 1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111010; // iC= -966 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101011; // iC=-1109 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101111; // iC=-1041 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000100; // iC=-1084 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010100; // iC=-1068 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101001; // iC=-1175 
vC = 14'b0000010000101100; // vC= 1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101001; // iC=-1047 
vC = 14'b0000001111000001; // vC=  961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101011; // iC=-1173 
vC = 14'b0000001111111110; // vC= 1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001010; // iC=-1078 
vC = 14'b0000010000100101; // vC= 1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110010; // iC=-1230 
vC = 14'b0000001110111111; // vC=  959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100100; // iC=-1180 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010111; // iC=-1257 
vC = 14'b0000010000100010; // vC= 1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100010; // iC=-1246 
vC = 14'b0000010000001000; // vC= 1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010000; // iC=-1264 
vC = 14'b0000001110010010; // vC=  914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110000; // iC=-1232 
vC = 14'b0000001110100011; // vC=  931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011001; // iC=-1255 
vC = 14'b0000001111101110; // vC= 1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110000; // iC=-1296 
vC = 14'b0000001110100100; // vC=  932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b0000010000010000; // vC= 1040 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101100; // iC=-1300 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100100; // iC=-1308 
vC = 14'b0000001111001000; // vC=  968 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100011; // iC=-1245 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110101; // iC=-1291 
vC = 14'b0000001111000001; // vC=  961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001101; // iC=-1395 
vC = 14'b0000001111101000; // vC= 1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100100; // iC=-1308 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101011; // iC=-1301 
vC = 14'b0000001110111111; // vC=  959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001001; // iC=-1399 
vC = 14'b0000001110110101; // vC=  949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b0000001111010110; // vC=  982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110111; // iC=-1353 
vC = 14'b0000001101001100; // vC=  844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b0000001111010111; // vC=  983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001100; // iC=-1396 
vC = 14'b0000001110011011; // vC=  923 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b0000001101000110; // vC=  838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001110; // iC=-1394 
vC = 14'b0000001101101001; // vC=  873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101011; // iC=-1365 
vC = 14'b0000001101010001; // vC=  849 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b0000001101100000; // vC=  864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b0000001101010010; // vC=  850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b0000001110100101; // vC=  933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110011; // iC=-1421 
vC = 14'b0000001100101000; // vC=  808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b0000001100111110; // vC=  830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110010; // iC=-1486 
vC = 14'b0000001110011100; // vC=  924 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b0000001100010101; // vC=  789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b0000001100001001; // vC=  777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001011; // iC=-1461 
vC = 14'b0000001100100010; // vC=  802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111001; // iC=-1479 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011000; // iC=-1448 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110111; // iC=-1545 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b0000001101011101; // vC=  861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b0000001100101010; // vC=  810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b0000001011110000; // vC=  752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010100; // iC=-1580 
vC = 14'b0000001100001010; // vC=  778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b0000001011010010; // vC=  722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b0000001011111111; // vC=  767 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100011; // iC=-1501 
vC = 14'b0000001011100110; // vC=  742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b0000001100101000; // vC=  808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001101; // iC=-1587 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110110; // iC=-1610 
vC = 14'b0000001100110110; // vC=  822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010111; // iC=-1449 
vC = 14'b0000001100001101; // vC=  781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b0000001100000111; // vC=  775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b0000001011110101; // vC=  757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b0000001010000111; // vC=  647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000100; // iC=-1468 
vC = 14'b0000001011101100; // vC=  748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b0000001011101010; // vC=  746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110101; // iC=-1483 
vC = 14'b0000001010111101; // vC=  701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000001011000100; // vC=  708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b0000001011011110; // vC=  734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b0000001011000101; // vC=  709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001101; // iC=-1459 
vC = 14'b0000001010100010; // vC=  674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b0000001010110010; // vC=  690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b0000001011101011; // vC=  747 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b0000001010000111; // vC=  647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b0000001010011001; // vC=  665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b0000001011010011; // vC=  723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101101; // iC=-1619 
vC = 14'b0000001001101000; // vC=  616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111111; // iC=-1537 
vC = 14'b0000001010110101; // vC=  693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b0000001010101111; // vC=  687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b0000001010000111; // vC=  647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110100; // iC=-1612 
vC = 14'b0000001010101100; // vC=  684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b0000001001100101; // vC=  613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101111; // iC=-1617 
vC = 14'b0000001000011000; // vC=  536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000110; // iC=-1466 
vC = 14'b0000001001111101; // vC=  637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b0000001001000001; // vC=  577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000001000100001; // vC=  545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010011; // iC=-1517 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b0000001001110000; // vC=  624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b0000001001111011; // vC=  635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b0000001001000110; // vC=  582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b0000001000110110; // vC=  566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b0000001000100011; // vC=  547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b0000000111110010; // vC=  498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010100; // iC=-1516 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b0000001001001101; // vC=  589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110111; // iC=-1545 
vC = 14'b0000000110111000; // vC=  440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b0000001000011001; // vC=  537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101001; // iC=-1623 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100011; // iC=-1501 
vC = 14'b0000000110110001; // vC=  433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111101; // iC=-1475 
vC = 14'b0000001000011111; // vC=  543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b0000001000000100; // vC=  516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010100; // iC=-1516 
vC = 14'b0000000110111000; // vC=  440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111001; // iC=-1479 
vC = 14'b0000001000100000; // vC=  544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101101; // iC=-1491 
vC = 14'b0000000110111100; // vC=  444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010001; // iC=-1583 
vC = 14'b0000000110110000; // vC=  432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b0000000110111010; // vC=  442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b0000000111101110; // vC=  494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110000; // iC=-1552 
vC = 14'b0000000111111001; // vC=  505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101111; // iC=-1553 
vC = 14'b0000000111101111; // vC=  495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b0000000110000100; // vC=  388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101011; // iC=-1557 
vC = 14'b0000000110111010; // vC=  442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000000110011111; // vC=  415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101011; // iC=-1557 
vC = 14'b0000000110100111; // vC=  423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b0000000101001101; // vC=  333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b0000000110011101; // vC=  413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010100; // iC=-1580 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b0000000110110011; // vC=  435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b0000000101000101; // vC=  325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b0000000101100001; // vC=  353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000000110000110; // vC=  390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b0000000110100110; // vC=  422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b0000000100100011; // vC=  291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001111; // iC=-1521 
vC = 14'b0000000101111101; // vC=  381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b0000000101111111; // vC=  383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100100; // iC=-1500 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b0000000100010011; // vC=  275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b0000000101011111; // vC=  351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000000100010001; // vC=  273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110010; // iC=-1486 
vC = 14'b0000000100101110; // vC=  302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001111; // iC=-1521 
vC = 14'b0000000101011101; // vC=  349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b0000000100110001; // vC=  305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000000101000000; // vC=  320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011011; // iC=-1445 
vC = 14'b0000000011100000; // vC=  224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b0000000011100111; // vC=  231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000000100110001; // vC=  305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110100; // iC=-1548 
vC = 14'b0000000101001001; // vC=  329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b0000000011010010; // vC=  210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010001; // iC=-1455 
vC = 14'b0000000100110110; // vC=  310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001000; // iC=-1464 
vC = 14'b0000000011110111; // vC=  247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001010; // iC=-1526 
vC = 14'b0000000011101110; // vC=  238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011101; // iC=-1507 
vC = 14'b0000000011100010; // vC=  226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010010; // iC=-1582 
vC = 14'b0000000011111110; // vC=  254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b0000000010110011; // vC=  179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001111; // iC=-1521 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010100; // iC=-1516 
vC = 14'b0000000001111101; // vC=  125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011000; // iC=-1448 
vC = 14'b0000000010010010; // vC=  146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b0000000011110010; // vC=  242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b0000000001101001; // vC=  105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101111; // iC=-1553 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011000; // iC=-1448 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001101; // iC=-1459 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111111; // iC=-1473 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b0000000001110100; // vC=  116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b0000000010111111; // vC=  191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000111; // iC=-1401 
vC = 14'b0000000010000100; // vC=  132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011011; // iC=-1445 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001111; // iC=-1457 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000000000100110; // vC=   38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b0000000010010110; // vC=  150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100101; // iC=-1435 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001110; // iC=-1394 
vC = 14'b0000000001001111; // vC=   79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000110; // iC=-1402 
vC = 14'b0000000000011101; // vC=   29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b0000000000100011; // vC=   35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000000000011000; // vC=   24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b1111111111100110; // vC=  -26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001100; // iC=-1396 
vC = 14'b1111111111110010; // vC=  -14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000010; // iC=-1470 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b0000000001011110; // vC=   94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010101; // iC=-1451 
vC = 14'b1111111111110011; // vC=  -13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101000; // iC=-1432 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b1111111111101111; // vC=  -17 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100010; // iC=-1374 
vC = 14'b1111111110101001; // vC=  -87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000011; // iC=-1469 
vC = 14'b0000000000111001; // vC=   57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b1111111110110101; // vC=  -75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b1111111111011010; // vC=  -38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010101; // iC=-1451 
vC = 14'b1111111110100001; // vC=  -95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000111; // iC=-1465 
vC = 14'b1111111110111011; // vC=  -69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100101; // iC=-1371 
vC = 14'b0000000000001010; // vC=   10 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b1111111111000101; // vC=  -59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111000; // iC=-1352 
vC = 14'b1111111111100111; // vC=  -25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000100; // iC=-1404 
vC = 14'b1111111110110100; // vC=  -76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b1111111110000010; // vC= -126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111101; // iC=-1347 
vC = 14'b1111111111000000; // vC=  -64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110011; // iC=-1421 
vC = 14'b1111111110100111; // vC=  -89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101001; // iC=-1367 
vC = 14'b1111111110100000; // vC=  -96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b1111111101011000; // vC= -168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b1111111111010001; // vC=  -47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111111110100000; // vC=  -96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011001; // iC=-1447 
vC = 14'b1111111111001000; // vC=  -56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010110; // iC=-1386 
vC = 14'b1111111111011111; // vC=  -33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101110; // iC=-1362 
vC = 14'b1111111101001000; // vC= -184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000101; // iC=-1339 
vC = 14'b1111111101111101; // vC= -131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011101; // iC=-1443 
vC = 14'b1111111110101010; // vC=  -86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111100; // iC=-1412 
vC = 14'b1111111110100010; // vC=  -94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000100; // iC=-1468 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b1111111110100110; // vC=  -90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001100; // iC=-1332 
vC = 14'b1111111101000010; // vC= -190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111111101001100; // vC= -180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b1111111110001010; // vC= -118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b1111111100011001; // vC= -231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111111110100101; // vC=  -91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b1111111100110010; // vC= -206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101111; // iC=-1297 
vC = 14'b1111111100101100; // vC= -212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011011; // iC=-1381 
vC = 14'b1111111100111101; // vC= -195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000011; // iC=-1405 
vC = 14'b1111111100011000; // vC= -232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b1111111100111111; // vC= -193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111111100101000; // vC= -216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000111; // iC=-1337 
vC = 14'b1111111101011111; // vC= -161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111011; // iC=-1285 
vC = 14'b1111111100010101; // vC= -235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011101; // iC=-1379 
vC = 14'b1111111100110001; // vC= -207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b1111111011011111; // vC= -289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010000; // iC=-1328 
vC = 14'b1111111100101001; // vC= -215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100101; // iC=-1371 
vC = 14'b1111111100110001; // vC= -207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b1111111011100111; // vC= -281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010110; // iC=-1386 
vC = 14'b1111111011111010; // vC= -262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010101; // iC=-1323 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b1111111100010001; // vC= -239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110000; // iC=-1360 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010000; // iC=-1328 
vC = 14'b1111111011000000; // vC= -320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101011; // iC=-1365 
vC = 14'b1111111011001110; // vC= -306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011000; // iC=-1256 
vC = 14'b1111111100100000; // vC= -224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010111; // iC=-1257 
vC = 14'b1111111100001100; // vC= -244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010000; // iC=-1328 
vC = 14'b1111111010100000; // vC= -352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101011; // iC=-1365 
vC = 14'b1111111100000000; // vC= -256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010101; // iC=-1259 
vC = 14'b1111111100100010; // vC= -222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011111; // iC=-1377 
vC = 14'b1111111010001101; // vC= -371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010000; // iC=-1264 
vC = 14'b1111111011100010; // vC= -286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111101; // iC=-1283 
vC = 14'b1111111100000000; // vC= -256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101110; // iC=-1234 
vC = 14'b1111111011011010; // vC= -294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110110; // iC=-1354 
vC = 14'b1111111010001001; // vC= -375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010110; // iC=-1322 
vC = 14'b1111111011010100; // vC= -300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101000; // iC=-1240 
vC = 14'b1111111011001010; // vC= -310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100000; // iC=-1312 
vC = 14'b1111111011100011; // vC= -285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010110; // iC=-1258 
vC = 14'b1111111001100111; // vC= -409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110000; // iC=-1360 
vC = 14'b1111111001110101; // vC= -395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101100; // iC=-1236 
vC = 14'b1111111001111100; // vC= -388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111111011000011; // vC= -317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110100; // iC=-1228 
vC = 14'b1111111011101101; // vC= -275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000011; // iC=-1213 
vC = 14'b1111111010010110; // vC= -362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010100; // iC=-1324 
vC = 14'b1111111010111000; // vC= -328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111111; // iC=-1281 
vC = 14'b1111111010100010; // vC= -350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001101; // iC=-1331 
vC = 14'b1111111011001100; // vC= -308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111101; // iC=-1347 
vC = 14'b1111111010011110; // vC= -354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111101; // iC=-1219 
vC = 14'b1111111001110010; // vC= -398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111000; // iC=-1224 
vC = 14'b1111111001110001; // vC= -399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111010; // iC=-1286 
vC = 14'b1111111010011001; // vC= -359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010010; // iC=-1326 
vC = 14'b1111111001011101; // vC= -419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010111; // iC=-1257 
vC = 14'b1111111000101011; // vC= -469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001100; // iC=-1268 
vC = 14'b1111111010010000; // vC= -368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001101; // iC=-1267 
vC = 14'b1111111010110011; // vC= -333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101100; // iC=-1300 
vC = 14'b1111111001100110; // vC= -410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000111; // iC=-1273 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110010; // iC=-1294 
vC = 14'b1111111000101111; // vC= -465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110010; // iC=-1230 
vC = 14'b1111111010100000; // vC= -352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110100; // iC=-1164 
vC = 14'b1111111000011011; // vC= -485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111101; // iC=-1283 
vC = 14'b1111111000000101; // vC= -507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001010; // iC=-1206 
vC = 14'b1111111000011011; // vC= -485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100111; // iC=-1241 
vC = 14'b1111111001100011; // vC= -413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100001; // iC=-1247 
vC = 14'b1111111001101101; // vC= -403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000110; // iC=-1210 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110100; // iC=-1292 
vC = 14'b1111111001110011; // vC= -397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101001; // iC=-1175 
vC = 14'b1111111001001011; // vC= -437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010111; // iC=-1129 
vC = 14'b1111111000010010; // vC= -494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111010; // iC=-1222 
vC = 14'b1111111001100000; // vC= -416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100001; // iC=-1183 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011101; // iC=-1251 
vC = 14'b1111111001010100; // vC= -428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001000; // iC=-1272 
vC = 14'b1111110111111101; // vC= -515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010011; // iC=-1133 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110000; // iC=-1232 
vC = 14'b1111110111101101; // vC= -531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010010; // iC=-1262 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011100; // iC=-1252 
vC = 14'b1111111000111101; // vC= -451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101110; // iC=-1170 
vC = 14'b1111110111110101; // vC= -523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001100; // iC=-1140 
vC = 14'b1111111000001100; // vC= -500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001001; // iC=-1207 
vC = 14'b1111111000101010; // vC= -470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101000; // iC=-1112 
vC = 14'b1111111000110011; // vC= -461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000000; // iC=-1088 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101101; // iC=-1171 
vC = 14'b1111110111110110; // vC= -522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000001; // iC=-1087 
vC = 14'b1111110111001000; // vC= -568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111100; // iC=-1220 
vC = 14'b1111110111100100; // vC= -540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111000; // iC=-1224 
vC = 14'b1111110111011001; // vC= -551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001100; // iC=-1204 
vC = 14'b1111110110000111; // vC= -633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111111; // iC=-1089 
vC = 14'b1111110110001111; // vC= -625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011111; // iC=-1185 
vC = 14'b1111110111111111; // vC= -513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011001; // iC=-1063 
vC = 14'b1111110111001001; // vC= -567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000110; // iC=-1210 
vC = 14'b1111110110010111; // vC= -617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b1111110110110001; // vC= -591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110111; // iC=-1097 
vC = 14'b1111110111101010; // vC= -534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111101; // iC=-1091 
vC = 14'b1111110111011011; // vC= -549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011011; // iC=-1189 
vC = 14'b1111110110001100; // vC= -628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001101; // iC=-1139 
vC = 14'b1111110111111001; // vC= -519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000000; // iC=-1088 
vC = 14'b1111110110101100; // vC= -596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110011; // iC=-1165 
vC = 14'b1111110111100100; // vC= -540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000000; // iC=-1152 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100011; // iC=-1117 
vC = 14'b1111110110100000; // vC= -608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000011; // iC=-1149 
vC = 14'b1111110111100000; // vC= -544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011001; // iC=-1063 
vC = 14'b1111110110111000; // vC= -584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010110; // iC=-1130 
vC = 14'b1111110111011010; // vC= -550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010110; // iC=-1066 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000110; // iC=-1146 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111110; // iC=-1154 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100001; // iC=-1055 
vC = 14'b1111110101000101; // vC= -699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110101; // iC=-1035 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100011; // iC=-1117 
vC = 14'b1111110110011111; // vC= -609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011001; // iC=-1127 
vC = 14'b1111110100110100; // vC= -716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010110; // iC=-1066 
vC = 14'b1111110110100111; // vC= -601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101011; // iC= -981 
vC = 14'b1111110100110000; // vC= -720 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110000; // iC=-1040 
vC = 14'b1111110101011001; // vC= -679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011111; // iC=-1121 
vC = 14'b1111110101010100; // vC= -684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111111; // iC=-1025 
vC = 14'b1111110101101111; // vC= -657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101010; // iC=-1110 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111010; // iC= -966 
vC = 14'b1111110110101110; // vC= -594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001001; // iC=-1015 
vC = 14'b1111110110010010; // vC= -622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110011; // iC=-1037 
vC = 14'b1111110100101101; // vC= -723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000101; // iC=-1083 
vC = 14'b1111110100011001; // vC= -743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101100; // iC= -980 
vC = 14'b1111110100001000; // vC= -760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000100; // iC=-1020 
vC = 14'b1111110101101010; // vC= -662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101001; // iC= -983 
vC = 14'b1111110110010100; // vC= -620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b1111110100111101; // vC= -707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110011; // iC= -973 
vC = 14'b1111110100110110; // vC= -714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000110; // iC=-1018 
vC = 14'b1111110101011111; // vC= -673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011101; // iC= -931 
vC = 14'b1111110110000100; // vC= -636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000000; // iC= -960 
vC = 14'b1111110100000011; // vC= -765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111011; // iC= -965 
vC = 14'b1111110101011110; // vC= -674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111010; // iC=-1030 
vC = 14'b1111110101100001; // vC= -671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111001; // iC=-1031 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010100; // iC=-1004 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b1111110011011111; // vC= -801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101111; // iC= -977 
vC = 14'b1111110101000100; // vC= -700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001101; // iC=-1011 
vC = 14'b1111110011101000; // vC= -792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111101; // iC= -963 
vC = 14'b1111110011110100; // vC= -780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111000; // iC=-1032 
vC = 14'b1111110011111010; // vC= -774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000011; // iC= -957 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011011; // iC= -933 
vC = 14'b1111110011101000; // vC= -792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010100; // iC= -876 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111100; // iC= -964 
vC = 14'b1111110101001011; // vC= -693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101000; // iC= -984 
vC = 14'b1111110011101000; // vC= -792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100011; // iC= -989 
vC = 14'b1111110101001010; // vC= -694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110001; // iC= -911 
vC = 14'b1111110010111010; // vC= -838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110111; // iC= -969 
vC = 14'b1111110011111110; // vC= -770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111010; // iC= -966 
vC = 14'b1111110100010000; // vC= -752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111011; // iC= -965 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111000; // iC= -840 
vC = 14'b1111110010100001; // vC= -863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101110; // iC= -914 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111111; // iC= -961 
vC = 14'b1111110011100110; // vC= -794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110101; // iC= -971 
vC = 14'b1111110011100011; // vC= -797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000011; // iC= -829 
vC = 14'b1111110100100001; // vC= -735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111110; // iC= -962 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000011; // iC= -893 
vC = 14'b1111110010101101; // vC= -851 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110111; // iC= -841 
vC = 14'b1111110011100010; // vC= -798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001110; // iC= -946 
vC = 14'b1111110010100111; // vC= -857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100001; // iC= -799 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100000; // iC= -864 
vC = 14'b1111110011110111; // vC= -777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100111; // iC= -921 
vC = 14'b1111110011001110; // vC= -818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001110; // iC= -882 
vC = 14'b1111110010000110; // vC= -890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101000; // iC= -856 
vC = 14'b1111110011100011; // vC= -797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100001; // iC= -863 
vC = 14'b1111110010010010; // vC= -878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101101; // iC= -787 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001011; // iC= -821 
vC = 14'b1111110011011110; // vC= -802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011001; // iC= -871 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101110; // iC= -850 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011111; // iC= -801 
vC = 14'b1111110010100001; // vC= -863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110011; // iC= -781 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101101; // iC= -787 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001101; // iC= -819 
vC = 14'b1111110011010010; // vC= -814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001001; // iC= -887 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101100; // iC= -852 
vC = 14'b1111110010010000; // vC= -880 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000110; // iC= -826 
vC = 14'b1111110011001001; // vC= -823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101101; // iC= -787 
vC = 14'b1111110010111000; // vC= -840 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101010; // iC= -854 
vC = 14'b1111110010001011; // vC= -885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110000; // iC= -848 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101000; // iC= -856 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110010; // iC= -782 
vC = 14'b1111110001111001; // vC= -903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001100; // iC= -820 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110010; // iC= -846 
vC = 14'b1111110001111100; // vC= -900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001110; // iC= -818 
vC = 14'b1111110001000011; // vC= -957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110111; // iC= -841 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111100; // iC= -708 
vC = 14'b1111110011001100; // vC= -820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110111; // iC= -841 
vC = 14'b1111110001110011; // vC= -909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100110; // iC= -794 
vC = 14'b1111110010101011; // vC= -853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101100; // iC= -724 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010000; // iC= -688 
vC = 14'b1111110000101001; // vC= -983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010101; // iC= -683 
vC = 14'b1111110001101101; // vC= -915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100110; // iC= -666 
vC = 14'b1111110011000000; // vC= -832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001101; // iC= -819 
vC = 14'b1111110000011111; // vC= -993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111101; // iC= -707 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011110; // iC= -802 
vC = 14'b1111110000100011; // vC= -989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111001; // iC= -647 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011001; // iC= -679 
vC = 14'b1111110001110011; // vC= -909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000111; // iC= -697 
vC = 14'b1111110000100100; // vC= -988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110111; // iC= -777 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011110; // iC= -738 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001100; // iC= -756 
vC = 14'b1111110010100011; // vC= -861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000100; // iC= -700 
vC = 14'b1111110000100101; // vC= -987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110100; // iC= -716 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100000; // iC= -672 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111001; // iC= -711 
vC = 14'b1111110010000110; // vC= -890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011110; // iC= -674 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110100; // iC= -652 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010010; // iC= -750 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000111; // iC= -697 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001011; // iC= -693 
vC = 14'b1111110000010001; // vC=-1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111111; // iC= -705 
vC = 14'b1111110001101000; // vC= -920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100010; // iC= -670 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110100; // iC= -588 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111010; // iC= -710 
vC = 14'b1111110001001111; // vC= -945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000010; // iC= -574 
vC = 14'b1111101111111111; // vC=-1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100001; // iC= -607 
vC = 14'b1111101111101100; // vC=-1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110110; // iC= -650 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111100; // iC= -580 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000000; // iC= -704 
vC = 14'b1111110001110110; // vC= -906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111010; // iC= -582 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111100; // iC= -580 
vC = 14'b1111110000101010; // vC= -982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100111; // iC= -537 
vC = 14'b1111110001110101; // vC= -907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111100; // iC= -580 
vC = 14'b1111101111010101; // vC=-1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011100; // iC= -548 
vC = 14'b1111110000110111; // vC= -969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101001; // iC= -599 
vC = 14'b1111110001000111; // vC= -953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111101; // iC= -579 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001101; // iC= -563 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b1111110000110011; // vC= -973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111101; // iC= -579 
vC = 14'b1111110001100000; // vC= -928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101100; // iC= -532 
vC = 14'b1111110001100110; // vC= -922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011011; // iC= -613 
vC = 14'b1111110001100100; // vC= -924 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111101111110111; // vC=-1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010011; // iC= -493 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100000; // iC= -480 
vC = 14'b1111101111110010; // vC=-1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101010; // iC= -534 
vC = 14'b1111110000110010; // vC= -974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110110; // iC= -586 
vC = 14'b1111101111000011; // vC=-1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010011; // iC= -621 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101111; // iC= -593 
vC = 14'b1111101110111001; // vC=-1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101101; // iC= -467 
vC = 14'b1111110000000011; // vC=-1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001001; // iC= -567 
vC = 14'b1111110000110101; // vC= -971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011011; // iC= -485 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111111; // iC= -577 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000011; // iC= -573 
vC = 14'b1111110000100001; // vC= -991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100000; // iC= -480 
vC = 14'b1111101110110001; // vC=-1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111010; // iC= -582 
vC = 14'b1111110000010100; // vC=-1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111101; // iC= -579 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010101; // iC= -427 
vC = 14'b1111101110111110; // vC=-1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001101; // iC= -563 
vC = 14'b1111101111111000; // vC=-1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b1111110000000010; // vC=-1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111100; // iC= -452 
vC = 14'b1111101111101001; // vC=-1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001000; // iC= -440 
vC = 14'b1111101111000001; // vC=-1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000111; // iC= -441 
vC = 14'b1111101110100001; // vC=-1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111010; // iC= -454 
vC = 14'b1111110000011101; // vC= -995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111001; // iC= -455 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110101; // iC= -523 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110011; // iC= -525 
vC = 14'b1111101110100110; // vC=-1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010001; // iC= -431 
vC = 14'b1111101111001000; // vC=-1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111101; // iC= -451 
vC = 14'b1111101110011100; // vC=-1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100011; // iC= -477 
vC = 14'b1111101110010101; // vC=-1131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011010; // iC= -358 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010100; // iC= -364 
vC = 14'b1111101110010000; // vC=-1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101010; // iC= -406 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001000; // iC= -376 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010101; // iC= -491 
vC = 14'b1111101111010001; // vC=-1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101100; // iC= -340 
vC = 14'b1111101110110111; // vC=-1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101111; // iC= -465 
vC = 14'b1111110000100100; // vC= -988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101101; // iC= -467 
vC = 14'b1111110000010000; // vC=-1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110001; // iC= -335 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110110; // iC= -394 
vC = 14'b1111110000001111; // vC=-1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110000; // iC= -400 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011110; // iC= -354 
vC = 14'b1111101110100010; // vC=-1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111101; // iC= -323 
vC = 14'b1111101110011010; // vC=-1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011000; // iC= -424 
vC = 14'b1111110000000001; // vC=-1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101111; // iC= -337 
vC = 14'b1111101111000100; // vC=-1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010010; // iC= -366 
vC = 14'b1111110000000011; // vC=-1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001111; // iC= -305 
vC = 14'b1111101111111110; // vC=-1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111001; // iC= -327 
vC = 14'b1111101111100010; // vC=-1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111100; // iC= -260 
vC = 14'b1111101110100100; // vC=-1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110010; // iC= -334 
vC = 14'b1111110000001111; // vC=-1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101111; // iC= -401 
vC = 14'b1111101110011010; // vC=-1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110000; // iC= -336 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001101; // iC= -307 
vC = 14'b1111101110011111; // vC=-1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100001; // iC= -351 
vC = 14'b1111101111101100; // vC=-1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101000; // iC= -280 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101101; // iC= -211 
vC = 14'b1111101110100110; // vC=-1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100010; // iC= -286 
vC = 14'b1111110000001001; // vC=-1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011010; // iC= -230 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010010; // iC= -238 
vC = 14'b1111101110111101; // vC=-1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011010; // iC= -294 
vC = 14'b1111101110010111; // vC=-1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010000; // iC= -176 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001010; // iC= -182 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101000; // iC= -216 
vC = 14'b1111101110110010; // vC=-1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000010; // iC= -254 
vC = 14'b1111101110010111; // vC=-1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011101; // iC= -227 
vC = 14'b1111101111000000; // vC=-1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000110; // iC= -186 
vC = 14'b1111101110111101; // vC=-1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110011; // iC=  -77 
vC = 14'b1111101111100110; // vC=-1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111111; // iC= -129 
vC = 14'b1111101111010100; // vC=-1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011101; // iC= -163 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010101; // iC= -171 
vC = 14'b1111101111101011; // vC=-1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110100; // iC=  -76 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010111; // iC= -105 
vC = 14'b1111101111100010; // vC=-1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101100; // iC=  -20 
vC = 14'b1111101110111100; // vC=-1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001001; // iC= -119 
vC = 14'b1111101111101011; // vC=-1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101000; // iC=  -24 
vC = 14'b1111101110001110; // vC=-1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101110; // iC=  -82 
vC = 14'b1111101110111010; // vC=-1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100000; // iC=  -32 
vC = 14'b1111101110111000; // vC=-1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111100; // iC=   -4 
vC = 14'b1111101111000001; // vC=-1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110111; // iC=   55 
vC = 14'b1111101111110001; // vC=-1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110101; // iC=   53 
vC = 14'b1111101110111111; // vC=-1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001110; // iC=   14 
vC = 14'b1111101101100100; // vC=-1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100100; // iC=  164 
vC = 14'b1111101110000011; // vC=-1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000110; // iC=  134 
vC = 14'b1111101111101000; // vC=-1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010000; // iC=   80 
vC = 14'b1111101111000000; // vC=-1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100101; // iC=  165 
vC = 14'b1111101101111001; // vC=-1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101000; // iC=  168 
vC = 14'b1111101110100010; // vC=-1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100001; // iC=  161 
vC = 14'b1111101110100101; // vC=-1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010110; // iC=  278 
vC = 14'b1111101111101001; // vC=-1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010101; // iC=  149 
vC = 14'b1111101101111001; // vC=-1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111100; // iC=  252 
vC = 14'b1111101111011111; // vC=-1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010000; // iC=  272 
vC = 14'b1111101110011001; // vC=-1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001111; // iC=  271 
vC = 14'b1111101111101000; // vC=-1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101010; // iC=  234 
vC = 14'b1111101111010111; // vC=-1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000001; // iC=  321 
vC = 14'b1111101110101100; // vC=-1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010011; // iC=  403 
vC = 14'b1111101111101111; // vC=-1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000001; // iC=  449 
vC = 14'b1111101111010011; // vC=-1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110001; // iC=  369 
vC = 14'b1111101111001011; // vC=-1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010101; // iC=  469 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011111; // iC=  479 
vC = 14'b1111101111100100; // vC=-1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010101; // iC=  405 
vC = 14'b1111101111100001; // vC=-1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101110; // iC=  558 
vC = 14'b1111101110001100; // vC=-1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011111; // iC=  479 
vC = 14'b1111110000010011; // vC=-1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000111; // iC=  455 
vC = 14'b1111101111110110; // vC=-1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011011; // iC=  539 
vC = 14'b1111101110111001; // vC=-1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010000; // iC=  592 
vC = 14'b1111101111101100; // vC=-1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110101; // iC=  629 
vC = 14'b1111101111010110; // vC=-1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010011; // iC=  595 
vC = 14'b1111101111010101; // vC=-1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110100; // iC=  564 
vC = 14'b1111101111010100; // vC=-1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001100; // iC=  588 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001110; // iC=  718 
vC = 14'b1111101110001101; // vC=-1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000011; // iC=  643 
vC = 14'b1111101111001000; // vC=-1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111100; // iC=  700 
vC = 14'b1111101111010011; // vC=-1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110000; // iC=  752 
vC = 14'b1111110000100010; // vC= -990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010000; // iC=  848 
vC = 14'b1111110000100011; // vC= -989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011010; // iC=  730 
vC = 14'b1111101110111001; // vC=-1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100000; // iC=  864 
vC = 14'b1111101111011111; // vC=-1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b1111101111010100; // vC=-1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001010; // iC=  906 
vC = 14'b1111110000011101; // vC= -995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101100; // iC=  876 
vC = 14'b1111110000000011; // vC=-1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100110; // iC=  870 
vC = 14'b1111101111010011; // vC=-1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111111; // iC=  831 
vC = 14'b1111101111111100; // vC=-1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101000; // iC=  872 
vC = 14'b1111110000101110; // vC= -978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011010; // iC=  986 
vC = 14'b1111110000101111; // vC= -977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010000; // iC= 1040 
vC = 14'b1111101111100011; // vC=-1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110000; // iC= 1072 
vC = 14'b1111110001000101; // vC= -955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101001; // iC= 1065 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100111; // iC= 1063 
vC = 14'b1111110000101111; // vC= -977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010010; // iC= 1042 
vC = 14'b1111101111010100; // vC=-1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001010; // iC= 1098 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010110; // iC= 1110 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000111; // iC= 1095 
vC = 14'b1111110000101010; // vC= -982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101000; // iC= 1064 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100100; // iC= 1060 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000110; // iC= 1094 
vC = 14'b1111101111100000; // vC=-1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011010; // iC= 1242 
vC = 14'b1111110001001101; // vC= -947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110011; // iC= 1267 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110110; // iC= 1206 
vC = 14'b1111110000110011; // vC= -973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100010; // iC= 1186 
vC = 14'b1111101111111011; // vC=-1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011100; // iC= 1180 
vC = 14'b1111110001010100; // vC= -940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100010; // iC= 1250 
vC = 14'b1111110010000101; // vC= -891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111110; // iC= 1278 
vC = 14'b1111110001110100; // vC= -908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001000; // iC= 1224 
vC = 14'b1111110000011000; // vC=-1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100110; // iC= 1318 
vC = 14'b1111110001000011; // vC= -957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110001; // iC= 1265 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001001; // iC= 1289 
vC = 14'b1111110010010011; // vC= -877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111111; // iC= 1407 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101011; // iC= 1323 
vC = 14'b1111110001110011; // vC= -909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000110; // iC= 1350 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100110; // iC= 1318 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001000; // iC= 1480 
vC = 14'b1111110000011110; // vC= -994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001110; // iC= 1358 
vC = 14'b1111110001000010; // vC= -958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001101; // iC= 1421 
vC = 14'b1111110010101100; // vC= -852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110110; // iC= 1462 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000110; // iC= 1414 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110111; // iC= 1399 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000011; // iC= 1539 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111101; // iC= 1533 
vC = 14'b1111110010101100; // vC= -852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001010; // iC= 1546 
vC = 14'b1111110001001101; // vC= -947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001111; // iC= 1487 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110001; // iC= 1457 
vC = 14'b1111110011000000; // vC= -832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011000; // iC= 1624 
vC = 14'b1111110010100001; // vC= -863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011010; // iC= 1562 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111110; // iC= 1662 
vC = 14'b1111110011110110; // vC= -778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001101; // iC= 1549 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110001; // iC= 1585 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101011; // iC= 1579 
vC = 14'b1111110011101010; // vC= -790 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b1111110011001000; // vC= -824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000001; // iC= 1601 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101010; // iC= 1578 
vC = 14'b1111110100011111; // vC= -737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b1111110100011011; // vC= -741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111100; // iC= 1596 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110000; // iC= 1648 
vC = 14'b1111110100011100; // vC= -740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011000; // iC= 1688 
vC = 14'b1111110011101010; // vC= -790 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010101; // iC= 1749 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b1111110100100100; // vC= -732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b1111110100001000; // vC= -760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111110; // iC= 1726 
vC = 14'b1111110011111011; // vC= -773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111110; // iC= 1726 
vC = 14'b1111110100100101; // vC= -731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b1111110100011000; // vC= -744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000110; // iC= 1670 
vC = 14'b1111110011110011; // vC= -781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b1111110100100101; // vC= -731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111110100111100; // vC= -708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b1111110101011000; // vC= -680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111111; // iC= 1663 
vC = 14'b1111110101000001; // vC= -703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000100; // iC= 1796 
vC = 14'b1111110110000110; // vC= -634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b1111110110011010; // vC= -614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011000; // iC= 1688 
vC = 14'b1111110101001000; // vC= -696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101011; // iC= 1707 
vC = 14'b1111110110100011; // vC= -605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b1111110110011110; // vC= -610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111110101010111; // vC= -681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000000; // iC= 1792 
vC = 14'b1111110110001001; // vC= -631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111110; // iC= 1726 
vC = 14'b1111110110010010; // vC= -622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b1111110101000011; // vC= -701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111110110000010; // vC= -638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b1111110101010111; // vC= -681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b1111110110001111; // vC= -625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b1111110101110001; // vC= -655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b1111110110100111; // vC= -601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100011; // iC= 1699 
vC = 14'b1111110110101000; // vC= -600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101001; // iC= 1833 
vC = 14'b1111110110100110; // vC= -602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111110111111101; // vC= -515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b1111110111000110; // vC= -570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101011; // iC= 1707 
vC = 14'b1111110111101010; // vC= -534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011111; // iC= 1759 
vC = 14'b1111110111110100; // vC= -524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000010; // iC= 1730 
vC = 14'b1111110101110101; // vC= -651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b1111111000010010; // vC= -494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b1111111000000111; // vC= -505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101011; // iC= 1835 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b1111110110010011; // vC= -621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101000; // iC= 1768 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010001; // iC= 1745 
vC = 14'b1111110110111010; // vC= -582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111110110101000; // vC= -600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b1111111000100010; // vC= -478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010111; // iC= 1751 
vC = 14'b1111110110101100; // vC= -596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110001; // iC= 1841 
vC = 14'b1111111000110001; // vC= -463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b1111111000110100; // vC= -460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011100; // iC= 1820 
vC = 14'b1111111000011100; // vC= -484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b1111111001000001; // vC= -447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b1111111001010001; // vC= -431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100010; // iC= 1762 
vC = 14'b1111110111101111; // vC= -529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b1111111001010000; // vC= -432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b1111111001101000; // vC= -408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b1111111001100101; // vC= -411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b1111111001111011; // vC= -389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011000; // iC= 1688 
vC = 14'b1111111000110001; // vC= -463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b1111111001101010; // vC= -406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100110; // iC= 1830 
vC = 14'b1111111010000000; // vC= -384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011000; // iC= 1752 
vC = 14'b1111111010011011; // vC= -357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b1111111001011101; // vC= -419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b1111111001111010; // vC= -390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b1111111000111011; // vC= -453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111111010001110; // vC= -370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111100; // iC= 1724 
vC = 14'b1111111001011000; // vC= -424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111111001101000; // vC= -408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b1111111011010000; // vC= -304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b1111111011000111; // vC= -313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010011; // iC= 1811 
vC = 14'b1111111001100111; // vC= -409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010011; // iC= 1811 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b1111111001001010; // vC= -438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101001; // iC= 1833 
vC = 14'b1111111011101011; // vC= -277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b1111111010001111; // vC= -369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b1111111001101001; // vC= -407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b1111111001111001; // vC= -391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101000; // iC= 1768 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110101; // iC= 1781 
vC = 14'b1111111001110101; // vC= -395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100000; // iC= 1824 
vC = 14'b1111111010011011; // vC= -357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b1111111010111100; // vC= -324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010011; // iC= 1747 
vC = 14'b1111111011010010; // vC= -302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b1111111010001001; // vC= -375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b1111111011110100; // vC= -268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110000; // iC= 1776 
vC = 14'b1111111100101011; // vC= -213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011100; // iC= 1820 
vC = 14'b1111111010100101; // vC= -347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b1111111100100100; // vC= -220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101101; // iC= 1709 
vC = 14'b1111111010111110; // vC= -322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110001; // iC= 1713 
vC = 14'b1111111101010100; // vC= -172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b1111111100000101; // vC= -251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b1111111011101000; // vC= -280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b1111111011101011; // vC= -277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b1111111101011111; // vC= -161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101100; // iC= 1772 
vC = 14'b1111111101000101; // vC= -187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b1111111101001111; // vC= -177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b1111111100110011; // vC= -205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b1111111101011000; // vC= -168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b1111111011101011; // vC= -277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111110; // iC= 1790 
vC = 14'b1111111100111110; // vC= -194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001000; // iC= 1672 
vC = 14'b1111111100011001; // vC= -231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110100; // iC= 1780 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111111; // iC= 1791 
vC = 14'b1111111101001000; // vC= -184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111001; // iC= 1657 
vC = 14'b1111111110101010; // vC=  -86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b1111111100001110; // vC= -242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b1111111100110100; // vC= -204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b1111111101000001; // vC= -191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b1111111110000101; // vC= -123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100110; // iC= 1766 
vC = 14'b1111111110111101; // vC=  -67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010011; // iC= 1747 
vC = 14'b1111111110111011; // vC=  -69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b1111111110011001; // vC= -103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b1111111101111110; // vC= -130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b1111111110110100; // vC=  -76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011101; // iC= 1693 
vC = 14'b1111111101001110; // vC= -178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b1111111101110110; // vC= -138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111111101111000; // vC= -136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b1111111111100110; // vC=  -26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b1111111111011101; // vC=  -35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b1111111110010101; // vC= -107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110011; // iC= 1651 
vC = 14'b1111111101101110; // vC= -146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001100; // iC= 1676 
vC = 14'b1111111110100101; // vC=  -91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b1111111111101011; // vC=  -21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101000; // iC= 1768 
vC = 14'b1111111110110000; // vC=  -80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101110; // iC= 1710 
vC = 14'b0000000000000100; // vC=    4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b1111111111110100; // vC=  -12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101000; // iC= 1768 
vC = 14'b1111111111100110; // vC=  -26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100111; // iC= 1639 
vC = 14'b1111111111110010; // vC=  -14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b1111111111100000; // vC=  -32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b0000000000001011; // vC=   11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100011; // iC= 1763 
vC = 14'b1111111111000000; // vC=  -64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b1111111110110011; // vC=  -77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110100; // iC= 1716 
vC = 14'b0000000000101110; // vC=   46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000111; // iC= 1671 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000000; // iC= 1664 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010100; // iC= 1620 
vC = 14'b0000000000101011; // vC=   43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111111111101110; // vC=  -18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011000; // iC= 1624 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001100; // iC= 1740 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001100; // iC= 1612 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000111; // iC= 1671 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010011; // iC= 1619 
vC = 14'b0000000000011011; // vC=   27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001011; // iC= 1739 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001000; // iC= 1672 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b0000000000000111; // vC=    7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b0000000000011100; // vC=   28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000000001010110; // vC=   86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000100; // iC= 1732 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001010; // iC= 1738 
vC = 14'b0000000000101001; // vC=   41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001111; // iC= 1679 
vC = 14'b0000000000100001; // vC=   33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010011; // iC= 1683 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b0000000010110001; // vC=  177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b0000000001110110; // vC=  118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b0000000010001110; // vC=  142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101101; // iC= 1581 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001110; // iC= 1614 
vC = 14'b0000000001110010; // vC=  114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000000011000111; // vC=  199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101111; // iC= 1583 
vC = 14'b0000000010000110; // vC=  134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000110; // iC= 1606 
vC = 14'b0000000010011001; // vC=  153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b0000000010111110; // vC=  190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b0000000010110000; // vC=  176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b0000000001111000; // vC=  120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000100; // iC= 1604 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111011; // iC= 1595 
vC = 14'b0000000100010100; // vC=  276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011010; // iC= 1626 
vC = 14'b0000000010111001; // vC=  185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111101; // iC= 1597 
vC = 14'b0000000011110100; // vC=  244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110010; // iC= 1650 
vC = 14'b0000000011000101; // vC=  197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111000; // iC= 1592 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b0000000100100101; // vC=  293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111011; // iC= 1595 
vC = 14'b0000000011101000; // vC=  232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b0000000100001001; // vC=  265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100101; // iC= 1573 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001100; // iC= 1548 
vC = 14'b0000000100010110; // vC=  278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011001; // iC= 1561 
vC = 14'b0000000100111011; // vC=  315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100101; // iC= 1573 
vC = 14'b0000000100010111; // vC=  279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011010; // iC= 1626 
vC = 14'b0000000011101001; // vC=  233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000111; // iC= 1543 
vC = 14'b0000000100011111; // vC=  287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101111; // iC= 1583 
vC = 14'b0000000101001011; // vC=  331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001000; // iC= 1544 
vC = 14'b0000000101001101; // vC=  333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101100; // iC= 1644 
vC = 14'b0000000011111010; // vC=  250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000101; // iC= 1541 
vC = 14'b0000000101100001; // vC=  353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000101; // iC= 1669 
vC = 14'b0000000100111010; // vC=  314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b0000000100101000; // vC=  296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111001; // iC= 1529 
vC = 14'b0000000101100100; // vC=  356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b0000000100100111; // vC=  295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100000; // iC= 1568 
vC = 14'b0000000011111110; // vC=  254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101000; // iC= 1576 
vC = 14'b0000000100010011; // vC=  275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b0000000101010011; // vC=  339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101010; // iC= 1578 
vC = 14'b0000000101000110; // vC=  326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b0000000101000001; // vC=  321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110110; // iC= 1526 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b0000000100111000; // vC=  312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010110; // iC= 1558 
vC = 14'b0000000100111101; // vC=  317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011101; // iC= 1501 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100101; // iC= 1573 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b0000000101000000; // vC=  320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b0000000110111000; // vC=  440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011011; // iC= 1499 
vC = 14'b0000000100110101; // vC=  309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100011; // iC= 1571 
vC = 14'b0000000110000001; // vC=  385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011000; // iC= 1624 
vC = 14'b0000000110101110; // vC=  430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b0000000110001101; // vC=  397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001100; // iC= 1612 
vC = 14'b0000000101111110; // vC=  382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110101; // iC= 1461 
vC = 14'b0000000110111101; // vC=  445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110010; // iC= 1458 
vC = 14'b0000000111101111; // vC=  495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101100; // iC= 1580 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010000; // iC= 1552 
vC = 14'b0000000101111110; // vC=  382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010111; // iC= 1559 
vC = 14'b0000000111001011; // vC=  459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101110; // iC= 1582 
vC = 14'b0000000101101111; // vC=  367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110011; // iC= 1587 
vC = 14'b0000001000001101; // vC=  525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101010; // iC= 1450 
vC = 14'b0000000101111001; // vC=  377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010001; // iC= 1489 
vC = 14'b0000001000010101; // vC=  533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011011; // iC= 1499 
vC = 14'b0000000110000100; // vC=  388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101010; // iC= 1514 
vC = 14'b0000001000001011; // vC=  523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111001; // iC= 1529 
vC = 14'b0000000111111101; // vC=  509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b0000000111011110; // vC=  478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b0000000110111000; // vC=  440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101100; // iC= 1452 
vC = 14'b0000001000011101; // vC=  541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111100; // iC= 1532 
vC = 14'b0000000111110100; // vC=  500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011011; // iC= 1563 
vC = 14'b0000000111111000; // vC=  504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010011; // iC= 1491 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101000; // iC= 1512 
vC = 14'b0000001000101001; // vC=  553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000010; // iC= 1410 
vC = 14'b0000000111011111; // vC=  479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001110; // iC= 1486 
vC = 14'b0000001000100000; // vC=  544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111110; // iC= 1406 
vC = 14'b0000001000011100; // vC=  540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b0000001001000101; // vC=  581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101101; // iC= 1517 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100101; // iC= 1509 
vC = 14'b0000001000101000; // vC=  552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111111; // iC= 1407 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101010; // iC= 1386 
vC = 14'b0000001001101100; // vC=  620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110001; // iC= 1521 
vC = 14'b0000000111110010; // vC=  498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111001; // iC= 1401 
vC = 14'b0000001000110000; // vC=  560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110111; // iC= 1463 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000000; // iC= 1408 
vC = 14'b0000001010001001; // vC=  649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100000; // iC= 1440 
vC = 14'b0000001010000000; // vC=  640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100011; // iC= 1507 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111100; // iC= 1404 
vC = 14'b0000001010010000; // vC=  656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010001; // iC= 1489 
vC = 14'b0000001000001011; // vC=  523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011010; // iC= 1434 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010010; // iC= 1426 
vC = 14'b0000001010011111; // vC=  671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001001; // iC= 1353 
vC = 14'b0000001001011101; // vC=  605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110100; // iC= 1460 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101110; // iC= 1454 
vC = 14'b0000001000010111; // vC=  535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010100; // iC= 1428 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000111; // iC= 1479 
vC = 14'b0000001010110010; // vC=  690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111000; // iC= 1464 
vC = 14'b0000001010110001; // vC=  689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001100; // iC= 1420 
vC = 14'b0000001010110001; // vC=  689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000100; // iC= 1348 
vC = 14'b0000001001011100; // vC=  604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100011; // iC= 1315 
vC = 14'b0000001011000011; // vC=  707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100011; // iC= 1379 
vC = 14'b0000001001110101; // vC=  629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101111; // iC= 1391 
vC = 14'b0000001010100100; // vC=  676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001000; // iC= 1352 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110101; // iC= 1397 
vC = 14'b0000001011000011; // vC=  707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010011; // iC= 1299 
vC = 14'b0000001001001110; // vC=  590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110110; // iC= 1398 
vC = 14'b0000001001100100; // vC=  612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110101; // iC= 1397 
vC = 14'b0000001010110011; // vC=  691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000101; // iC= 1413 
vC = 14'b0000001010001111; // vC=  655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011011; // iC= 1307 
vC = 14'b0000001011011010; // vC=  730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110111; // iC= 1399 
vC = 14'b0000001010001000; // vC=  648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110010; // iC= 1394 
vC = 14'b0000001001111101; // vC=  637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001101; // iC= 1357 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111101; // iC= 1277 
vC = 14'b0000001011100001; // vC=  737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001010; // iC= 1354 
vC = 14'b0000001010001111; // vC=  655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011010; // iC= 1370 
vC = 14'b0000001011110000; // vC=  752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100101; // iC= 1253 
vC = 14'b0000001100010001; // vC=  785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110110; // iC= 1398 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011010; // iC= 1370 
vC = 14'b0000001010010001; // vC=  657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101001; // iC= 1257 
vC = 14'b0000001010110011; // vC=  691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101111; // iC= 1327 
vC = 14'b0000001011100001; // vC=  737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110011; // iC= 1267 
vC = 14'b0000001100100000; // vC=  800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000000; // iC= 1280 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000111; // iC= 1351 
vC = 14'b0000001010100101; // vC=  677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110110; // iC= 1334 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010011; // iC= 1363 
vC = 14'b0000001011011001; // vC=  729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010011; // iC= 1299 
vC = 14'b0000001100010110; // vC=  790 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010110; // iC= 1366 
vC = 14'b0000001101001000; // vC=  840 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010110; // iC= 1302 
vC = 14'b0000001100101000; // vC=  808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001010; // iC= 1290 
vC = 14'b0000001100101100; // vC=  812 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110011; // iC= 1267 
vC = 14'b0000001011010010; // vC=  722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101101; // iC= 1261 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111011; // iC= 1275 
vC = 14'b0000001010111111; // vC=  703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110001; // iC= 1201 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111011; // iC= 1275 
vC = 14'b0000001101010111; // vC=  855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101101; // iC= 1325 
vC = 14'b0000001101001011; // vC=  843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111110; // iC= 1278 
vC = 14'b0000001100000001; // vC=  769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001001; // iC= 1289 
vC = 14'b0000001100001101; // vC=  781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111111; // iC= 1279 
vC = 14'b0000001100101110; // vC=  814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100110; // iC= 1254 
vC = 14'b0000001101111000; // vC=  888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010111; // iC= 1239 
vC = 14'b0000001101101001; // vC=  873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100101; // iC= 1317 
vC = 14'b0000001101011001; // vC=  857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101010; // iC= 1194 
vC = 14'b0000001100000100; // vC=  772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011001; // iC= 1241 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011110; // iC= 1182 
vC = 14'b0000001011110000; // vC=  752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111110; // iC= 1214 
vC = 14'b0000001110001010; // vC=  906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000110; // iC= 1286 
vC = 14'b0000001101100011; // vC=  867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010100; // iC= 1236 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100010; // iC= 1250 
vC = 14'b0000001110010010; // vC=  914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111001; // iC= 1209 
vC = 14'b0000001110011111; // vC=  927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011000; // iC= 1176 
vC = 14'b0000001101100101; // vC=  869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010010; // iC= 1234 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100011; // iC= 1251 
vC = 14'b0000001101110001; // vC=  881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000001; // iC= 1217 
vC = 14'b0000001100101110; // vC=  814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001010; // iC= 1162 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100100; // iC= 1124 
vC = 14'b0000001101011111; // vC=  863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100000; // iC= 1120 
vC = 14'b0000001101111011; // vC=  891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010100; // iC= 1172 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000011; // iC= 1155 
vC = 14'b0000001110011100; // vC=  924 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011110; // iC= 1118 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010010; // iC= 1170 
vC = 14'b0000001101001101; // vC=  845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110000; // iC= 1200 
vC = 14'b0000001101001111; // vC=  847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010010; // iC= 1106 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000001; // iC= 1153 
vC = 14'b0000001101111011; // vC=  891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000000; // iC= 1088 
vC = 14'b0000001101011010; // vC=  858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b0000001101001100; // vC=  844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111101; // iC= 1085 
vC = 14'b0000001110000111; // vC=  903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000001; // iC= 1153 
vC = 14'b0000001110001101; // vC=  909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b0000001110000101; // vC=  901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000001; // iC= 1089 
vC = 14'b0000001101001000; // vC=  840 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001111; // iC= 1167 
vC = 14'b0000001110010100; // vC=  916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010010; // iC= 1106 
vC = 14'b0000001101110011; // vC=  883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011001; // iC= 1049 
vC = 14'b0000001111101000; // vC= 1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010100; // iC= 1172 
vC = 14'b0000001110111001; // vC=  953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011000; // iC= 1176 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010110; // iC= 1110 
vC = 14'b0000001110010100; // vC=  916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111100; // iC= 1084 
vC = 14'b0000010000000010; // vC= 1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110011; // iC= 1139 
vC = 14'b0000001110000011; // vC=  899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100000; // iC= 1056 
vC = 14'b0000001111111011; // vC= 1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001110; // iC= 1038 
vC = 14'b0000001111111000; // vC= 1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000000; // iC= 1152 
vC = 14'b0000001111100011; // vC=  995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010000; // iC= 1040 
vC = 14'b0000001111011100; // vC=  988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110010; // iC= 1074 
vC = 14'b0000001110100001; // vC=  929 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110101; // iC= 1013 
vC = 14'b0000001111010011; // vC=  979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101000; // iC= 1128 
vC = 14'b0000001110010100; // vC=  916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010101; // iC= 1109 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100100; // iC= 1060 
vC = 14'b0000001111000001; // vC=  961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011110; // iC=  990 
vC = 14'b0000001110111111; // vC=  959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010110; // iC=  982 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110001; // iC= 1009 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110110; // iC= 1078 
vC = 14'b0000001110100101; // vC=  933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010011; // iC=  979 
vC = 14'b0000001110101011; // vC=  939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100111; // iC= 1063 
vC = 14'b0000010000000000; // vC= 1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100010; // iC=  994 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001001; // iC= 1033 
vC = 14'b0000010000000010; // vC= 1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011110; // iC= 1054 
vC = 14'b0000010000100001; // vC= 1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101011; // iC=  939 
vC = 14'b0000010000100111; // vC= 1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110011; // iC= 1075 
vC = 14'b0000001111111011; // vC= 1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100001; // iC=  993 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011001; // iC=  921 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010111; // iC=  983 
vC = 14'b0000010000011100; // vC= 1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010010; // iC= 1042 
vC = 14'b0000010000010001; // vC= 1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001001; // iC= 1033 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000010; // iC=  898 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101110; // iC=  942 
vC = 14'b0000010000101011; // vC= 1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101101; // iC=  941 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010110; // iC=  982 
vC = 14'b0000010001011111; // vC= 1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111001; // iC=  889 
vC = 14'b0000010000001100; // vC= 1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101100; // iC=  876 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110001; // iC= 1009 
vC = 14'b0000010000111000; // vC= 1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111010; // iC=  954 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101010; // iC= 1002 
vC = 14'b0000010000000110; // vC= 1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110101; // iC= 1013 
vC = 14'b0000010000001110; // vC= 1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100110; // iC=  998 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011111; // iC=  991 
vC = 14'b0000010000111101; // vC= 1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101000; // iC=  872 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011101; // iC=  925 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101100; // iC=  940 
vC = 14'b0000010001010100; // vC= 1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100000; // iC=  928 
vC = 14'b0000010001010110; // vC= 1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000100; // iC=  964 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011100; // iC=  924 
vC = 14'b0000010000110000; // vC= 1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011100; // iC=  924 
vC = 14'b0000010000000101; // vC= 1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110111; // iC=  823 
vC = 14'b0000010000001000; // vC= 1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001000; // iC=  904 
vC = 14'b0000010001111010; // vC= 1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011111; // iC=  863 
vC = 14'b0000010010001100; // vC= 1164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000011; // iC=  835 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010110; // iC=  918 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000000; // iC=  896 
vC = 14'b0000010001100101; // vC= 1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001111; // iC=  911 
vC = 14'b0000010000101100; // vC= 1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001000; // iC=  840 
vC = 14'b0000010000000001; // vC= 1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100111; // iC=  871 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010011; // iC=  787 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100001; // iC=  865 
vC = 14'b0000010010011101; // vC= 1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110111; // iC=  759 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000101; // iC=  901 
vC = 14'b0000010010010011; // vC= 1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110001; // iC=  881 
vC = 14'b0000010010101011; // vC= 1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010111; // iC=  791 
vC = 14'b0000010001101100; // vC= 1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111100; // iC=  828 
vC = 14'b0000010001011111; // vC= 1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111000; // iC=  760 
vC = 14'b0000010000010111; // vC= 1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111011; // iC=  763 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011100; // iC=  796 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011000; // iC=  728 
vC = 14'b0000010000100010; // vC= 1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001110; // iC=  718 
vC = 14'b0000010001110111; // vC= 1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100010; // iC=  802 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101010; // iC=  746 
vC = 14'b0000010000101000; // vC= 1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101110; // iC=  750 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001101; // iC=  781 
vC = 14'b0000010000101100; // vC= 1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001000; // iC=  712 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000010; // iC=  834 
vC = 14'b0000010001100001; // vC= 1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011010; // iC=  730 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101010; // iC=  746 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011101; // iC=  797 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001000; // iC=  776 
vC = 14'b0000010010000011; // vC= 1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101110; // iC=  750 
vC = 14'b0000010011010110; // vC= 1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000100; // iC=  772 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010000; // iC=  784 
vC = 14'b0000010001111001; // vC= 1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100100; // iC=  804 
vC = 14'b0000010011010011; // vC= 1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000100; // iC=  772 
vC = 14'b0000010001011001; // vC= 1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110101; // iC=  693 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000111; // iC=  711 
vC = 14'b0000010001101001; // vC= 1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010011; // iC=  787 
vC = 14'b0000010010011101; // vC= 1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111010; // iC=  698 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011000; // iC=  728 
vC = 14'b0000010010011010; // vC= 1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011111; // iC=  671 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101100; // iC=  620 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010011; // iC=  659 
vC = 14'b0000010001010100; // vC= 1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010001; // iC=  657 
vC = 14'b0000010011100110; // vC= 1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000111; // iC=  711 
vC = 14'b0000010010100010; // vC= 1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010010; // iC=  658 
vC = 14'b0000010001110011; // vC= 1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111011; // iC=  699 
vC = 14'b0000010011111001; // vC= 1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011010; // iC=  602 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011101; // iC=  733 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010010; // iC=  658 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000010; // iC=  706 
vC = 14'b0000010001100011; // vC= 1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100100; // iC=  676 
vC = 14'b0000010011011000; // vC= 1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011010; // iC=  666 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111001; // iC=  569 
vC = 14'b0000010011100001; // vC= 1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011110; // iC=  606 
vC = 14'b0000010011100010; // vC= 1250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100010; // iC=  610 
vC = 14'b0000010011100001; // vC= 1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100100; // iC=  612 
vC = 14'b0000010011100001; // vC= 1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000111; // iC=  583 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100111; // iC=  679 
vC = 14'b0000010011110111; // vC= 1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101100; // iC=  556 
vC = 14'b0000010011101001; // vC= 1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100000; // iC=  544 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000110; // iC=  582 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110000; // iC=  624 
vC = 14'b0000010010100101; // vC= 1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010001; // iC=  593 
vC = 14'b0000010011111000; // vC= 1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100101; // iC=  613 
vC = 14'b0000010010001101; // vC= 1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110101; // iC=  565 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001111; // iC=  591 
vC = 14'b0000010011111010; // vC= 1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101011; // iC=  555 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111000; // iC=  632 
vC = 14'b0000010010110101; // vC= 1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110100; // iC=  564 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110000; // iC=  624 
vC = 14'b0000010011110011; // vC= 1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010111; // iC=  599 
vC = 14'b0000010011110011; // vC= 1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100000; // iC=  608 
vC = 14'b0000010100001000; // vC= 1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001101; // iC=  461 
vC = 14'b0000010010010011; // vC= 1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111010; // iC=  570 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110100; // iC=  500 
vC = 14'b0000010011111010; // vC= 1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011000; // iC=  600 
vC = 14'b0000010010110010; // vC= 1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000110; // iC=  454 
vC = 14'b0000010011110110; // vC= 1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011000; // iC=  472 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010011; // iC=  531 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101110; // iC=  494 
vC = 14'b0000010011110000; // vC= 1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000000; // iC=  576 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110000; // iC=  432 
vC = 14'b0000010010111001; // vC= 1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010000; // iC=  528 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010010; // iC=  466 
vC = 14'b0000010100011100; // vC= 1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010111; // iC=  471 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001100; // iC=  524 
vC = 14'b0000010010011001; // vC= 1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100000; // iC=  544 
vC = 14'b0000010100101010; // vC= 1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111111; // iC=  383 
vC = 14'b0000010100010100; // vC= 1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010000; // iC=  528 
vC = 14'b0000010011000001; // vC= 1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000101; // iC=  517 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011110; // iC=  414 
vC = 14'b0000010100111000; // vC= 1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000001; // iC=  449 
vC = 14'b0000010011100011; // vC= 1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110101; // iC=  373 
vC = 14'b0000010011101011; // vC= 1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100011; // iC=  419 
vC = 14'b0000010010101100; // vC= 1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010101; // iC=  469 
vC = 14'b0000010011101011; // vC= 1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111110; // iC=  446 
vC = 14'b0000010100110110; // vC= 1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101111; // iC=  495 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101110; // iC=  430 
vC = 14'b0000010011000111; // vC= 1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001110; // iC=  398 
vC = 14'b0000010100110110; // vC= 1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010001; // iC=  401 
vC = 14'b0000010011101110; // vC= 1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011111; // iC=  351 
vC = 14'b0000010011111101; // vC= 1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100100; // iC=  356 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101111; // iC=  367 
vC = 14'b0000010100000010; // vC= 1282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111011; // iC=  315 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100110; // iC=  358 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101010; // iC=  362 
vC = 14'b0000010011000011; // vC= 1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011010; // iC=  346 
vC = 14'b0000010100110000; // vC= 1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100101; // iC=  357 
vC = 14'b0000010011100111; // vC= 1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001001; // iC=  265 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011001; // iC=  281 
vC = 14'b0000010011110000; // vC= 1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110101; // iC=  245 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001010; // iC=  394 
vC = 14'b0000010100111000; // vC= 1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011111; // iC=  287 
vC = 14'b0000010100000101; // vC= 1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101010; // iC=  362 
vC = 14'b0000010101001100; // vC= 1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100010; // iC=  354 
vC = 14'b0000010011100101; // vC= 1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010011; // iC=  339 
vC = 14'b0000010101001000; // vC= 1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110011; // iC=  243 
vC = 14'b0000010010101110; // vC= 1198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100110; // iC=  166 
vC = 14'b0000010011111000; // vC= 1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000011; // iC=  259 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010100; // iC=  148 
vC = 14'b0000010011101101; // vC= 1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110100; // iC=  180 
vC = 14'b0000010011001001; // vC= 1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010000; // iC=  144 
vC = 14'b0000010010111000; // vC= 1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111111; // iC=  255 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111000; // iC=  248 
vC = 14'b0000010011111011; // vC= 1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011100; // iC=  156 
vC = 14'b0000010100111101; // vC= 1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001101; // iC=  141 
vC = 14'b0000010011100100; // vC= 1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011011; // iC=   91 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100101; // iC=  165 
vC = 14'b0000010100011101; // vC= 1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110011; // iC=  115 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001011; // iC=   75 
vC = 14'b0000010101001000; // vC= 1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101101; // iC=   45 
vC = 14'b0000010101000110; // vC= 1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111010; // iC=   58 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101001; // iC=   41 
vC = 14'b0000010100011110; // vC= 1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001001; // iC=   73 
vC = 14'b0000010010110110; // vC= 1206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001010; // iC=  -54 
vC = 14'b0000010011011001; // vC= 1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111111; // iC=  -65 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000111; // iC=    7 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110010; // iC=  -78 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100110; // iC=  -90 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010111; // iC=  -41 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101010; // iC=  -22 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100010; // iC=  -30 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011011; // iC= -101 
vC = 14'b0000010100111110; // vC= 1342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111101; // iC= -195 
vC = 14'b0000010011010000; // vC= 1232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011100; // iC= -164 
vC = 14'b0000010011110100; // vC= 1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110000; // iC= -208 
vC = 14'b0000010011111111; // vC= 1279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010011; // iC= -173 
vC = 14'b0000010011010101; // vC= 1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011100; // iC= -228 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100110; // iC= -218 
vC = 14'b0000010100010110; // vC= 1302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001001; // iC= -183 
vC = 14'b0000010011001100; // vC= 1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100011; // iC= -221 
vC = 14'b0000010100010101; // vC= 1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000011; // iC= -317 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110000; // iC= -336 
vC = 14'b0000010100001111; // vC= 1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010011; // iC= -365 
vC = 14'b0000010010111000; // vC= 1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000011; // iC= -445 
vC = 14'b0000010100010100; // vC= 1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001010; // iC= -438 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011001; // iC= -487 
vC = 14'b0000010011000011; // vC= 1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010100; // iC= -492 
vC = 14'b0000010100100101; // vC= 1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001001; // iC= -503 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000011; // iC= -509 
vC = 14'b0000010100011000; // vC= 1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010110; // iC= -426 
vC = 14'b0000010011010111; // vC= 1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111101; // iC= -579 
vC = 14'b0000010011010000; // vC= 1232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100110; // iC= -602 
vC = 14'b0000010100010100; // vC= 1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110011; // iC= -589 
vC = 14'b0000010011000100; // vC= 1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101111; // iC= -593 
vC = 14'b0000010010000000; // vC= 1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011110; // iC= -674 
vC = 14'b0000010010101100; // vC= 1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000100; // iC= -636 
vC = 14'b0000010011100101; // vC= 1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110011; // iC= -653 
vC = 14'b0000010001111010; // vC= 1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110000; // iC= -720 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101110; // iC= -594 
vC = 14'b0000010010011001; // vC= 1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001001; // iC= -759 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100011; // iC= -797 
vC = 14'b0000010011011001; // vC= 1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100100; // iC= -732 
vC = 14'b0000010011001011; // vC= 1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110010; // iC= -718 
vC = 14'b0000010011010000; // vC= 1232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000001; // iC= -767 
vC = 14'b0000010011011010; // vC= 1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101100; // iC= -788 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001111; // iC= -881 
vC = 14'b0000010010110011; // vC= 1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010101; // iC= -811 
vC = 14'b0000010001111111; // vC= 1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110110; // iC= -778 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110001; // iC= -847 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100010; // iC= -926 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000001; // iC= -895 
vC = 14'b0000010001101001; // vC= 1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100111; // iC= -985 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111100; // iC= -964 
vC = 14'b0000010001000001; // vC= 1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111001; // iC=-1031 
vC = 14'b0000010010110101; // vC= 1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000110; // iC=-1018 
vC = 14'b0000010001000010; // vC= 1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111000; // iC=-1032 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000110; // iC=-1082 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100010; // iC= -990 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111000; // iC=-1096 
vC = 14'b0000010010110010; // vC= 1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110101; // iC=-1099 
vC = 14'b0000010001110000; // vC= 1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100111; // iC=-1113 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010100; // iC=-1004 
vC = 14'b0000010001100000; // vC= 1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110110; // iC=-1162 
vC = 14'b0000010010110110; // vC= 1206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100011; // iC=-1117 
vC = 14'b0000010001010110; // vC= 1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100110; // iC=-1050 
vC = 14'b0000010000111011; // vC= 1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001110; // iC=-1138 
vC = 14'b0000010010101011; // vC= 1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010100; // iC=-1132 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110001; // iC=-1167 
vC = 14'b0000010001101011; // vC= 1131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011101; // iC=-1187 
vC = 14'b0000010000001110; // vC= 1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010000; // iC=-1136 
vC = 14'b0000010001011100; // vC= 1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101111; // iC=-1233 
vC = 14'b0000010001101000; // vC= 1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001011; // iC=-1269 
vC = 14'b0000001111110101; // vC= 1013 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100011; // iC=-1309 
vC = 14'b0000010000110110; // vC= 1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010010; // iC=-1262 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000101; // iC=-1339 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000000; // iC=-1216 
vC = 14'b0000010001010110; // vC= 1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011010; // iC=-1318 
vC = 14'b0000010000101110; // vC= 1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111001; // iC=-1287 
vC = 14'b0000010000001100; // vC= 1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b0000010000100010; // vC= 1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010010; // iC=-1262 
vC = 14'b0000010000010100; // vC= 1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101110; // iC=-1362 
vC = 14'b0000010001000011; // vC= 1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000010; // iC=-1278 
vC = 14'b0000001110110110; // vC=  950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010010; // iC=-1326 
vC = 14'b0000001110110111; // vC=  951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011001; // iC=-1383 
vC = 14'b0000001110101001; // vC=  937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010010; // iC=-1326 
vC = 14'b0000010000010110; // vC= 1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001000; // iC=-1464 
vC = 14'b0000010000100010; // vC= 1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011100; // iC=-1444 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b0000010000110100; // vC= 1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011001; // iC=-1383 
vC = 14'b0000001110111110; // vC=  958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111000; // iC=-1416 
vC = 14'b0000001111011010; // vC=  986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110111; // iC=-1353 
vC = 14'b0000001111011110; // vC=  990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010100; // iC=-1516 
vC = 14'b0000001111000100; // vC=  964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b0000001111001111; // vC=  975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000100; // iC=-1404 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110101; // iC=-1483 
vC = 14'b0000001101110100; // vC=  884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111111; // iC=-1537 
vC = 14'b0000001111011010; // vC=  986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001011; // iC=-1461 
vC = 14'b0000001110110011; // vC=  947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b0000001111110110; // vC= 1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b0000001110111000; // vC=  952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100101; // iC=-1435 
vC = 14'b0000001101101011; // vC=  875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000100; // iC=-1468 
vC = 14'b0000001101011000; // vC=  856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b0000001110111010; // vC=  954 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b0000001110100100; // vC=  932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111101; // iC=-1539 
vC = 14'b0000001110111001; // vC=  953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b0000001101100001; // vC=  865 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b0000001110010111; // vC=  919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b0000001101110011; // vC=  883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110111; // iC=-1481 
vC = 14'b0000001100101010; // vC=  810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100011; // iC=-1565 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011000; // iC=-1448 
vC = 14'b0000001101100100; // vC=  868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000001100100111; // vC=  807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100110; // iC=-1562 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000001100000001; // vC=  769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b0000001110001001; // vC=  905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110101; // iC=-1611 
vC = 14'b0000001100011000; // vC=  792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b0000001100110101; // vC=  821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b0000001101100110; // vC=  870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101011; // iC=-1621 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b0000001100001111; // vC=  783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110101; // iC=-1483 
vC = 14'b0000001100001000; // vC=  776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010111; // iC=-1577 
vC = 14'b0000001011000100; // vC=  708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b0000001011000001; // vC=  705 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111101; // iC=-1539 
vC = 14'b0000001101001110; // vC=  846 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111001; // iC=-1479 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b0000001010101100; // vC=  684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b0000001011101010; // vC=  746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b0000001100000011; // vC=  771 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b0000001100010111; // vC=  791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b0000001100001000; // vC=  776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b0000001100100101; // vC=  805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011101; // iC=-1507 
vC = 14'b0000001010101101; // vC=  685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101010; // iC=-1558 
vC = 14'b0000001011001101; // vC=  717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000001010010101; // vC=  661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b0000001010001110; // vC=  654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b0000001010101000; // vC=  680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b0000001010000001; // vC=  641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b0000001001010010; // vC=  594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b0000001001100011; // vC=  611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b0000001010111110; // vC=  702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000001011000111; // vC=  711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110000; // iC=-1488 
vC = 14'b0000001001011001; // vC=  601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000101; // iC=-1595 
vC = 14'b0000001011010001; // vC=  721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b0000001001111010; // vC=  634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b0000001000101101; // vC=  557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111111; // iC=-1537 
vC = 14'b0000001010000010; // vC=  642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b0000001001110101; // vC=  629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001101; // iC=-1651 
vC = 14'b0000001010000001; // vC=  641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b0000001001001101; // vC=  589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b0000001010011011; // vC=  667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b0000001000011101; // vC=  541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000001010001101; // vC=  653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001100; // iC=-1524 
vC = 14'b0000001000000101; // vC=  517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010010; // iC=-1582 
vC = 14'b0000000111101110; // vC=  494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b0000001000000001; // vC=  513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010010; // iC=-1646 
vC = 14'b0000001001000110; // vC=  582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000001000100011; // vC=  547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b0000000111011000; // vC=  472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b0000000111110111; // vC=  503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000001001001010; // vC=  586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100100; // iC=-1564 
vC = 14'b0000001000011100; // vC=  540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111100; // iC=-1540 
vC = 14'b0000000111010111; // vC=  471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101010; // iC=-1558 
vC = 14'b0000001000011011; // vC=  539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b0000000111111000; // vC=  504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000010; // iC=-1534 
vC = 14'b0000000110111001; // vC=  441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b0000000111110011; // vC=  499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000000111100110; // vC=  486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b0000000111011011; // vC=  475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011101; // iC=-1571 
vC = 14'b0000000111110111; // vC=  503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b0000000111011010; // vC=  474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b0000001000010101; // vC=  533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b0000000111110011; // vC=  499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b0000000111101010; // vC=  490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000000111011110; // vC=  478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010111; // iC=-1513 
vC = 14'b0000000110000111; // vC=  391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010100; // iC=-1644 
vC = 14'b0000000110011011; // vC=  411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b0000000110001101; // vC=  397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b0000000101011000; // vC=  344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011001; // iC=-1639 
vC = 14'b0000000101100110; // vC=  358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b0000000110101101; // vC=  429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100111; // iC=-1497 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b0000000101001010; // vC=  330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101111; // iC=-1617 
vC = 14'b0000000110010110; // vC=  406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b0000000101000100; // vC=  324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101110; // iC=-1618 
vC = 14'b0000000110011111; // vC=  415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b0000000110101101; // vC=  429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111011; // iC=-1541 
vC = 14'b0000000100010011; // vC=  275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b0000000100110011; // vC=  307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b0000000100011001; // vC=  281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b0000000110001101; // vC=  397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000000100111110; // vC=  318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b0000000101100110; // vC=  358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b0000000011111110; // vC=  254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110001; // iC=-1487 
vC = 14'b0000000101101011; // vC=  363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011111; // iC=-1505 
vC = 14'b0000000100111000; // vC=  312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001111; // iC=-1521 
vC = 14'b0000000011010111; // vC=  215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111110; // iC=-1538 
vC = 14'b0000000100101110; // vC=  302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b0000000101000110; // vC=  326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101111; // iC=-1553 
vC = 14'b0000000101001001; // vC=  329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b0000000101010111; // vC=  343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000000011010100; // vC=  212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b0000000100000000; // vC=  256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b0000000100110001; // vC=  305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000010; // iC=-1534 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001100; // iC=-1524 
vC = 14'b0000000100001011; // vC=  267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b0000000011000101; // vC=  197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000001; // iC=-1599 
vC = 14'b0000000011110010; // vC=  242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b0000000100011010; // vC=  282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b0000000011001100; // vC=  204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101011; // iC=-1493 
vC = 14'b0000000010100100; // vC=  164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b0000000100010011; // vC=  275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101101; // iC=-1491 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b0000000011000000; // vC=  192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b0000000001111010; // vC=  122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110100; // iC=-1548 
vC = 14'b0000000011111111; // vC=  255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b0000000011010011; // vC=  211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b0000000011101000; // vC=  232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110100; // iC=-1612 
vC = 14'b0000000011100011; // vC=  227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110100; // iC=-1548 
vC = 14'b0000000001111111; // vC=  127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110001; // iC=-1551 
vC = 14'b0000000001100101; // vC=  101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001111; // iC=-1521 
vC = 14'b0000000000111110; // vC=   62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b0000000010110110; // vC=  182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b0000000001011110; // vC=   94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b0000000000111011; // vC=   59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b0000000001001110; // vC=   78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b0000000000000110; // vC=    6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b0000000000111011; // vC=   59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101101; // iC=-1555 
vC = 14'b0000000001011000; // vC=   88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b0000000000010001; // vC=   17 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000011; // iC=-1469 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b1111111111100111; // vC=  -25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010100; // iC=-1516 
vC = 14'b0000000000101010; // vC=   42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b1111111111110110; // vC=  -10 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101101; // iC=-1491 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000000000101100; // vC=   44 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101010; // iC=-1430 
vC = 14'b1111111111101001; // vC=  -23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011000; // iC=-1448 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011101; // iC=-1443 
vC = 14'b0000000000100001; // vC=   33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b0000000000011000; // vC=   24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b0000000001000111; // vC=   71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b1111111111011111; // vC=  -33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010101; // iC=-1451 
vC = 14'b0000000000110000; // vC=   48 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b1111111110110111; // vC=  -73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b0000000000000001; // vC=    1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b0000000000011101; // vC=   29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b1111111110011111; // vC=  -97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b1111111111001110; // vC=  -50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011111; // iC=-1505 
vC = 14'b1111111111101110; // vC=  -18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b1111111111000101; // vC=  -59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b1111111111001011; // vC=  -53 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001111; // iC=-1457 
vC = 14'b1111111110011001; // vC= -103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100100; // iC=-1436 
vC = 14'b1111111111010101; // vC=  -43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011101; // iC=-1443 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b1111111101011110; // vC= -162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b1111111110110110; // vC=  -74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b1111111110010110; // vC= -106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b1111111101101110; // vC= -146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b1111111101011000; // vC= -168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111110; // iC=-1538 
vC = 14'b1111111101101011; // vC= -149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b1111111110000100; // vC= -124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b1111111111001100; // vC=  -52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110100; // iC=-1420 
vC = 14'b1111111101001000; // vC= -184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000100; // iC=-1468 
vC = 14'b1111111101110001; // vC= -143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110011; // iC=-1421 
vC = 14'b1111111101101101; // vC= -147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b1111111110100101; // vC=  -91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b1111111101011110; // vC= -162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000010; // iC=-1470 
vC = 14'b1111111100101100; // vC= -212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011110; // iC=-1378 
vC = 14'b1111111101101010; // vC= -150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100011; // iC=-1437 
vC = 14'b1111111100111111; // vC= -193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b1111111101110100; // vC= -140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100100; // iC=-1372 
vC = 14'b1111111101000010; // vC= -190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101011; // iC=-1429 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000110; // iC=-1466 
vC = 14'b1111111011101011; // vC= -277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b1111111100011011; // vC= -229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001100; // iC=-1396 
vC = 14'b1111111011101010; // vC= -278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b1111111101110000; // vC= -144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000001; // iC=-1407 
vC = 14'b1111111100111000; // vC= -200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b1111111101001001; // vC= -183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101010; // iC=-1366 
vC = 14'b1111111100000001; // vC= -255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111101; // iC=-1347 
vC = 14'b1111111101001010; // vC= -182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101000; // iC=-1368 
vC = 14'b1111111011010000; // vC= -304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001001; // iC=-1399 
vC = 14'b1111111011111011; // vC= -261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111111011000010; // vC= -318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011011; // iC=-1445 
vC = 14'b1111111011101100; // vC= -276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b1111111100000101; // vC= -251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000010; // iC=-1342 
vC = 14'b1111111011100110; // vC= -282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101100; // iC=-1428 
vC = 14'b1111111011010100; // vC= -300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110101; // iC=-1483 
vC = 14'b1111111100001011; // vC= -245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011111; // iC=-1377 
vC = 14'b1111111100000011; // vC= -253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000111; // iC=-1337 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100101; // iC=-1435 
vC = 14'b1111111010000110; // vC= -378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b1111111011010111; // vC= -297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101011; // iC=-1365 
vC = 14'b1111111010010001; // vC= -367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110110; // iC=-1354 
vC = 14'b1111111011011010; // vC= -294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111100; // iC=-1348 
vC = 14'b1111111010001111; // vC= -369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100000; // iC=-1312 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111111010101101; // vC= -339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001101; // iC=-1395 
vC = 14'b1111111011011001; // vC= -295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010101; // iC=-1387 
vC = 14'b1111111011010111; // vC= -297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111110; // iC=-1346 
vC = 14'b1111111010001011; // vC= -373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b1111111010010110; // vC= -362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000110; // iC=-1402 
vC = 14'b1111111011100011; // vC= -285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101100; // iC=-1364 
vC = 14'b1111111010010001; // vC= -367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101110; // iC=-1362 
vC = 14'b1111111010110001; // vC= -335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b1111111001011110; // vC= -418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011101; // iC=-1379 
vC = 14'b1111111010101010; // vC= -342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001111; // iC=-1329 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000001; // iC=-1279 
vC = 14'b1111111010111011; // vC= -325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111111001000111; // vC= -441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001001; // iC=-1271 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100101; // iC=-1307 
vC = 14'b1111111010100101; // vC= -347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101111; // iC=-1297 
vC = 14'b1111111000011111; // vC= -481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000010; // iC=-1278 
vC = 14'b1111111000101101; // vC= -467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110100; // iC=-1356 
vC = 14'b1111111001010101; // vC= -427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001101; // iC=-1267 
vC = 14'b1111111001110101; // vC= -395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010001; // iC=-1327 
vC = 14'b1111111001101011; // vC= -405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001111; // iC=-1329 
vC = 14'b1111110111110110; // vC= -522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110110; // iC=-1290 
vC = 14'b1111111010000011; // vC= -381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000101; // iC=-1275 
vC = 14'b1111111001001010; // vC= -438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100110; // iC=-1370 
vC = 14'b1111111001100010; // vC= -414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101000; // iC=-1304 
vC = 14'b1111111000001011; // vC= -501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101011; // iC=-1237 
vC = 14'b1111111001101001; // vC= -407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011011; // iC=-1317 
vC = 14'b1111111000111111; // vC= -449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001101; // iC=-1267 
vC = 14'b1111110111010100; // vC= -556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101001; // iC=-1239 
vC = 14'b1111111000011111; // vC= -481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111001; // iC=-1351 
vC = 14'b1111110111101100; // vC= -532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111111; // iC=-1281 
vC = 14'b1111110111111110; // vC= -514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000001; // iC=-1215 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110000; // iC=-1232 
vC = 14'b1111111000000101; // vC= -507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010111; // iC=-1321 
vC = 14'b1111110110111100; // vC= -580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111110111111011; // vC= -517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110101; // iC=-1355 
vC = 14'b1111111000100011; // vC= -477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111001; // iC=-1223 
vC = 14'b1111111000111101; // vC= -451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001101; // iC=-1267 
vC = 14'b1111110111100100; // vC= -540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011101; // iC=-1251 
vC = 14'b1111110110100000; // vC= -608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100111; // iC=-1305 
vC = 14'b1111110111110010; // vC= -526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111010; // iC=-1222 
vC = 14'b1111110110101100; // vC= -596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010000; // iC=-1200 
vC = 14'b1111110111101011; // vC= -533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b1111110110101101; // vC= -595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101010; // iC=-1174 
vC = 14'b1111110111110111; // vC= -521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100111; // iC=-1305 
vC = 14'b1111111000000001; // vC= -511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000110; // iC=-1210 
vC = 14'b1111110111000111; // vC= -569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111001; // iC=-1287 
vC = 14'b1111110111101100; // vC= -532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110001; // iC=-1167 
vC = 14'b1111110110111000; // vC= -584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111011; // iC=-1221 
vC = 14'b1111110110000011; // vC= -637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101110; // iC=-1298 
vC = 14'b1111110111011111; // vC= -545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110001; // iC=-1167 
vC = 14'b1111110101111010; // vC= -646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001001; // iC=-1143 
vC = 14'b1111110110100001; // vC= -607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101001; // iC=-1239 
vC = 14'b1111110111111000; // vC= -520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011100; // iC=-1188 
vC = 14'b1111110110011100; // vC= -612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010010; // iC=-1134 
vC = 14'b1111110110011010; // vC= -614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101100; // iC=-1172 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001101; // iC=-1139 
vC = 14'b1111110101010101; // vC= -683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000010; // iC=-1214 
vC = 14'b1111110101110001; // vC= -655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100100; // iC=-1180 
vC = 14'b1111110101001010; // vC= -694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111010; // iC=-1222 
vC = 14'b1111110110111100; // vC= -580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101110; // iC=-1234 
vC = 14'b1111110101100010; // vC= -670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011110; // iC=-1122 
vC = 14'b1111110110110101; // vC= -587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101101; // iC=-1171 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100010; // iC=-1246 
vC = 14'b1111110101001111; // vC= -689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001011; // iC=-1205 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111101; // iC=-1155 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b1111110100100010; // vC= -734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110011; // iC=-1229 
vC = 14'b1111110100110101; // vC= -715 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000100; // iC=-1148 
vC = 14'b1111110110011011; // vC= -613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010110; // iC=-1194 
vC = 14'b1111110101100110; // vC= -666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110110; // iC=-1226 
vC = 14'b1111110110001101; // vC= -627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110001; // iC=-1103 
vC = 14'b1111110110011111; // vC= -609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110100; // iC=-1100 
vC = 14'b1111110110000001; // vC= -639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000000; // iC=-1088 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b1111110110001100; // vC= -628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111100; // iC=-1156 
vC = 14'b1111110110011010; // vC= -614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000100; // iC=-1148 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011101; // iC=-1187 
vC = 14'b1111110110001111; // vC= -625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001110; // iC=-1074 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111110100101010; // vC= -726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010010; // iC=-1198 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010011; // iC=-1133 
vC = 14'b1111110100000001; // vC= -767 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011011; // iC=-1125 
vC = 14'b1111110101010111; // vC= -681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001100; // iC=-1140 
vC = 14'b1111110101111100; // vC= -644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101111; // iC=-1105 
vC = 14'b1111110100001101; // vC= -755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001101; // iC=-1139 
vC = 14'b1111110100110111; // vC= -713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111101; // iC=-1091 
vC = 14'b1111110011110110; // vC= -778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110001; // iC=-1039 
vC = 14'b1111110011110100; // vC= -780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011000; // iC=-1128 
vC = 14'b1111110100000011; // vC= -765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101010; // iC=-1110 
vC = 14'b1111110011000101; // vC= -827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110011; // iC=-1037 
vC = 14'b1111110101001100; // vC= -692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011111; // iC=-1057 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111001; // iC=-1159 
vC = 14'b1111110100101011; // vC= -725 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011100; // iC=-1124 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011000; // iC=-1128 
vC = 14'b1111110011000101; // vC= -827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010000; // iC=-1072 
vC = 14'b1111110011000010; // vC= -830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101101; // iC=-1107 
vC = 14'b1111110100001110; // vC= -754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101000; // iC=-1048 
vC = 14'b1111110011011100; // vC= -804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100100; // iC= -988 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000010; // iC=-1022 
vC = 14'b1111110011010100; // vC= -812 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010010; // iC=-1006 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100110; // iC= -986 
vC = 14'b1111110010010101; // vC= -875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100010; // iC= -990 
vC = 14'b1111110011101000; // vC= -792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011110; // iC=-1058 
vC = 14'b1111110100100110; // vC= -730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111110; // iC=-1026 
vC = 14'b1111110100000001; // vC= -767 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011010; // iC= -998 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100001; // iC=-1055 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011101; // iC=-1059 
vC = 14'b1111110010000110; // vC= -890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010000; // iC= -944 
vC = 14'b1111110010111110; // vC= -834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000111; // iC=-1017 
vC = 14'b1111110010000011; // vC= -893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010000; // iC= -944 
vC = 14'b1111110010110111; // vC= -841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101110; // iC= -978 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000011; // iC= -957 
vC = 14'b1111110010101110; // vC= -850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001001; // iC= -951 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111100; // iC= -964 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000011; // iC= -957 
vC = 14'b1111110011000101; // vC= -827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100010; // iC=-1054 
vC = 14'b1111110010000101; // vC= -891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010100; // iC= -940 
vC = 14'b1111110010011110; // vC= -866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111110; // iC= -962 
vC = 14'b1111110011110000; // vC= -784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111000; // iC= -904 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010111; // iC= -937 
vC = 14'b1111110010000001; // vC= -895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101000; // iC= -920 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111100; // iC=-1028 
vC = 14'b1111110001100110; // vC= -922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110110; // iC= -906 
vC = 14'b1111110001000101; // vC= -955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111101; // iC= -899 
vC = 14'b1111110010001100; // vC= -884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110110; // iC= -906 
vC = 14'b1111110001110111; // vC= -905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100100; // iC= -860 
vC = 14'b1111110001010100; // vC= -940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110111; // iC= -905 
vC = 14'b1111110001001110; // vC= -946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011100; // iC= -932 
vC = 14'b1111110010001110; // vC= -882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001011; // iC= -949 
vC = 14'b1111110000101011; // vC= -981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110000; // iC= -912 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110000; // iC= -976 
vC = 14'b1111110001011111; // vC= -929 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111011; // iC= -965 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010110; // iC= -874 
vC = 14'b1111110010110110; // vC= -842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111001; // iC= -967 
vC = 14'b1111110010101000; // vC= -856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101100; // iC= -852 
vC = 14'b1111110000110001; // vC= -975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011001; // iC= -871 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011001; // iC= -871 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000010; // iC= -830 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100101; // iC= -923 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000111; // iC= -953 
vC = 14'b1111110010010110; // vC= -874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110000; // iC= -912 
vC = 14'b1111110000001000; // vC=-1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001010; // iC= -822 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101110; // iC= -850 
vC = 14'b1111110001001010; // vC= -950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010001; // iC= -815 
vC = 14'b1111110001110110; // vC= -906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110010; // iC= -910 
vC = 14'b1111101111110110; // vC=-1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011101; // iC= -867 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110111; // iC= -777 
vC = 14'b1111110000001111; // vC=-1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100111; // iC= -857 
vC = 14'b1111110000111111; // vC= -961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100111; // iC= -857 
vC = 14'b1111101111110010; // vC=-1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001010; // iC= -822 
vC = 14'b1111101111110010; // vC=-1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111000; // iC= -904 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011010; // iC= -806 
vC = 14'b1111110010000100; // vC= -892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010010; // iC= -814 
vC = 14'b1111101111111010; // vC=-1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100011; // iC= -797 
vC = 14'b1111101111110101; // vC=-1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101100; // iC= -788 
vC = 14'b1111110000100111; // vC= -985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111110001001000; // vC= -952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101011; // iC= -853 
vC = 14'b1111110001101100; // vC= -916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011101; // iC= -739 
vC = 14'b1111101111111011; // vC=-1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111110; // iC= -834 
vC = 14'b1111110000011110; // vC= -994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111001; // iC= -839 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011010; // iC= -742 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010101; // iC= -811 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000101; // iC= -763 
vC = 14'b1111110000100111; // vC= -985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001011; // iC= -821 
vC = 14'b1111110001000110; // vC= -954 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010111; // iC= -745 
vC = 14'b1111101111110101; // vC=-1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101000; // iC= -728 
vC = 14'b1111110001011100; // vC= -932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010111; // iC= -745 
vC = 14'b1111101111010101; // vC=-1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101110; // iC= -786 
vC = 14'b1111101111001111; // vC=-1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010101; // iC= -747 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100100; // iC= -668 
vC = 14'b1111110000101001; // vC= -983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100101; // iC= -795 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010011; // iC= -685 
vC = 14'b1111110000011111; // vC= -993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011011; // iC= -677 
vC = 14'b1111101111000011; // vC=-1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100001; // iC= -735 
vC = 14'b1111110000011000; // vC=-1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011011; // iC= -677 
vC = 14'b1111110000101011; // vC= -981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110100; // iC= -652 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101110; // iC= -786 
vC = 14'b1111110000110101; // vC= -971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111001; // iC= -711 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001010; // iC= -694 
vC = 14'b1111101111010010; // vC=-1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011101; // iC= -739 
vC = 14'b1111101110010111; // vC=-1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000010; // iC= -638 
vC = 14'b1111101111010111; // vC=-1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100000; // iC= -736 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100000; // iC= -608 
vC = 14'b1111101111100110; // vC=-1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101001; // iC= -727 
vC = 14'b1111101111000111; // vC=-1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010000; // iC= -752 
vC = 14'b1111101110011110; // vC=-1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111011; // iC= -709 
vC = 14'b1111101110001010; // vC=-1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011100; // iC= -612 
vC = 14'b1111101110001001; // vC=-1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101011; // iC= -725 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111001; // iC= -583 
vC = 14'b1111101111110111; // vC=-1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111000; // iC= -584 
vC = 14'b1111101111110101; // vC=-1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110010; // iC= -590 
vC = 14'b1111101111011000; // vC=-1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011110; // iC= -610 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010101; // iC= -619 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011110; // iC= -674 
vC = 14'b1111101110100001; // vC=-1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000100; // iC= -636 
vC = 14'b1111101111010001; // vC=-1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111100; // iC= -644 
vC = 14'b1111101111010010; // vC=-1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111100; // iC= -580 
vC = 14'b1111101110111101; // vC=-1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101110; // iC= -594 
vC = 14'b1111101101110110; // vC=-1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111001; // iC= -647 
vC = 14'b1111101110001101; // vC=-1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101000; // iC= -536 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010010; // iC= -558 
vC = 14'b1111101110000011; // vC=-1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100110; // iC= -538 
vC = 14'b1111101111101011; // vC=-1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001001; // iC= -631 
vC = 14'b1111101111101100; // vC=-1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111110; // iC= -578 
vC = 14'b1111101101011101; // vC=-1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101100; // iC= -596 
vC = 14'b1111101101100110; // vC=-1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001011; // iC= -501 
vC = 14'b1111101111000001; // vC=-1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110010; // iC= -526 
vC = 14'b1111101110100010; // vC=-1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001001; // iC= -567 
vC = 14'b1111101101111011; // vC=-1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101001; // iC= -599 
vC = 14'b1111101111011101; // vC=-1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110101; // iC= -587 
vC = 14'b1111101110011110; // vC=-1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111000; // iC= -584 
vC = 14'b1111101101101011; // vC=-1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010011; // iC= -621 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110111; // iC= -585 
vC = 14'b1111101101110011; // vC=-1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b1111101110001011; // vC=-1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110100; // iC= -524 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101111; // iC= -593 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101110; // iC= -466 
vC = 14'b1111101110101010; // vC=-1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000011; // iC= -445 
vC = 14'b1111101110111000; // vC=-1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010100; // iC= -556 
vC = 14'b1111101111011111; // vC=-1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001001; // iC= -503 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000100; // iC= -572 
vC = 14'b1111101101110111; // vC=-1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010110; // iC= -554 
vC = 14'b1111101110111110; // vC=-1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111001; // iC= -455 
vC = 14'b1111101110110000; // vC=-1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011001; // iC= -423 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011001; // iC= -487 
vC = 14'b1111101110010100; // vC=-1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101000; // iC= -536 
vC = 14'b1111101101100100; // vC=-1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010011; // iC= -429 
vC = 14'b1111101110100111; // vC=-1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001100; // iC= -436 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000011; // iC= -509 
vC = 14'b1111101110000001; // vC=-1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100000; // iC= -480 
vC = 14'b1111101101011000; // vC=-1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100110; // iC= -410 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010100; // iC= -428 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110101; // iC= -459 
vC = 14'b1111101110010110; // vC=-1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111000; // iC= -520 
vC = 14'b1111101110111000; // vC=-1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000111; // iC= -441 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101011; // iC= -405 
vC = 14'b1111101110101011; // vC=-1109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111000; // iC= -392 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011010; // iC= -486 
vC = 14'b1111101100111011; // vC=-1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010110; // iC= -362 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010101; // iC= -491 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110001; // iC= -335 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110111; // iC= -329 
vC = 14'b1111101101010000; // vC=-1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000100; // iC= -380 
vC = 14'b1111101101101010; // vC=-1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001001; // iC= -439 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111100; // iC= -324 
vC = 14'b1111101100111111; // vC=-1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011101; // iC= -355 
vC = 14'b1111101101000110; // vC=-1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011001; // iC= -295 
vC = 14'b1111101101110101; // vC=-1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110011; // iC= -333 
vC = 14'b1111101100111101; // vC=-1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111101; // iC= -323 
vC = 14'b1111101101010100; // vC=-1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111100; // iC= -388 
vC = 14'b1111101101011100; // vC=-1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100010; // iC= -286 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001100; // iC= -308 
vC = 14'b1111101101101101; // vC=-1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010010; // iC= -366 
vC = 14'b1111101110000011; // vC=-1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101001; // iC= -343 
vC = 14'b1111101110010011; // vC=-1133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100100; // iC= -412 
vC = 14'b1111101101010001; // vC=-1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000101; // iC= -251 
vC = 14'b1111101100010100; // vC=-1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110110; // iC= -266 
vC = 14'b1111101101110101; // vC=-1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011111; // iC= -225 
vC = 14'b1111101100010100; // vC=-1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110000; // iC= -336 
vC = 14'b1111101100011011; // vC=-1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111000; // iC= -264 
vC = 14'b1111101011111111; // vC=-1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110011; // iC= -269 
vC = 14'b1111101101101111; // vC=-1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101010; // iC= -342 
vC = 14'b1111101101011011; // vC=-1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010100; // iC= -172 
vC = 14'b1111101100000111; // vC=-1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010010; // iC= -174 
vC = 14'b1111101110011011; // vC=-1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101100; // iC= -212 
vC = 14'b1111101100110101; // vC=-1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001000; // iC= -248 
vC = 14'b1111101101111000; // vC=-1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010100; // iC= -172 
vC = 14'b1111101100001001; // vC=-1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011010; // iC= -166 
vC = 14'b1111101100110011; // vC=-1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001010; // iC= -118 
vC = 14'b1111101100011001; // vC=-1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010101; // iC= -235 
vC = 14'b1111101101010101; // vC=-1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011111; // iC= -161 
vC = 14'b1111101101011100; // vC=-1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100010; // iC=  -94 
vC = 14'b1111101101101101; // vC=-1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010011; // iC= -109 
vC = 14'b1111101101011010; // vC=-1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111111; // iC= -193 
vC = 14'b1111101101100011; // vC=-1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010111; // iC=  -41 
vC = 14'b1111101100001001; // vC=-1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001000; // iC= -120 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111100; // iC=   -4 
vC = 14'b1111101110001110; // vC=-1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000000; // iC=  -64 
vC = 14'b1111101101000010; // vC=-1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011000; // iC=   24 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110111; // iC=   -9 
vC = 14'b1111101110010010; // vC=-1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011100; // iC=  -36 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001111; // iC=  -49 
vC = 14'b1111101100111101; // vC=-1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010011; // iC=   83 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101111; // iC=  111 
vC = 14'b1111101110000000; // vC=-1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001010; // iC=  138 
vC = 14'b1111101100101110; // vC=-1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010001; // iC=  145 
vC = 14'b1111101110010000; // vC=-1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011110; // iC=   94 
vC = 14'b1111101101011000; // vC=-1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000000; // iC=   64 
vC = 14'b1111101101110111; // vC=-1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001010; // iC=  202 
vC = 14'b1111101100110011; // vC=-1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010100; // iC=  212 
vC = 14'b1111101101111100; // vC=-1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100011; // iC=  227 
vC = 14'b1111101100010011; // vC=-1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110101; // iC=  245 
vC = 14'b1111101110000111; // vC=-1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001100; // iC=  268 
vC = 14'b1111101110000110; // vC=-1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110001; // iC=  305 
vC = 14'b1111101100110100; // vC=-1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101001; // iC=  297 
vC = 14'b1111101101011110; // vC=-1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010110; // iC=  342 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110001; // iC=  241 
vC = 14'b1111101101100111; // vC=-1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010001; // iC=  337 
vC = 14'b1111101100001111; // vC=-1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001010; // iC=  330 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111100; // iC=  316 
vC = 14'b1111101110000111; // vC=-1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000111; // iC=  327 
vC = 14'b1111101110010100; // vC=-1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101110; // iC=  494 
vC = 14'b1111101101011101; // vC=-1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001110; // iC=  462 
vC = 14'b1111101110010011; // vC=-1133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011011; // iC=  411 
vC = 14'b1111101101111011; // vC=-1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101101; // iC=  493 
vC = 14'b1111101100100111; // vC=-1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110001; // iC=  561 
vC = 14'b1111101100101110; // vC=-1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100100; // iC=  484 
vC = 14'b1111101110101011; // vC=-1109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111010; // iC=  570 
vC = 14'b1111101110101101; // vC=-1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110101; // iC=  565 
vC = 14'b1111101101101000; // vC=-1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110110; // iC=  630 
vC = 14'b1111101110001000; // vC=-1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011011; // iC=  667 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011001; // iC=  601 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b1111101101010100; // vC=-1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000011; // iC=  707 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111110; // iC=  766 
vC = 14'b1111101110100010; // vC=-1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011111; // iC=  735 
vC = 14'b1111101100101110; // vC=-1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111010; // iC=  826 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110101; // iC=  757 
vC = 14'b1111101100101100; // vC=-1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100010; // iC=  802 
vC = 14'b1111101101110011; // vC=-1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101100; // iC=  748 
vC = 14'b1111101111000101; // vC=-1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000100; // iC=  900 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000110; // iC=  902 
vC = 14'b1111101101110110; // vC=-1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101011; // iC=  939 
vC = 14'b1111101111001111; // vC=-1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001010; // iC=  906 
vC = 14'b1111101101010100; // vC=-1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111000; // iC=  952 
vC = 14'b1111101110001000; // vC=-1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000110; // iC=  902 
vC = 14'b1111101110101111; // vC=-1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001100; // iC= 1036 
vC = 14'b1111101110111100; // vC=-1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001001; // iC= 1033 
vC = 14'b1111101110110100; // vC=-1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110101; // iC=  949 
vC = 14'b1111101111101000; // vC=-1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101001; // iC= 1065 
vC = 14'b1111101110100111; // vC=-1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010011; // iC=  979 
vC = 14'b1111101111101011; // vC=-1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000100; // iC= 1092 
vC = 14'b1111101111101110; // vC=-1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111011; // iC= 1147 
vC = 14'b1111101110010001; // vC=-1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011111; // iC= 1055 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001010; // iC= 1098 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101100; // iC= 1132 
vC = 14'b1111101111010110; // vC=-1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001101; // iC= 1229 
vC = 14'b1111101111111111; // vC=-1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010101; // iC= 1109 
vC = 14'b1111101110110010; // vC=-1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011000; // iC= 1112 
vC = 14'b1111101110110100; // vC=-1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101001; // iC= 1193 
vC = 14'b1111101111110000; // vC=-1040 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101000; // iC= 1192 
vC = 14'b1111101111101010; // vC=-1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001111; // iC= 1295 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001101; // iC= 1229 
vC = 14'b1111101111110011; // vC=-1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100000; // iC= 1312 
vC = 14'b1111101110100110; // vC=-1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010011; // iC= 1299 
vC = 14'b1111101110001111; // vC=-1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111011; // iC= 1403 
vC = 14'b1111101111011001; // vC=-1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101000; // iC= 1320 
vC = 14'b1111110000110011; // vC= -973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111010; // iC= 1338 
vC = 14'b1111101111001000; // vC=-1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001110; // iC= 1358 
vC = 14'b1111101111101010; // vC=-1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100000; // iC= 1376 
vC = 14'b1111101110111001; // vC=-1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110001; // iC= 1393 
vC = 14'b1111110000100000; // vC= -992 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001001; // iC= 1417 
vC = 14'b1111110000000001; // vC=-1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111111; // iC= 1407 
vC = 14'b1111101111000000; // vC=-1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000111; // iC= 1415 
vC = 14'b1111110000111011; // vC= -965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100011; // iC= 1379 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010110; // iC= 1494 
vC = 14'b1111110000101010; // vC= -982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000100; // iC= 1476 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011011; // iC= 1499 
vC = 14'b1111110000011011; // vC= -997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b1111101111110010; // vC=-1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011110; // iC= 1502 
vC = 14'b1111110000110101; // vC= -971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101100; // iC= 1452 
vC = 14'b1111101111100110; // vC=-1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000001; // iC= 1601 
vC = 14'b1111110001000101; // vC= -955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101111; // iC= 1583 
vC = 14'b1111110000110110; // vC= -970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b1111101111110010; // vC=-1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010011; // iC= 1491 
vC = 14'b1111110010010010; // vC= -878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001011; // iC= 1547 
vC = 14'b1111110010011001; // vC= -871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110101; // iC= 1653 
vC = 14'b1111110000000011; // vC=-1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100101; // iC= 1637 
vC = 14'b1111110001000101; // vC= -955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101110; // iC= 1646 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111010; // iC= 1658 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101010; // iC= 1578 
vC = 14'b1111110001000111; // vC= -953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b1111110000111000; // vC= -968 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001101; // iC= 1677 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011100; // iC= 1628 
vC = 14'b1111110010001110; // vC= -882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b1111110000110001; // vC= -975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000000; // iC= 1600 
vC = 14'b1111110010010011; // vC= -877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000111; // iC= 1671 
vC = 14'b1111110010110110; // vC= -842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100001; // iC= 1633 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011011; // iC= 1627 
vC = 14'b1111110010000110; // vC= -890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b1111110001100001; // vC= -927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010001; // iC= 1745 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011000; // iC= 1688 
vC = 14'b1111110010011101; // vC= -867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111110; // iC= 1662 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010001; // iC= 1745 
vC = 14'b1111110011111100; // vC= -772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b1111110001110101; // vC= -907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111001; // iC= 1785 
vC = 14'b1111110011110001; // vC= -783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111111; // iC= 1791 
vC = 14'b1111110011001110; // vC= -818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000110; // iC= 1798 
vC = 14'b1111110011011101; // vC= -803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b1111110011010100; // vC= -812 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b1111110011000110; // vC= -826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b1111110010110110; // vC= -842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011000; // iC= 1752 
vC = 14'b1111110100111100; // vC= -708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b1111110100100110; // vC= -730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111110011001101; // vC= -819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b1111110011101010; // vC= -790 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110010; // iC= 1778 
vC = 14'b1111110011111110; // vC= -770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000010; // iC= 1858 
vC = 14'b1111110101101011; // vC= -661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110100; // iC= 1716 
vC = 14'b1111110100101111; // vC= -721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000100; // iC= 1796 
vC = 14'b1111110100101001; // vC= -727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b1111110101101010; // vC= -662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111110100000111; // vC= -761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b1111110100110110; // vC= -714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000010; // iC= 1794 
vC = 14'b1111110100111010; // vC= -710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110001; // iC= 1713 
vC = 14'b1111110110101110; // vC= -594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111110101001010; // vC= -694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b1111110101001111; // vC= -689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011111; // iC= 1759 
vC = 14'b1111110110000111; // vC= -633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111101; // iC= 1789 
vC = 14'b1111110110010010; // vC= -622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000110; // iC= 1798 
vC = 14'b1111110100101111; // vC= -721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b1111110110100111; // vC= -601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111001; // iC= 1785 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b1111110110111000; // vC= -584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b1111110110001000; // vC= -632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b1111110110001010; // vC= -630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b1111110111000011; // vC= -573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b1111110101110100; // vC= -652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000010; // iC= 1730 
vC = 14'b1111110110001011; // vC= -629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010000; // iC= 1808 
vC = 14'b1111110110000011; // vC= -637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101111; // iC= 1839 
vC = 14'b1111110110010110; // vC= -618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101111; // iC= 1839 
vC = 14'b1111110111011011; // vC= -549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b1111110111001010; // vC= -566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b1111110110110010; // vC= -590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001100; // iC= 1740 
vC = 14'b1111110111100000; // vC= -544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b1111111000111011; // vC= -453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b1111110111111011; // vC= -517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110000; // iC= 1776 
vC = 14'b1111111000100011; // vC= -477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b1111111000001111; // vC= -497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111111000100010; // vC= -478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b1111110111110000; // vC= -528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010101; // iC= 1749 
vC = 14'b1111110111100110; // vC= -538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111111001010111; // vC= -425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b1111111001001001; // vC= -439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b1111110111100111; // vC= -537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010101; // iC= 1749 
vC = 14'b1111111001010011; // vC= -429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b1111111000111101; // vC= -451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000100; // iC= 1796 
vC = 14'b1111111000001000; // vC= -504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000001; // iC= 1729 
vC = 14'b1111111001011000; // vC= -424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000010; // iC= 1794 
vC = 14'b1111111001011011; // vC= -421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b1111111001100000; // vC= -416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b1111111001111011; // vC= -389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100000; // iC= 1824 
vC = 14'b1111111000111110; // vC= -450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b1111111000110100; // vC= -460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111101; // iC= 1853 
vC = 14'b1111111001101010; // vC= -406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011100; // iC= 1884 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b1111111000101010; // vC= -470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b1111111011000011; // vC= -317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b1111111001010010; // vC= -430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001001; // iC= 1737 
vC = 14'b1111111010111011; // vC= -325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000100; // iC= 1860 
vC = 14'b1111111010000101; // vC= -379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110001; // iC= 1841 
vC = 14'b1111111010001001; // vC= -375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b1111111001100000; // vC= -416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b1111111011010000; // vC= -304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100011; // iC= 1763 
vC = 14'b1111111010011001; // vC= -359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101101; // iC= 1837 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b1111111001100011; // vC= -413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b1111111011011001; // vC= -295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b1111111010011000; // vC= -360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100101; // iC= 1765 
vC = 14'b1111111011101010; // vC= -278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111111001111010; // vC= -390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b1111111010010001; // vC= -367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000001; // iC= 1729 
vC = 14'b1111111011000010; // vC= -318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b1111111011111000; // vC= -264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b1111111010100111; // vC= -345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b1111111010011100; // vC= -356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b1111111011110100; // vC= -268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b1111111011101100; // vC= -276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111111011110111; // vC= -265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b1111111100000000; // vC= -256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101000; // iC= 1832 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b1111111011000010; // vC= -318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000101; // iC= 1861 
vC = 14'b1111111011010001; // vC= -303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b1111111100101101; // vC= -211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111111100011011; // vC= -229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b1111111100000011; // vC= -253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b1111111100010001; // vC= -239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111111100101011; // vC= -213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b1111111100100010; // vC= -222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b1111111101000010; // vC= -190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b1111111100101101; // vC= -211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111110; // iC= 1726 
vC = 14'b1111111110011001; // vC= -103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111001; // iC= 1849 
vC = 14'b1111111100000011; // vC= -253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b1111111101111001; // vC= -135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101110; // iC= 1838 
vC = 14'b1111111101111111; // vC= -129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b1111111100110111; // vC= -201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b1111111110001100; // vC= -116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000100; // iC= 1860 
vC = 14'b1111111101101010; // vC= -150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b1111111110011100; // vC= -100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101110; // iC= 1710 
vC = 14'b1111111110000000; // vC= -128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000100; // iC= 1860 
vC = 14'b1111111101000110; // vC= -186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b1111111110110111; // vC=  -73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010001; // iC= 1745 
vC = 14'b1111111101011110; // vC= -162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b1111111101011100; // vC= -164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b1111111110110011; // vC=  -77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101001; // iC= 1833 
vC = 14'b1111111111001010; // vC=  -54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111111; // iC= 1791 
vC = 14'b1111111111110100; // vC=  -12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001100; // iC= 1740 
vC = 14'b1111111111101111; // vC=  -17 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b1111111110100000; // vC=  -96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b1111111101111101; // vC= -131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b1111111110000100; // vC= -124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b1111111110010110; // vC= -106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b1111111110111111; // vC=  -65 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b1111111111110100; // vC=  -12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110000; // iC= 1840 
vC = 14'b1111111111010111; // vC=  -41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000000000000010; // vC=    2 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b1111111110101011; // vC=  -85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b1111111111111000; // vC=   -8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b1111111110110100; // vC=  -76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011000; // iC= 1752 
vC = 14'b0000000000000011; // vC=    3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b1111111111011100; // vC=  -36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100100; // iC= 1764 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100110; // iC= 1702 
vC = 14'b1111111111000101; // vC=  -59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111111111111000; // vC=   -8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010101; // iC= 1749 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b1111111111110011; // vC=  -13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b0000000001010110; // vC=   86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000000000000011; // vC=    3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100111; // iC= 1703 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b0000000000000110; // vC=    6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b0000000001101111; // vC=  111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010011; // iC= 1747 
vC = 14'b0000000000010111; // vC=   23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110100; // iC= 1780 
vC = 14'b0000000001100000; // vC=   96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110101; // iC= 1781 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000000000111101; // vC=   61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111001; // iC= 1657 
vC = 14'b0000000001111001; // vC=  121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010101; // iC= 1749 
vC = 14'b0000000010010010; // vC=  146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001011; // iC= 1675 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000110; // iC= 1734 
vC = 14'b0000000000110000; // vC=   48 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b0000000010110111; // vC=  183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b0000000000111101; // vC=   61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001110; // iC= 1678 
vC = 14'b0000000011001001; // vC=  201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101100; // iC= 1772 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010101; // iC= 1685 
vC = 14'b0000000011010110; // vC=  214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000000010011100; // vC=  156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011111; // iC= 1759 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100011; // iC= 1699 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101000; // iC= 1640 
vC = 14'b0000000100000101; // vC=  261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b0000000011011001; // vC=  217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111010; // iC= 1658 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b0000000100000100; // vC=  260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111111; // iC= 1663 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b0000000011100110; // vC=  230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b0000000011100000; // vC=  224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b0000000011100011; // vC=  227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101101; // iC= 1709 
vC = 14'b0000000011010011; // vC=  211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100101; // iC= 1637 
vC = 14'b0000000011110111; // vC=  247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100100; // iC= 1636 
vC = 14'b0000000100110111; // vC=  311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110111; // iC= 1655 
vC = 14'b0000000100011001; // vC=  281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b0000000011101100; // vC=  236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100101; // iC= 1637 
vC = 14'b0000000011100111; // vC=  231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b0000000101001011; // vC=  331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111101; // iC= 1597 
vC = 14'b0000000011111111; // vC=  255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111111; // iC= 1599 
vC = 14'b0000000011110010; // vC=  242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010010; // iC= 1618 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011000; // iC= 1624 
vC = 14'b0000000100011000; // vC=  280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100001; // iC= 1633 
vC = 14'b0000000101000011; // vC=  323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010000; // iC= 1616 
vC = 14'b0000000100011111; // vC=  287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b0000000101000000; // vC=  320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000100; // iC= 1604 
vC = 14'b0000000011110101; // vC=  245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011111; // iC= 1695 
vC = 14'b0000000110000111; // vC=  391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b0000000011111011; // vC=  251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000000; // iC= 1600 
vC = 14'b0000000101000011; // vC=  323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b0000000100001011; // vC=  267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100110; // iC= 1638 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b0000000101011011; // vC=  347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101110; // iC= 1646 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110111; // iC= 1655 
vC = 14'b0000000110001001; // vC=  393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b0000000101011011; // vC=  347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b0000000110011001; // vC=  409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110101; // iC= 1653 
vC = 14'b0000000100110001; // vC=  305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011110; // iC= 1630 
vC = 14'b0000000101001101; // vC=  333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b0000000111000001; // vC=  449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100111; // iC= 1575 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001100; // iC= 1612 
vC = 14'b0000000101010111; // vC=  343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010011; // iC= 1555 
vC = 14'b0000000110011100; // vC=  412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010110; // iC= 1686 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101101; // iC= 1581 
vC = 14'b0000000101111110; // vC=  382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001111; // iC= 1551 
vC = 14'b0000000110100011; // vC=  419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001010; // iC= 1610 
vC = 14'b0000000111010110; // vC=  470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b0000001000000100; // vC=  516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111100; // iC= 1596 
vC = 14'b0000000111011010; // vC=  474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010010; // iC= 1618 
vC = 14'b0000001000010011; // vC=  531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000101; // iC= 1605 
vC = 14'b0000000110000011; // vC=  387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111111; // iC= 1663 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100100; // iC= 1572 
vC = 14'b0000000110111010; // vC=  442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000110; // iC= 1542 
vC = 14'b0000001000001001; // vC=  521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011001; // iC= 1625 
vC = 14'b0000000111010001; // vC=  465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001011; // iC= 1547 
vC = 14'b0000001000001010; // vC=  522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b0000000110111000; // vC=  440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111110; // iC= 1534 
vC = 14'b0000001000110111; // vC=  567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100000; // iC= 1632 
vC = 14'b0000001001001000; // vC=  584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001001; // iC= 1545 
vC = 14'b0000000110101110; // vC=  430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001110; // iC= 1550 
vC = 14'b0000000111001011; // vC=  459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b0000000111000100; // vC=  452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001011; // iC= 1547 
vC = 14'b0000000111111111; // vC=  511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110000; // iC= 1520 
vC = 14'b0000000111001001; // vC=  457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001110; // iC= 1486 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000010; // iC= 1538 
vC = 14'b0000001000000111; // vC=  519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110110; // iC= 1526 
vC = 14'b0000001001001101; // vC=  589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001001; // iC= 1609 
vC = 14'b0000001001011101; // vC=  605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101010; // iC= 1578 
vC = 14'b0000001000010111; // vC=  535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111001; // iC= 1529 
vC = 14'b0000001010000000; // vC=  640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b0000000111110101; // vC=  501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000110; // iC= 1478 
vC = 14'b0000001001101000; // vC=  616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110000; // iC= 1584 
vC = 14'b0000001000001110; // vC=  526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001011; // iC= 1547 
vC = 14'b0000001001000110; // vC=  582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110111; // iC= 1591 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101111; // iC= 1455 
vC = 14'b0000001001111001; // vC=  633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111001; // iC= 1529 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110011; // iC= 1523 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011100; // iC= 1436 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010110; // iC= 1494 
vC = 14'b0000001001011011; // vC=  603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010100; // iC= 1492 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010111; // iC= 1431 
vC = 14'b0000001010010110; // vC=  662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000110; // iC= 1478 
vC = 14'b0000001010111001; // vC=  697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110010; // iC= 1458 
vC = 14'b0000001010000101; // vC=  645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010100; // iC= 1556 
vC = 14'b0000001001010111; // vC=  599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000110; // iC= 1414 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111110; // iC= 1534 
vC = 14'b0000001001101110; // vC=  622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110000; // iC= 1456 
vC = 14'b0000001010100010; // vC=  674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011111; // iC= 1439 
vC = 14'b0000001010110001; // vC=  689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101010; // iC= 1450 
vC = 14'b0000001011010110; // vC=  726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000101; // iC= 1413 
vC = 14'b0000001011001001; // vC=  713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010011; // iC= 1427 
vC = 14'b0000001011001100; // vC=  716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100110; // iC= 1510 
vC = 14'b0000001011011000; // vC=  728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011111; // iC= 1503 
vC = 14'b0000001011100100; // vC=  740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010101; // iC= 1429 
vC = 14'b0000001011010100; // vC=  724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010101; // iC= 1493 
vC = 14'b0000001010011011; // vC=  667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000101; // iC= 1477 
vC = 14'b0000001010100011; // vC=  675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111010; // iC= 1402 
vC = 14'b0000001100001100; // vC=  780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010110; // iC= 1494 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001111; // iC= 1423 
vC = 14'b0000001010110001; // vC=  689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001111; // iC= 1487 
vC = 14'b0000001010000101; // vC=  645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101100; // iC= 1516 
vC = 14'b0000001010111101; // vC=  701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000110; // iC= 1478 
vC = 14'b0000001011010111; // vC=  727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000100; // iC= 1412 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111010; // iC= 1402 
vC = 14'b0000001100101010; // vC=  810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010100; // iC= 1364 
vC = 14'b0000001100000111; // vC=  775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000111; // iC= 1479 
vC = 14'b0000001100110001; // vC=  817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000000; // iC= 1472 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001101; // iC= 1485 
vC = 14'b0000001011010011; // vC=  723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110011; // iC= 1331 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110010; // iC= 1330 
vC = 14'b0000001100001100; // vC=  780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101000; // iC= 1448 
vC = 14'b0000001010111110; // vC=  702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101011; // iC= 1387 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b0000001100100101; // vC=  805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001101; // iC= 1421 
vC = 14'b0000001101001101; // vC=  845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111000; // iC= 1464 
vC = 14'b0000001101011000; // vC=  856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110101; // iC= 1461 
vC = 14'b0000001011100100; // vC=  740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100111; // iC= 1447 
vC = 14'b0000001101011101; // vC=  861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010111; // iC= 1367 
vC = 14'b0000001100110010; // vC=  818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001011; // iC= 1291 
vC = 14'b0000001100010001; // vC=  785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101000; // iC= 1384 
vC = 14'b0000001101100100; // vC=  868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110011; // iC= 1395 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110101; // iC= 1333 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011111; // iC= 1375 
vC = 14'b0000001100111100; // vC=  828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110111; // iC= 1335 
vC = 14'b0000001110000000; // vC=  896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010000; // iC= 1424 
vC = 14'b0000001110001100; // vC=  908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101111; // iC= 1327 
vC = 14'b0000001101100100; // vC=  868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111111; // iC= 1343 
vC = 14'b0000001101011001; // vC=  857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111100; // iC= 1340 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100111; // iC= 1255 
vC = 14'b0000001100010001; // vC=  785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111001; // iC= 1337 
vC = 14'b0000001110000010; // vC=  898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001011; // iC= 1355 
vC = 14'b0000001100011000; // vC=  792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011000; // iC= 1304 
vC = 14'b0000001100101100; // vC=  812 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110100; // iC= 1396 
vC = 14'b0000001110000100; // vC=  900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010100; // iC= 1236 
vC = 14'b0000001110101001; // vC=  937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110100; // iC= 1332 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101110; // iC= 1262 
vC = 14'b0000001101010101; // vC=  853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001011; // iC= 1355 
vC = 14'b0000001101101011; // vC=  875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001101; // iC= 1293 
vC = 14'b0000001100100101; // vC=  805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011010; // iC= 1306 
vC = 14'b0000001101010100; // vC=  852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110101; // iC= 1269 
vC = 14'b0000001101111001; // vC=  889 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111001; // iC= 1209 
vC = 14'b0000001101000000; // vC=  832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001001; // iC= 1353 
vC = 14'b0000001101100000; // vC=  864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000001110100110; // vC=  934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000100; // iC= 1220 
vC = 14'b0000001101011010; // vC=  858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111011; // iC= 1339 
vC = 14'b0000001101011100; // vC=  860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000000; // iC= 1344 
vC = 14'b0000001110001111; // vC=  911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010001; // iC= 1297 
vC = 14'b0000001101011110; // vC=  862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110101; // iC= 1205 
vC = 14'b0000001110001110; // vC=  910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110011; // iC= 1267 
vC = 14'b0000001101111110; // vC=  894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010011; // iC= 1235 
vC = 14'b0000001111100001; // vC=  993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011010; // iC= 1306 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100100; // iC= 1252 
vC = 14'b0000001101111010; // vC=  890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010110; // iC= 1302 
vC = 14'b0000001110010110; // vC=  918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101100; // iC= 1260 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100110; // iC= 1254 
vC = 14'b0000001101111000; // vC=  888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100000; // iC= 1184 
vC = 14'b0000001101110101; // vC=  885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111001; // iC= 1145 
vC = 14'b0000001110111010; // vC=  954 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000011; // iC= 1283 
vC = 14'b0000001110111001; // vC=  953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111100; // iC= 1212 
vC = 14'b0000001111000110; // vC=  966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000111; // iC= 1287 
vC = 14'b0000001111100011; // vC=  995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b0000001111110010; // vC= 1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100101; // iC= 1253 
vC = 14'b0000010000001100; // vC= 1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000001111110010; // vC= 1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010000; // iC= 1168 
vC = 14'b0000001111010111; // vC=  983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100011; // iC= 1123 
vC = 14'b0000001111110111; // vC= 1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110001; // iC= 1137 
vC = 14'b0000010000010110; // vC= 1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101000; // iC= 1128 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110101; // iC= 1205 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110000; // iC= 1136 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000111; // iC= 1159 
vC = 14'b0000001111110101; // vC= 1013 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001110; // iC= 1102 
vC = 14'b0000001111011111; // vC=  991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110011; // iC= 1139 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001101; // iC= 1101 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100110; // iC= 1190 
vC = 14'b0000010000111000; // vC= 1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000001; // iC= 1217 
vC = 14'b0000010000011101; // vC= 1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111101; // iC= 1149 
vC = 14'b0000010000100111; // vC= 1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000000; // iC= 1216 
vC = 14'b0000010001000101; // vC= 1093 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101101; // iC= 1069 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000100; // iC= 1092 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001000; // iC= 1160 
vC = 14'b0000010000001101; // vC= 1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100001; // iC= 1185 
vC = 14'b0000010000101111; // vC= 1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101011; // iC= 1067 
vC = 14'b0000010000010000; // vC= 1040 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100100; // iC= 1060 
vC = 14'b0000010001101000; // vC= 1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000011; // iC= 1027 
vC = 14'b0000001111101101; // vC= 1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000110; // iC= 1030 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111010; // iC= 1146 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011100; // iC= 1116 
vC = 14'b0000001111100110; // vC=  998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000110; // iC= 1094 
vC = 14'b0000010001111010; // vC= 1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010101; // iC= 1045 
vC = 14'b0000010000111000; // vC= 1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011010; // iC= 1050 
vC = 14'b0000010001110011; // vC= 1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100111; // iC= 1063 
vC = 14'b0000010000001001; // vC= 1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101101; // iC= 1005 
vC = 14'b0000010001100101; // vC= 1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110100; // iC= 1076 
vC = 14'b0000010001101111; // vC= 1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111101; // iC= 1021 
vC = 14'b0000010001111101; // vC= 1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011011; // iC= 1115 
vC = 14'b0000001111111111; // vC= 1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100001; // iC= 1121 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000100; // iC= 1028 
vC = 14'b0000010010000001; // vC= 1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010000; // iC=  976 
vC = 14'b0000010001010010; // vC= 1106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001000; // iC=  968 
vC = 14'b0000010001011111; // vC= 1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111111; // iC=  959 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101000; // iC= 1000 
vC = 14'b0000010000110011; // vC= 1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000000; // iC=  960 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011111; // iC= 1055 
vC = 14'b0000010001110010; // vC= 1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011000; // iC= 1048 
vC = 14'b0000010010101011; // vC= 1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011011; // iC= 1051 
vC = 14'b0000010010100111; // vC= 1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110111; // iC= 1079 
vC = 14'b0000010001000111; // vC= 1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100101; // iC=  997 
vC = 14'b0000010001000001; // vC= 1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011111; // iC= 1055 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100100; // iC= 1060 
vC = 14'b0000010001101001; // vC= 1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011100; // iC= 1052 
vC = 14'b0000010000111111; // vC= 1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000000; // iC=  960 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001000; // iC= 1032 
vC = 14'b0000010001000000; // vC= 1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001101; // iC= 1037 
vC = 14'b0000010001011010; // vC= 1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000101; // iC=  965 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000101; // iC= 1029 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110011; // iC=  883 
vC = 14'b0000010011011000; // vC= 1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111100; // iC= 1020 
vC = 14'b0000010011010011; // vC= 1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110010; // iC=  946 
vC = 14'b0000010001011110; // vC= 1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000000; // iC= 1024 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110101; // iC= 1013 
vC = 14'b0000010010000100; // vC= 1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101010; // iC=  938 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011011; // iC=  923 
vC = 14'b0000010001010010; // vC= 1106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110011; // iC=  947 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110101; // iC=  885 
vC = 14'b0000010001010101; // vC= 1109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000101; // iC=  965 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000010; // iC=  962 
vC = 14'b0000010010011010; // vC= 1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001110; // iC=  974 
vC = 14'b0000010010110011; // vC= 1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011111; // iC=  863 
vC = 14'b0000010010011010; // vC= 1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010001; // iC=  849 
vC = 14'b0000010011010001; // vC= 1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001100; // iC=  908 
vC = 14'b0000010001111010; // vC= 1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100010; // iC=  930 
vC = 14'b0000010011010010; // vC= 1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010110; // iC=  854 
vC = 14'b0000010011010101; // vC= 1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110011; // iC=  819 
vC = 14'b0000010010010111; // vC= 1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110011; // iC=  819 
vC = 14'b0000010010001100; // vC= 1164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011111; // iC=  927 
vC = 14'b0000010100000110; // vC= 1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101110; // iC=  878 
vC = 14'b0000010011101011; // vC= 1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001010; // iC=  906 
vC = 14'b0000010010110010; // vC= 1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111111; // iC=  895 
vC = 14'b0000010100000111; // vC= 1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011000; // iC=  856 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101111; // iC=  879 
vC = 14'b0000010011100001; // vC= 1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100111; // iC=  871 
vC = 14'b0000010100000101; // vC= 1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111101; // iC=  829 
vC = 14'b0000010100000011; // vC= 1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001101; // iC=  845 
vC = 14'b0000010010111001; // vC= 1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001110; // iC=  782 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011101; // iC=  733 
vC = 14'b0000010100000110; // vC= 1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110001; // iC=  881 
vC = 14'b0000010100100100; // vC= 1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110001; // iC=  881 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101111; // iC=  815 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111001; // iC=  825 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001001; // iC=  777 
vC = 14'b0000010010101111; // vC= 1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011100; // iC=  732 
vC = 14'b0000010011000011; // vC= 1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010011; // iC=  787 
vC = 14'b0000010100111001; // vC= 1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111111; // iC=  831 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010011; // iC=  723 
vC = 14'b0000010100110101; // vC= 1333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110101; // iC=  693 
vC = 14'b0000010011000010; // vC= 1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111100; // iC=  700 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000110; // iC=  774 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011010; // iC=  730 
vC = 14'b0000010100000111; // vC= 1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011101; // iC=  797 
vC = 14'b0000010100100000; // vC= 1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110011; // iC=  755 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010111; // iC=  663 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101001; // iC=  681 
vC = 14'b0000010011000001; // vC= 1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011001; // iC=  665 
vC = 14'b0000010011010000; // vC= 1232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101101; // iC=  749 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001010; // iC=  714 
vC = 14'b0000010011011100; // vC= 1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000000; // iC=  768 
vC = 14'b0000010011001001; // vC= 1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001011; // iC=  715 
vC = 14'b0000010100101011; // vC= 1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101100; // iC=  748 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110101; // iC=  629 
vC = 14'b0000010011100100; // vC= 1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100010; // iC=  674 
vC = 14'b0000010011001001; // vC= 1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001011; // iC=  651 
vC = 14'b0000010011010001; // vC= 1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011001; // iC=  601 
vC = 14'b0000010101001101; // vC= 1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111010; // iC=  698 
vC = 14'b0000010100100000; // vC= 1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111011; // iC=  699 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011110; // iC=  606 
vC = 14'b0000010100100111; // vC= 1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101110; // iC=  622 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111111; // iC=  575 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111111; // iC=  703 
vC = 14'b0000010101101001; // vC= 1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111100; // iC=  700 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110111; // iC=  631 
vC = 14'b0000010100110111; // vC= 1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000101; // iC=  709 
vC = 14'b0000010101001001; // vC= 1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111011; // iC=  699 
vC = 14'b0000010101011110; // vC= 1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111001; // iC=  697 
vC = 14'b0000010100110111; // vC= 1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001111; // iC=  655 
vC = 14'b0000010100000011; // vC= 1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001100; // iC=  652 
vC = 14'b0000010011111001; // vC= 1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110000; // iC=  624 
vC = 14'b0000010101001000; // vC= 1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001101; // iC=  653 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001100; // iC=  588 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110111; // iC=  567 
vC = 14'b0000010101001000; // vC= 1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111000; // iC=  568 
vC = 14'b0000010011100111; // vC= 1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010001; // iC=  657 
vC = 14'b0000010101000000; // vC= 1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100111; // iC=  551 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000010; // iC=  578 
vC = 14'b0000010101101111; // vC= 1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000100; // iC=  580 
vC = 14'b0000010100001101; // vC= 1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110110; // iC=  502 
vC = 14'b0000010101000110; // vC= 1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101101; // iC=  621 
vC = 14'b0000010101001110; // vC= 1358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010101; // iC=  597 
vC = 14'b0000010100010101; // vC= 1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110010; // iC=  626 
vC = 14'b0000010100010111; // vC= 1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100000; // iC=  544 
vC = 14'b0000010101001010; // vC= 1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100111; // iC=  615 
vC = 14'b0000010100001010; // vC= 1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100010; // iC=  610 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001101; // iC=  589 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010001; // iC=  465 
vC = 14'b0000010101001110; // vC= 1358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111110; // iC=  446 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000010; // iC=  450 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111110; // iC=  574 
vC = 14'b0000010100100001; // vC= 1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100010; // iC=  546 
vC = 14'b0000010100010111; // vC= 1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111111; // iC=  575 
vC = 14'b0000010100010111; // vC= 1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000010; // iC=  514 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110001; // iC=  497 
vC = 14'b0000010101011100; // vC= 1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001111; // iC=  527 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110110; // iC=  502 
vC = 14'b0000010100001111; // vC= 1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011100; // iC=  476 
vC = 14'b0000010101001111; // vC= 1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000100; // iC=  452 
vC = 14'b0000010110001111; // vC= 1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101100; // iC=  492 
vC = 14'b0000010101010101; // vC= 1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111110; // iC=  510 
vC = 14'b0000010101010111; // vC= 1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011010; // iC=  474 
vC = 14'b0000010100001010; // vC= 1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000000; // iC=  384 
vC = 14'b0000010110000101; // vC= 1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011101; // iC=  413 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111100; // iC=  444 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010100; // iC=  340 
vC = 14'b0000010101110111; // vC= 1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100010; // iC=  354 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100110; // iC=  358 
vC = 14'b0000010101011000; // vC= 1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100010; // iC=  418 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011010; // iC=  346 
vC = 14'b0000010101111000; // vC= 1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001000; // iC=  328 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101101; // iC=  301 
vC = 14'b0000010100101110; // vC= 1326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110100; // iC=  372 
vC = 14'b0000010100111000; // vC= 1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100100; // iC=  292 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011001; // iC=  281 
vC = 14'b0000010110001101; // vC= 1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100000; // iC=  352 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101000; // iC=  232 
vC = 14'b0000010110011001; // vC= 1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100000; // iC=  288 
vC = 14'b0000010100110101; // vC= 1333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001001; // iC=  329 
vC = 14'b0000010100110010; // vC= 1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101001; // iC=  297 
vC = 14'b0000010101000110; // vC= 1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101001; // iC=  297 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000101; // iC=  261 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100100; // iC=  164 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110011; // iC=  179 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010111; // iC=  215 
vC = 14'b0000010110011001; // vC= 1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111101; // iC=  125 
vC = 14'b0000010101101010; // vC= 1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001111; // iC=  207 
vC = 14'b0000010101101001; // vC= 1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101101; // iC=  173 
vC = 14'b0000010110010001; // vC= 1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000011; // iC=   67 
vC = 14'b0000010100111000; // vC= 1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101010; // iC=  106 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101001; // iC=  169 
vC = 14'b0000010100101010; // vC= 1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011110; // iC=   94 
vC = 14'b0000010110100000; // vC= 1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101111; // iC=   47 
vC = 14'b0000010101001000; // vC= 1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011100; // iC=   28 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110101; // iC=  -11 
vC = 14'b0000010110001100; // vC= 1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101000; // iC=  -24 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110111; // iC=   -9 
vC = 14'b0000010110000100; // vC= 1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010100; // iC=  -44 
vC = 14'b0000010101011000; // vC= 1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110010; // iC=  -14 
vC = 14'b0000010110001010; // vC= 1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100110; // iC=  -26 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000011; // iC=    3 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011101; // iC=  -99 
vC = 14'b0000010100001110; // vC= 1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010101; // iC=  -43 
vC = 14'b0000010100111101; // vC= 1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110000; // iC=  -80 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101011; // iC=  -85 
vC = 14'b0000010100010100; // vC= 1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111000; // iC= -136 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000100; // iC= -124 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000100; // iC= -188 
vC = 14'b0000010110100000; // vC= 1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010111; // iC= -169 
vC = 14'b0000010101001001; // vC= 1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010001; // iC= -303 
vC = 14'b0000010101111000; // vC= 1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011010; // iC= -294 
vC = 14'b0000010100100011; // vC= 1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110000; // iC= -208 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011110; // iC= -354 
vC = 14'b0000010100000001; // vC= 1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111100; // iC= -260 
vC = 14'b0000010101111100; // vC= 1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011000; // iC= -424 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110111; // iC= -329 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000110; // iC= -378 
vC = 14'b0000010101011010; // vC= 1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100111; // iC= -345 
vC = 14'b0000010101110001; // vC= 1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011111; // iC= -417 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100100; // iC= -412 
vC = 14'b0000010100100000; // vC= 1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100100; // iC= -540 
vC = 14'b0000010101001101; // vC= 1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001001; // iC= -439 
vC = 14'b0000010101000100; // vC= 1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101100; // iC= -468 
vC = 14'b0000010011111011; // vC= 1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110011; // iC= -589 
vC = 14'b0000010101011001; // vC= 1369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b0000010110000001; // vC= 1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101100; // iC= -596 
vC = 14'b0000010100101011; // vC= 1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010100; // iC= -684 
vC = 14'b0000010100000011; // vC= 1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101011; // iC= -597 
vC = 14'b0000010100010111; // vC= 1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110101; // iC= -651 
vC = 14'b0000010011111000; // vC= 1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110010; // iC= -718 
vC = 14'b0000010101110101; // vC= 1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001011; // iC= -693 
vC = 14'b0000010011010110; // vC= 1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011111; // iC= -673 
vC = 14'b0000010011011010; // vC= 1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101110; // iC= -786 
vC = 14'b0000010100011100; // vC= 1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101000; // iC= -792 
vC = 14'b0000010100001110; // vC= 1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001110; // iC= -818 
vC = 14'b0000010011011000; // vC= 1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000000; // iC= -832 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110100; // iC= -844 
vC = 14'b0000010011000011; // vC= 1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101101; // iC= -787 
vC = 14'b0000010100010111; // vC= 1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100001; // iC= -927 
vC = 14'b0000010100110001; // vC= 1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000000; // iC= -896 
vC = 14'b0000010011010011; // vC= 1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010001; // iC= -815 
vC = 14'b0000010100001101; // vC= 1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111011; // iC= -965 
vC = 14'b0000010010110101; // vC= 1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011101; // iC= -931 
vC = 14'b0000010100000010; // vC= 1282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101110; // iC= -978 
vC = 14'b0000010011110010; // vC= 1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100100; // iC= -924 
vC = 14'b0000010010101111; // vC= 1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100110; // iC= -986 
vC = 14'b0000010100001000; // vC= 1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001001; // iC=-1015 
vC = 14'b0000010011111100; // vC= 1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010110; // iC= -938 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010000; // iC=-1008 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101100; // iC=-1044 
vC = 14'b0000010011011010; // vC= 1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010010; // iC=-1134 
vC = 14'b0000010100010011; // vC= 1299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011011; // iC=-1061 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100101; // iC=-1051 
vC = 14'b0000010010001111; // vC= 1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011111; // iC=-1185 
vC = 14'b0000010011001011; // vC= 1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101011; // iC=-1109 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001001; // iC=-1143 
vC = 14'b0000010011010111; // vC= 1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011110; // iC=-1186 
vC = 14'b0000010011101010; // vC= 1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111011; // iC=-1221 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011010; // iC=-1190 
vC = 14'b0000010100000011; // vC= 1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011110; // iC=-1122 
vC = 14'b0000010011001010; // vC= 1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110101; // iC=-1163 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011011; // iC=-1253 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100111; // iC=-1305 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001101; // iC=-1267 
vC = 14'b0000010011001101; // vC= 1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101000; // iC=-1240 
vC = 14'b0000010011000111; // vC= 1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110010; // iC=-1230 
vC = 14'b0000010011001001; // vC= 1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b0000010010010011; // vC= 1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110001; // iC=-1295 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111110; // iC=-1282 
vC = 14'b0000010010000010; // vC= 1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010111; // iC=-1385 
vC = 14'b0000010000111010; // vC= 1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000000; // iC=-1280 
vC = 14'b0000010001100001; // vC= 1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110011; // iC=-1293 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101010; // iC=-1366 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b0000010001011001; // vC= 1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001101; // iC=-1395 
vC = 14'b0000010001111000; // vC= 1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111000; // iC=-1416 
vC = 14'b0000010010001101; // vC= 1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b0000010000000010; // vC= 1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b0000010001101110; // vC= 1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000100; // iC=-1468 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b0000010000101010; // vC= 1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b0000001111101011; // vC= 1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b0000010000001010; // vC= 1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b0000001111011010; // vC=  986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100110; // iC=-1562 
vC = 14'b0000010000111101; // vC= 1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011111; // iC=-1505 
vC = 14'b0000010000000001; // vC= 1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001101; // iC=-1587 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b0000010000110100; // vC= 1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b0000001111000101; // vC=  965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b0000010000110111; // vC= 1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011111; // iC=-1505 
vC = 14'b0000010000100111; // vC= 1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b0000010000110110; // vC= 1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b0000001110010100; // vC=  916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b0000001111011111; // vC=  991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b0000001110110011; // vC=  947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b0000001111111001; // vC= 1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000001111010000; // vC=  976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001101; // iC=-1587 
vC = 14'b0000001110111011; // vC=  955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111001; // iC=-1607 
vC = 14'b0000001111000110; // vC=  966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b0000001110101010; // vC=  938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000001111100001; // vC=  993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b0000001101111110; // vC=  894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b0000001101000101; // vC=  837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111100; // iC=-1540 
vC = 14'b0000001111010111; // vC=  983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b0000001111010101; // vC=  981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000001101100001; // vC=  865 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111101; // iC=-1667 
vC = 14'b0000001101110101; // vC=  885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000001; // iC=-1663 
vC = 14'b0000001101010101; // vC=  853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010010; // iC=-1646 
vC = 14'b0000001110001100; // vC=  908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111010; // iC=-1670 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b0000001101111100; // vC=  892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110001; // iC=-1615 
vC = 14'b0000001100001110; // vC=  782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000001110001010; // vC=  906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111001; // iC=-1607 
vC = 14'b0000001101011000; // vC=  856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101100; // iC=-1556 
vC = 14'b0000001101011111; // vC=  863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b0000001101100110; // vC=  870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b0000001011111111; // vC=  767 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101000; // iC=-1688 
vC = 14'b0000001101111011; // vC=  891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b0000001100011100; // vC=  796 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b0000001100001000; // vC=  776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110100; // iC=-1548 
vC = 14'b0000001101100010; // vC=  866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000001; // iC=-1599 
vC = 14'b0000001011110000; // vC=  752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b0000001101001011; // vC=  843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111100; // iC=-1604 
vC = 14'b0000001100000100; // vC=  772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110100; // iC=-1548 
vC = 14'b0000001101001101; // vC=  845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000001011101100; // vC=  748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101101; // iC=-1555 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b0000001011100001; // vC=  737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111010; // iC=-1670 
vC = 14'b0000001011000001; // vC=  705 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100100; // iC=-1564 
vC = 14'b0000001100000001; // vC=  769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b0000001100011111; // vC=  799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b0000001010011000; // vC=  664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b0000001010100000; // vC=  672 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000001011111001; // vC=  761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b0000001011011110; // vC=  734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100011; // iC=-1565 
vC = 14'b0000001011010001; // vC=  721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001101; // iC=-1651 
vC = 14'b0000001011000111; // vC=  711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000001011011101; // vC=  733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b0000001001001110; // vC=  590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b0000001011000101; // vC=  709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b0000001001111000; // vC=  632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b0000001010101100; // vC=  684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001101; // iC=-1651 
vC = 14'b0000001000011110; // vC=  542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b0000001000110000; // vC=  560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000001000101011; // vC=  555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b0000001000110111; // vC=  567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b0000001001111011; // vC=  635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000001001100000; // vC=  608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b0000001000000101; // vC=  517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100101; // iC=-1627 
vC = 14'b0000000111111110; // vC=  510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101110; // iC=-1618 
vC = 14'b0000001001100101; // vC=  613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011110; // iC=-1634 
vC = 14'b0000001000101010; // vC=  554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b0000001001110000; // vC=  624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110111; // iC=-1673 
vC = 14'b0000000111111100; // vC=  508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000111; // iC=-1657 
vC = 14'b0000000111100010; // vC=  482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000001000100100; // vC=  548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b0000001000011110; // vC=  542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b0000001000101010; // vC=  554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b0000001000000100; // vC=  516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000001000101110; // vC=  558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000001; // iC=-1663 
vC = 14'b0000000111100010; // vC=  482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110001; // iC=-1679 
vC = 14'b0000000111110001; // vC=  497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000000110010110; // vC=  406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b0000000111111111; // vC=  511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000001000010000; // vC=  528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001110; // iC=-1586 
vC = 14'b0000000110001111; // vC=  399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110111; // iC=-1609 
vC = 14'b0000000110011000; // vC=  408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b0000000110101101; // vC=  429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011101; // iC=-1699 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b0000000110001000; // vC=  392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b0000000110001000; // vC=  392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000000111101000; // vC=  488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b0000000110100110; // vC=  422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b0000000110110011; // vC=  435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b0000000110011100; // vC=  412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111101; // iC=-1667 
vC = 14'b0000000101011001; // vC=  345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b0000000110001001; // vC=  393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b0000000111000010; // vC=  450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000000100111101; // vC=  317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b0000000101100001; // vC=  353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111111; // iC=-1665 
vC = 14'b0000000101010110; // vC=  342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000010; // iC=-1662 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110110; // iC=-1674 
vC = 14'b0000000100111010; // vC=  314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b0000000100100101; // vC=  293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b0000000100111100; // vC=  316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b0000000101001111; // vC=  335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b0000000101000011; // vC=  323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010111; // iC=-1641 
vC = 14'b0000000101011001; // vC=  345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011010; // iC=-1702 
vC = 14'b0000000100110101; // vC=  309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111010; // iC=-1670 
vC = 14'b0000000100010101; // vC=  277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110111; // iC=-1673 
vC = 14'b0000000101000100; // vC=  324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b0000000011100100; // vC=  228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b0000000101000100; // vC=  324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000000101001011; // vC=  331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b0000000100110000; // vC=  304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b0000000010101110; // vC=  174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101000; // iC=-1688 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b0000000100011010; // vC=  282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b0000000100011111; // vC=  287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b0000000011001011; // vC=  203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b0000000100100010; // vC=  290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011110; // iC=-1634 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b0000000011110010; // vC=  242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b0000000100001011; // vC=  267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111100; // iC=-1668 
vC = 14'b0000000011111010; // vC=  250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b0000000011101000; // vC=  232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b0000000010000101; // vC=  133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101010; // iC=-1558 
vC = 14'b0000000011100101; // vC=  229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b0000000010100010; // vC=  162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b0000000010111011; // vC=  187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010111; // iC=-1577 
vC = 14'b0000000011001001; // vC=  201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b0000000010010010; // vC=  146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000000011000111; // vC=  199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b0000000000111111; // vC=   63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b0000000010011011; // vC=  155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b0000000000111001; // vC=   57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000000010010010; // vC=  146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110000; // iC=-1552 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110110; // iC=-1674 
vC = 14'b0000000000011000; // vC=   24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b0000000001011110; // vC=   94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b0000000001011110; // vC=   94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b0000000001000100; // vC=   68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b0000000000111101; // vC=   61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000000000100010; // vC=   34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b0000000001011100; // vC=   92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b0000000001110111; // vC=  119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b0000000001011111; // vC=   95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b0000000000001111; // vC=   15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000000000000101; // vC=    5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110001; // iC=-1679 
vC = 14'b0000000001011111; // vC=   95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b1111111111011100; // vC=  -36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000000001000101; // vC=   69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b1111111111000010; // vC=  -62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b0000000000010001; // vC=   17 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001000; // iC=-1656 
vC = 14'b1111111111111100; // vC=   -4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100000; // iC=-1632 
vC = 14'b1111111111110111; // vC=   -9 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b1111111111100011; // vC=  -29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b0000000000000110; // vC=    6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b1111111110011010; // vC= -102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100011; // iC=-1565 
vC = 14'b0000000000010011; // vC=   19 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b0000000000001010; // vC=   10 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001100; // iC=-1524 
vC = 14'b1111111110100011; // vC=  -93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010001; // iC=-1583 
vC = 14'b1111111110001110; // vC= -114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000111; // iC=-1657 
vC = 14'b0000000000000010; // vC=    2 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100011; // iC=-1629 
vC = 14'b1111111110101101; // vC=  -83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b1111111111011111; // vC=  -33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b1111111101101111; // vC= -145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010001; // iC=-1583 
vC = 14'b1111111111101111; // vC=  -17 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b1111111110000001; // vC= -127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b1111111111010001; // vC=  -47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b1111111110110011; // vC=  -77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b1111111111010110; // vC=  -42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b1111111111010010; // vC=  -46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b1111111110001010; // vC= -118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b1111111101110010; // vC= -142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b1111111101001001; // vC= -183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b1111111110011101; // vC=  -99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b1111111100101110; // vC= -210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b1111111101100010; // vC= -158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010111; // iC=-1577 
vC = 14'b1111111101001010; // vC= -182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b1111111110001010; // vC= -118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101101; // iC=-1619 
vC = 14'b1111111100001000; // vC= -248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b1111111101000011; // vC= -189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111001; // iC=-1479 
vC = 14'b1111111100100110; // vC= -218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b1111111011110100; // vC= -268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001110; // iC=-1586 
vC = 14'b1111111011110001; // vC= -271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b1111111100101110; // vC= -210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111100; // iC=-1540 
vC = 14'b1111111100000111; // vC= -249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b1111111011100011; // vC= -285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b1111111101101001; // vC= -151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b1111111101001111; // vC= -177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100110; // iC=-1562 
vC = 14'b1111111100101101; // vC= -211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b1111111100010110; // vC= -234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b1111111011011100; // vC= -292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b1111111100100110; // vC= -218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b1111111100010011; // vC= -237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010011; // iC=-1581 
vC = 14'b1111111011101100; // vC= -276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011001; // iC=-1447 
vC = 14'b1111111100011001; // vC= -231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b1111111100011001; // vC= -231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b1111111100001111; // vC= -241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b1111111100101101; // vC= -211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b1111111100000100; // vC= -252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b1111111011011001; // vC= -295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b1111111011011111; // vC= -289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011001; // iC=-1447 
vC = 14'b1111111011111001; // vC= -263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101000; // iC=-1432 
vC = 14'b1111111100010111; // vC= -233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b1111111011111111; // vC= -257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b1111111001101110; // vC= -402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111101; // iC=-1475 
vC = 14'b1111111011100000; // vC= -288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000011; // iC=-1533 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111100; // iC=-1476 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b1111111010110001; // vC= -335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b1111111010110000; // vC= -336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b1111111010110100; // vC= -332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010100; // iC=-1388 
vC = 14'b1111111010011101; // vC= -355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b1111111001001010; // vC= -438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b1111111001001110; // vC= -434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b1111111001111001; // vC= -391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b1111111010000101; // vC= -379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101000; // iC=-1432 
vC = 14'b1111111010000110; // vC= -378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b1111111000100100; // vC= -476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101101; // iC=-1491 
vC = 14'b1111111010000100; // vC= -380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101011; // iC=-1429 
vC = 14'b1111111000110000; // vC= -464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110001; // iC=-1487 
vC = 14'b1111111010100110; // vC= -346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100101; // iC=-1371 
vC = 14'b1111111001110100; // vC= -396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b1111111000000011; // vC= -509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b1111111001001111; // vC= -433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b1111111000010011; // vC= -493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010001; // iC=-1455 
vC = 14'b1111111010000111; // vC= -377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110110; // iC=-1354 
vC = 14'b1111111001101100; // vC= -404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101011; // iC=-1365 
vC = 14'b1111111001101101; // vC= -403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101110; // iC=-1362 
vC = 14'b1111111000011001; // vC= -487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001101; // iC=-1459 
vC = 14'b1111111001110100; // vC= -396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001101; // iC=-1395 
vC = 14'b1111110111010011; // vC= -557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001011; // iC=-1333 
vC = 14'b1111111001101001; // vC= -407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001011; // iC=-1397 
vC = 14'b1111111000100101; // vC= -475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b1111111000010101; // vC= -491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011011; // iC=-1445 
vC = 14'b1111110111101100; // vC= -532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111010; // iC=-1414 
vC = 14'b1111111000100010; // vC= -478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001100; // iC=-1332 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110100; // iC=-1356 
vC = 14'b1111110111000010; // vC= -574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011100; // iC=-1316 
vC = 14'b1111110111111101; // vC= -515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110000; // iC=-1360 
vC = 14'b1111111001000010; // vC= -446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100101; // iC=-1435 
vC = 14'b1111111000101101; // vC= -467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100001; // iC=-1375 
vC = 14'b1111110111110010; // vC= -526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010111; // iC=-1321 
vC = 14'b1111110111100110; // vC= -538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111100; // iC=-1348 
vC = 14'b1111110111000011; // vC= -573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101010; // iC=-1430 
vC = 14'b1111110111010010; // vC= -558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b1111110110101100; // vC= -596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110000; // iC=-1296 
vC = 14'b1111110110001010; // vC= -630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110101; // iC=-1291 
vC = 14'b1111110111100101; // vC= -539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111101; // iC=-1347 
vC = 14'b1111110110101100; // vC= -596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001101; // iC=-1395 
vC = 14'b1111110110011100; // vC= -612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101011; // iC=-1429 
vC = 14'b1111110111001101; // vC= -563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110100; // iC=-1356 
vC = 14'b1111110110001010; // vC= -630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111100; // iC=-1348 
vC = 14'b1111110111111110; // vC= -514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010101; // iC=-1387 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010100; // iC=-1324 
vC = 14'b1111110110010111; // vC= -617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000000; // iC=-1344 
vC = 14'b1111110111001011; // vC= -565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000111; // iC=-1337 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b1111110110010001; // vC= -623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101001; // iC=-1239 
vC = 14'b1111110110011001; // vC= -615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001111; // iC=-1393 
vC = 14'b1111110101010001; // vC= -687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010000; // iC=-1264 
vC = 14'b1111110101101010; // vC= -662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110011; // iC=-1357 
vC = 14'b1111110110000111; // vC= -633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110101; // iC=-1291 
vC = 14'b1111110101001111; // vC= -689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b1111110101100011; // vC= -669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100110; // iC=-1242 
vC = 14'b1111110101011111; // vC= -673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011001; // iC=-1255 
vC = 14'b1111110101111111; // vC= -641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101011; // iC=-1301 
vC = 14'b1111110100100000; // vC= -736 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101111; // iC=-1233 
vC = 14'b1111110110000110; // vC= -634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000011; // iC=-1213 
vC = 14'b1111110110011100; // vC= -612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110111; // iC=-1353 
vC = 14'b1111110100101110; // vC= -722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010110; // iC=-1194 
vC = 14'b1111110100100011; // vC= -733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000100; // iC=-1212 
vC = 14'b1111110101110100; // vC= -652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b1111110100110001; // vC= -719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000000; // iC=-1280 
vC = 14'b1111110011110100; // vC= -780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110011; // iC=-1293 
vC = 14'b1111110110000001; // vC= -639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111001; // iC=-1223 
vC = 14'b1111110100100101; // vC= -731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111011; // iC=-1285 
vC = 14'b1111110011110110; // vC= -778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001011; // iC=-1269 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011101; // iC=-1187 
vC = 14'b1111110100111010; // vC= -710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110001; // iC=-1231 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111011; // iC=-1285 
vC = 14'b1111110011010001; // vC= -815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100010; // iC=-1310 
vC = 14'b1111110011111011; // vC= -773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001000; // iC=-1144 
vC = 14'b1111110100001110; // vC= -754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101110; // iC=-1298 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011011; // iC=-1189 
vC = 14'b1111110100110011; // vC= -717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110100; // iC=-1164 
vC = 14'b1111110101010010; // vC= -686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011101; // iC=-1123 
vC = 14'b1111110101001101; // vC= -691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110110; // iC=-1162 
vC = 14'b1111110101001010; // vC= -694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101111; // iC=-1169 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110000; // iC=-1168 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100011; // iC=-1181 
vC = 14'b1111110010111010; // vC= -838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000001; // iC=-1151 
vC = 14'b1111110011010110; // vC= -810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101100; // iC=-1172 
vC = 14'b1111110011111110; // vC= -770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101000; // iC=-1112 
vC = 14'b1111110100101000; // vC= -728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010001; // iC=-1199 
vC = 14'b1111110011001110; // vC= -818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100110; // iC=-1242 
vC = 14'b1111110010110101; // vC= -843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111010; // iC=-1094 
vC = 14'b1111110100000110; // vC= -762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111110; // iC=-1090 
vC = 14'b1111110011111110; // vC= -770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101100; // iC=-1108 
vC = 14'b1111110010011110; // vC= -866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011100; // iC=-1124 
vC = 14'b1111110100000010; // vC= -766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010000; // iC=-1136 
vC = 14'b1111110011100111; // vC= -793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101010; // iC=-1110 
vC = 14'b1111110010110110; // vC= -842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011110; // iC=-1186 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010101; // iC=-1067 
vC = 14'b1111110011000000; // vC= -832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001001; // iC=-1143 
vC = 14'b1111110001111110; // vC= -898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101000; // iC=-1112 
vC = 14'b1111110011010001; // vC= -815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100001; // iC=-1055 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001110; // iC=-1202 
vC = 14'b1111110010111100; // vC= -836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111111; // iC=-1153 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110010; // iC=-1038 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101101; // iC=-1043 
vC = 14'b1111110001001101; // vC= -947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100111; // iC=-1113 
vC = 14'b1111110010000111; // vC= -889 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101110; // iC=-1042 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011111; // iC=-1121 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000101; // iC=-1147 
vC = 14'b1111110001111111; // vC= -897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000110; // iC=-1018 
vC = 14'b1111110011010110; // vC= -810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111101; // iC=-1091 
vC = 14'b1111110001101101; // vC= -915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010100; // iC=-1132 
vC = 14'b1111110010101101; // vC= -851 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011100; // iC= -996 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110010; // iC=-1102 
vC = 14'b1111110000101110; // vC= -978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001011; // iC=-1141 
vC = 14'b1111110010010111; // vC= -873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110011; // iC=-1101 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110000; // iC=-1104 
vC = 14'b1111110010010010; // vC= -878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011000; // iC=-1128 
vC = 14'b1111110010000100; // vC= -892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011101; // iC= -995 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011010; // iC=-1126 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101110; // iC= -978 
vC = 14'b1111110000101010; // vC= -982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110010; // iC=-1038 
vC = 14'b1111110000011000; // vC=-1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101100; // iC= -980 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101110; // iC= -978 
vC = 14'b1111110010001000; // vC= -888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010000; // iC=-1072 
vC = 14'b1111110001001010; // vC= -950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101011; // iC=-1045 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111001; // iC=-1031 
vC = 14'b1111110001000000; // vC= -960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111110001001000; // vC= -952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100101; // iC= -923 
vC = 14'b1111101111111111; // vC=-1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100111; // iC=-1049 
vC = 14'b1111101111110100; // vC=-1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100001; // iC= -991 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011000; // iC=-1000 
vC = 14'b1111110001001000; // vC= -952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101111; // iC=-1041 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001110; // iC= -946 
vC = 14'b1111110001011001; // vC= -935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010100; // iC= -940 
vC = 14'b1111110000000100; // vC=-1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001010; // iC= -950 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101100; // iC= -916 
vC = 14'b1111110001101010; // vC= -918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111000; // iC=-1032 
vC = 14'b1111110000100011; // vC= -989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111100; // iC= -964 
vC = 14'b1111101111100000; // vC=-1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100101; // iC= -923 
vC = 14'b1111110001001110; // vC= -946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001101; // iC= -947 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011100; // iC= -996 
vC = 14'b1111110000011110; // vC= -994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100001; // iC= -863 
vC = 14'b1111110001010111; // vC= -937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011001; // iC= -935 
vC = 14'b1111101110111101; // vC=-1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010100; // iC=-1004 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010001; // iC= -879 
vC = 14'b1111110000011010; // vC= -998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100000; // iC= -864 
vC = 14'b1111101111111001; // vC=-1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010110; // iC= -938 
vC = 14'b1111101111011101; // vC=-1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111111; // iC= -961 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100000; // iC= -992 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100101; // iC= -987 
vC = 14'b1111101110011100; // vC=-1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100111; // iC= -857 
vC = 14'b1111101111011100; // vC=-1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111001; // iC= -839 
vC = 14'b1111101111011001; // vC=-1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010010; // iC= -814 
vC = 14'b1111101110111101; // vC=-1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111011; // iC= -965 
vC = 14'b1111101110101111; // vC=-1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100101; // iC= -923 
vC = 14'b1111110000101001; // vC= -983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100011; // iC= -861 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011000; // iC= -936 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101000; // iC= -856 
vC = 14'b1111101111110111; // vC=-1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101100; // iC= -852 
vC = 14'b1111101111010100; // vC=-1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010011; // iC= -813 
vC = 14'b1111101110111110; // vC=-1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011101; // iC= -931 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111001; // iC= -839 
vC = 14'b1111101110100111; // vC=-1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100001; // iC= -927 
vC = 14'b1111101111011100; // vC=-1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000000; // iC= -896 
vC = 14'b1111101110001110; // vC=-1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101110; // iC= -850 
vC = 14'b1111101110011011; // vC=-1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101100; // iC= -852 
vC = 14'b1111101110000011; // vC=-1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101111; // iC= -849 
vC = 14'b1111101110000000; // vC=-1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101100; // iC= -852 
vC = 14'b1111101110101111; // vC=-1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100100; // iC= -860 
vC = 14'b1111101110111100; // vC=-1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010011; // iC= -813 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111110; // iC= -770 
vC = 14'b1111101110110101; // vC=-1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011100; // iC= -740 
vC = 14'b1111101110000001; // vC=-1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001010; // iC= -822 
vC = 14'b1111101110000110; // vC=-1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101110; // iC= -722 
vC = 14'b1111101111001110; // vC=-1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100110; // iC= -794 
vC = 14'b1111101111100111; // vC=-1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110000; // iC= -848 
vC = 14'b1111101111010111; // vC=-1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000100; // iC= -764 
vC = 14'b1111101110100110; // vC=-1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111110; // iC= -770 
vC = 14'b1111101110011100; // vC=-1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010110; // iC= -746 
vC = 14'b1111101101110100; // vC=-1164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010000; // iC= -816 
vC = 14'b1111101111011100; // vC=-1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101110; // iC= -722 
vC = 14'b1111101101110101; // vC=-1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011100; // iC= -740 
vC = 14'b1111101110010000; // vC=-1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001000; // iC= -760 
vC = 14'b1111101100111011; // vC=-1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010000; // iC= -688 
vC = 14'b1111101101101001; // vC=-1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100010; // iC= -798 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010001; // iC= -751 
vC = 14'b1111101110101011; // vC=-1109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101000; // iC= -728 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111101110001000; // vC=-1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110000; // iC= -656 
vC = 14'b1111101101111000; // vC=-1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110101; // iC= -715 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100110; // iC= -730 
vC = 14'b1111101110001011; // vC=-1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010010; // iC= -686 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101011; // iC= -725 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101101; // iC= -723 
vC = 14'b1111101101111000; // vC=-1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110001; // iC= -655 
vC = 14'b1111101100110111; // vC=-1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101000; // iC= -664 
vC = 14'b1111101110001010; // vC=-1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111000; // iC= -648 
vC = 14'b1111101101100000; // vC=-1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101001; // iC= -663 
vC = 14'b1111101101100110; // vC=-1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001000; // iC= -696 
vC = 14'b1111101100010110; // vC=-1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011011; // iC= -677 
vC = 14'b1111101110001011; // vC=-1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111000; // iC= -584 
vC = 14'b1111101101000010; // vC=-1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111101; // iC= -707 
vC = 14'b1111101110010111; // vC=-1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011010; // iC= -678 
vC = 14'b1111101100111100; // vC=-1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011001; // iC= -615 
vC = 14'b1111101100111000; // vC=-1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101011; // iC= -597 
vC = 14'b1111101101101001; // vC=-1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111101101101110; // vC=-1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110101; // iC= -651 
vC = 14'b1111101101101011; // vC=-1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101001; // iC= -599 
vC = 14'b1111101100010001; // vC=-1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101011; // iC= -661 
vC = 14'b1111101100111110; // vC=-1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011001; // iC= -615 
vC = 14'b1111101100100101; // vC=-1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100001; // iC= -607 
vC = 14'b1111101011111111; // vC=-1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000101; // iC= -635 
vC = 14'b1111101100101011; // vC=-1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001101; // iC= -627 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000101; // iC= -571 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110010; // iC= -654 
vC = 14'b1111101110001010; // vC=-1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110011; // iC= -653 
vC = 14'b1111101100001110; // vC=-1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001101; // iC= -499 
vC = 14'b1111101101100110; // vC=-1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111001; // iC= -583 
vC = 14'b1111101100101111; // vC=-1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111010; // iC= -518 
vC = 14'b1111101100011101; // vC=-1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010001; // iC= -623 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101110; // iC= -530 
vC = 14'b1111101101010000; // vC=-1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100101; // iC= -475 
vC = 14'b1111101101100111; // vC=-1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b1111101101010011; // vC=-1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010110; // iC= -554 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011001; // iC= -551 
vC = 14'b1111101011011100; // vC=-1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101010; // iC= -534 
vC = 14'b1111101100000111; // vC=-1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111101101100111; // vC=-1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111011; // iC= -581 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110101; // iC= -459 
vC = 14'b1111101011011000; // vC=-1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100101; // iC= -539 
vC = 14'b1111101011110011; // vC=-1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110011; // iC= -461 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110011; // iC= -525 
vC = 14'b1111101100001000; // vC=-1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001101; // iC= -499 
vC = 14'b1111101011100111; // vC=-1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111000; // iC= -456 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100000; // iC= -416 
vC = 14'b1111101100010100; // vC=-1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111010; // iC= -454 
vC = 14'b1111101101011101; // vC=-1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100011; // iC= -413 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111001; // iC= -519 
vC = 14'b1111101100001010; // vC=-1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011011; // iC= -485 
vC = 14'b1111101101001001; // vC=-1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111100; // iC= -516 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101011; // iC= -533 
vC = 14'b1111101011110100; // vC=-1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011011; // iC= -421 
vC = 14'b1111101101010000; // vC=-1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110101; // iC= -459 
vC = 14'b1111101011100011; // vC=-1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000010; // iC= -382 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010001; // iC= -431 
vC = 14'b1111101100000011; // vC=-1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010111; // iC= -489 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101111; // iC= -401 
vC = 14'b1111101011001100; // vC=-1332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110110; // iC= -394 
vC = 14'b1111101100111000; // vC=-1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011011; // iC= -421 
vC = 14'b1111101011111001; // vC=-1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110111; // iC= -329 
vC = 14'b1111101011010101; // vC=-1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100001; // iC= -479 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010100; // iC= -428 
vC = 14'b1111101100011111; // vC=-1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111011; // iC= -325 
vC = 14'b1111101100110000; // vC=-1232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110010; // iC= -462 
vC = 14'b1111101011101101; // vC=-1299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111010; // iC= -390 
vC = 14'b1111101011010101; // vC=-1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000000; // iC= -384 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100011; // iC= -285 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110000; // iC= -400 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011000; // iC= -296 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011101; // iC= -291 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111101; // iC= -259 
vC = 14'b1111101100010000; // vC=-1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011011; // iC= -229 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100111; // iC= -281 
vC = 14'b1111101010110001; // vC=-1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111001; // iC= -327 
vC = 14'b1111101100010000; // vC=-1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001001; // iC= -311 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100001; // iC= -223 
vC = 14'b1111101011101001; // vC=-1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010010; // iC= -302 
vC = 14'b1111101100100011; // vC=-1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000001; // iC= -255 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000111; // iC= -185 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001100; // iC= -116 
vC = 14'b1111101100101001; // vC=-1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011001; // iC= -167 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010101; // iC= -107 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111100; // iC= -196 
vC = 14'b1111101011001101; // vC=-1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011010; // iC= -166 
vC = 14'b1111101100101000; // vC=-1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000101; // iC= -187 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100000; // iC= -160 
vC = 14'b1111101010011010; // vC=-1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010000; // iC= -112 
vC = 14'b1111101100000011; // vC=-1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111101; // iC=   -3 
vC = 14'b1111101100101011; // vC=-1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001111; // iC=  -49 
vC = 14'b1111101100100010; // vC=-1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110100; // iC=  -76 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011010; // iC=   26 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010100; // iC=   20 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111000; // iC=   56 
vC = 14'b1111101011110000; // vC=-1296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000111; // iC=    7 
vC = 14'b1111101100010110; // vC=-1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111001; // iC=   -7 
vC = 14'b1111101100001110; // vC=-1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010101; // iC=   21 
vC = 14'b1111101010110101; // vC=-1355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111000; // iC=  120 
vC = 14'b1111101100100101; // vC=-1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111011; // iC=  123 
vC = 14'b1111101011001001; // vC=-1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010100; // iC=  148 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111000; // iC=  184 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001001; // iC=  137 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101101; // iC=  109 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000000; // iC=  128 
vC = 14'b1111101011110010; // vC=-1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110010; // iC=  242 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100011; // iC=  163 
vC = 14'b1111101011010001; // vC=-1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100101; // iC=  229 
vC = 14'b1111101100001111; // vC=-1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100000; // iC=  224 
vC = 14'b1111101011010000; // vC=-1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100000; // iC=  288 
vC = 14'b1111101011011110; // vC=-1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011110; // iC=  286 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110011; // iC=  243 
vC = 14'b1111101011000101; // vC=-1339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010111; // iC=  407 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110110; // iC=  438 
vC = 14'b1111101100111010; // vC=-1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001001; // iC=  393 
vC = 14'b1111101011110010; // vC=-1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101011; // iC=  427 
vC = 14'b1111101100100011; // vC=-1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100110; // iC=  358 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111101; // iC=  381 
vC = 14'b1111101100001000; // vC=-1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101010; // iC=  426 
vC = 14'b1111101100101111; // vC=-1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001110; // iC=  462 
vC = 14'b1111101011001101; // vC=-1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000001; // iC=  449 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010110; // iC=  598 
vC = 14'b1111101011111100; // vC=-1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010001; // iC=  529 
vC = 14'b1111101100100000; // vC=-1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000000; // iC=  576 
vC = 14'b1111101100001111; // vC=-1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010010; // iC=  594 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000001; // iC=  641 
vC = 14'b1111101101000101; // vC=-1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011101; // iC=  733 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111010; // iC=  698 
vC = 14'b1111101011010001; // vC=-1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100010; // iC=  674 
vC = 14'b1111101100001010; // vC=-1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011010; // iC=  730 
vC = 14'b1111101011010001; // vC=-1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101110; // iC=  814 
vC = 14'b1111101100011011; // vC=-1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000111; // iC=  775 
vC = 14'b1111101011101110; // vC=-1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110000; // iC=  752 
vC = 14'b1111101011010010; // vC=-1326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001010; // iC=  842 
vC = 14'b1111101011111001; // vC=-1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010111; // iC=  791 
vC = 14'b1111101100110011; // vC=-1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000000; // iC=  896 
vC = 14'b1111101011101111; // vC=-1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011011; // iC=  923 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000100; // iC=  964 
vC = 14'b1111101101101110; // vC=-1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000000; // iC=  896 
vC = 14'b1111101101000110; // vC=-1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001010; // iC=  906 
vC = 14'b1111101100001110; // vC=-1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011001; // iC=  985 
vC = 14'b1111101100010110; // vC=-1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011011; // iC=  987 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010011; // iC=  915 
vC = 14'b1111101101000110; // vC=-1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100110; // iC= 1062 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011001; // iC= 1049 
vC = 14'b1111101101111010; // vC=-1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001011; // iC= 1099 
vC = 14'b1111101110001110; // vC=-1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111100; // iC= 1084 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010010; // iC= 1042 
vC = 14'b1111101100100111; // vC=-1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000000; // iC= 1088 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111011; // iC= 1147 
vC = 14'b1111101100001000; // vC=-1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001110; // iC= 1102 
vC = 14'b1111101100110011; // vC=-1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010010; // iC= 1170 
vC = 14'b1111101100111100; // vC=-1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101011; // iC= 1131 
vC = 14'b1111101100110001; // vC=-1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000111; // iC= 1223 
vC = 14'b1111101101100000; // vC=-1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010111; // iC= 1175 
vC = 14'b1111101110000110; // vC=-1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011011; // iC= 1307 
vC = 14'b1111101110010000; // vC=-1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110101; // iC= 1269 
vC = 14'b1111101110101111; // vC=-1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010011; // iC= 1299 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111111; // iC= 1215 
vC = 14'b1111101101011110; // vC=-1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000000; // iC= 1280 
vC = 14'b1111101100101110; // vC=-1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011110; // iC= 1246 
vC = 14'b1111101101001011; // vC=-1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111011; // iC= 1275 
vC = 14'b1111101111001011; // vC=-1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100110; // iC= 1318 
vC = 14'b1111101101001011; // vC=-1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011010; // iC= 1306 
vC = 14'b1111101111011100; // vC=-1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101000; // iC= 1320 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100100; // iC= 1380 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100001; // iC= 1441 
vC = 14'b1111101110001101; // vC=-1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111011; // iC= 1403 
vC = 14'b1111101110101000; // vC=-1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000010; // iC= 1410 
vC = 14'b1111101101111011; // vC=-1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101011; // iC= 1515 
vC = 14'b1111101111101101; // vC=-1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101110; // iC= 1518 
vC = 14'b1111101111100011; // vC=-1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010111; // iC= 1431 
vC = 14'b1111101110110111; // vC=-1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010100; // iC= 1428 
vC = 14'b1111101111101110; // vC=-1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000101; // iC= 1477 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100000; // iC= 1568 
vC = 14'b1111101111010010; // vC=-1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111011; // iC= 1595 
vC = 14'b1111101110001001; // vC=-1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010011; // iC= 1491 
vC = 14'b1111101110111010; // vC=-1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101110; // iC= 1518 
vC = 14'b1111110000010111; // vC=-1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110001; // iC= 1585 
vC = 14'b1111101111011010; // vC=-1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001001; // iC= 1609 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101111; // iC= 1583 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011001; // iC= 1625 
vC = 14'b1111110000011010; // vC= -998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100011; // iC= 1571 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110010; // iC= 1650 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111011; // iC= 1659 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b1111101111001110; // vC=-1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b1111110001011001; // vC= -935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010100; // iC= 1620 
vC = 14'b1111101111100110; // vC=-1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100010; // iC= 1762 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b1111110001010101; // vC= -939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b1111110001100100; // vC= -924 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110001; // iC= 1713 
vC = 14'b1111110010000010; // vC= -894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101000; // iC= 1640 
vC = 14'b1111110010001110; // vC= -882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000010; // iC= 1730 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111110001110101; // vC= -907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010101; // iC= 1685 
vC = 14'b1111110000110101; // vC= -971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111110000100011; // vC= -989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111100; // iC= 1788 
vC = 14'b1111110000110101; // vC= -971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001011; // iC= 1739 
vC = 14'b1111110010010110; // vC= -874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011100; // iC= 1820 
vC = 14'b1111110010101110; // vC= -850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110000; // iC= 1776 
vC = 14'b1111110011000110; // vC= -826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001101; // iC= 1869 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b1111110010011110; // vC= -866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101111; // iC= 1839 
vC = 14'b1111110001110010; // vC= -910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b1111110010100101; // vC= -859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b1111110011111101; // vC= -771 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b1111110010101000; // vC= -856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100100; // iC= 1764 
vC = 14'b1111110011010011; // vC= -813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b1111110100100000; // vC= -736 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000011; // iC= 1859 
vC = 14'b1111110010110011; // vC= -845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010000; // iC= 1808 
vC = 14'b1111110010110010; // vC= -846 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b1111110100101101; // vC= -723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b1111110011110010; // vC= -782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111110011111010; // vC= -774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111110100000111; // vC= -761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b1111110100110110; // vC= -714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000111; // iC= 1799 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010011; // iC= 1811 
vC = 14'b1111110100111010; // vC= -710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111110011111011; // vC= -773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b1111110100111100; // vC= -708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b1111110100111000; // vC= -712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111110101100001; // vC= -671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010001; // iC= 1873 
vC = 14'b1111110100010001; // vC= -751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b1111110100011110; // vC= -738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b1111110101101011; // vC= -661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b1111110101001010; // vC= -694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b1111110100111010; // vC= -710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110101; // iC= 1781 
vC = 14'b1111110111000010; // vC= -574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b1111110100110100; // vC= -716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b1111110101101000; // vC= -664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b1111110101010010; // vC= -686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b1111110101111100; // vC= -644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b1111110101101001; // vC= -663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b1111110111100101; // vC= -539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b1111110110001100; // vC= -628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001010; // iC= 1866 
vC = 14'b1111110111101000; // vC= -536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100011; // iC= 1827 
vC = 14'b1111110110110100; // vC= -588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111110110100010; // vC= -606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110110; // iC= 1846 
vC = 14'b1111110111110101; // vC= -523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101101; // iC= 1837 
vC = 14'b1111111000010011; // vC= -493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b1111110111000001; // vC= -575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001100; // iC= 1804 
vC = 14'b1111111000011101; // vC= -483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111001; // iC= 1785 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111110111111000; // vC= -520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b1111110111101111; // vC= -529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b1111111000110110; // vC= -458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b1111110111110110; // vC= -522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111110111111100; // vC= -516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b1111111000001101; // vC= -499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000100; // iC= 1860 
vC = 14'b1111110111010111; // vC= -553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b1111111000011100; // vC= -484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b1111110111100100; // vC= -540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111110111111000; // vC= -520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b1111111000111110; // vC= -450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111111000111111; // vC= -449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111111000001001; // vC= -503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111111001011011; // vC= -421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111111; // iC= 1791 
vC = 14'b1111111000001001; // vC= -503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111111000000111; // vC= -505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b1111111010001000; // vC= -376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b1111111001111001; // vC= -391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111111010110001; // vC= -335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b1111111000100101; // vC= -475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b1111111000101001; // vC= -471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b1111111001011111; // vC= -417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111111010110011; // vC= -333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b1111111011000111; // vC= -313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110110; // iC= 1846 
vC = 14'b1111111001011111; // vC= -417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111111001010001; // vC= -431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b1111111010000111; // vC= -377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110001; // iC= 1841 
vC = 14'b1111111011010111; // vC= -297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b1111111010011110; // vC= -354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b1111111010110010; // vC= -334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b1111111010110001; // vC= -335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b1111111011001010; // vC= -310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b1111111011111101; // vC= -259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111111100010101; // vC= -235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b1111111010111101; // vC= -323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111111011111001; // vC= -263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000010; // iC= 1858 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b1111111011111100; // vC= -260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110010; // iC= 1906 
vC = 14'b1111111100110010; // vC= -206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b1111111010110100; // vC= -332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101111; // iC= 1839 
vC = 14'b1111111100001000; // vC= -248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101111; // iC= 1839 
vC = 14'b1111111100110101; // vC= -203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111111100111111; // vC= -193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101110; // iC= 1838 
vC = 14'b1111111100101100; // vC= -212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011100; // iC= 1884 
vC = 14'b1111111100111100; // vC= -196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111100001001; // vC= -247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111111101011011; // vC= -165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b1111111011101011; // vC= -277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b1111111100110000; // vC= -208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b1111111100110111; // vC= -201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b1111111100111100; // vC= -196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b1111111110010000; // vC= -112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111111101101100; // vC= -148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101101; // iC= 1837 
vC = 14'b1111111100001101; // vC= -243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b1111111101101010; // vC= -150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111111110011011; // vC= -101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101010; // iC= 1898 
vC = 14'b1111111110010010; // vC= -110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001001; // iC= 1865 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111100111110; // vC= -194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111111111000000; // vC=  -64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110000; // iC= 1840 
vC = 14'b1111111111000111; // vC=  -57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011011; // iC= 1819 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101100; // iC= 1772 
vC = 14'b1111111110111110; // vC=  -66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010000; // iC= 1808 
vC = 14'b1111111111000001; // vC=  -63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111111110011100; // vC= -100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b1111111110000011; // vC= -125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b1111111101110010; // vC= -142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111111111111101; // vC=   -3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000000; // iC= 1792 
vC = 14'b1111111111001101; // vC=  -51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010011; // iC= 1811 
vC = 14'b1111111110100110; // vC=  -90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100110; // iC= 1830 
vC = 14'b0000000000010100; // vC=   20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111111110110100; // vC=  -76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000011; // iC= 1795 
vC = 14'b0000000000101010; // vC=   42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111100; // iC= 1788 
vC = 14'b1111111110101001; // vC=  -87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b1111111110111100; // vC=  -68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b0000000000011001; // vC=   25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111101; // iC= 1853 
vC = 14'b1111111110101101; // vC=  -83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b0000000000001000; // vC=    8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b0000000001010010; // vC=   82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b0000000001010010; // vC=   82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b0000000000110100; // vC=   52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110100; // iC= 1780 
vC = 14'b1111111111101000; // vC=  -24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b0000000000101001; // vC=   41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100110; // iC= 1830 
vC = 14'b0000000000010001; // vC=   17 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b1111111111101011; // vC=  -21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110110; // iC= 1846 
vC = 14'b0000000000110001; // vC=   49 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b0000000001110101; // vC=  117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b0000000000101000; // vC=   40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000111; // iC= 1799 
vC = 14'b1111111111111001; // vC=   -7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b0000000010011100; // vC=  156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000000000010110; // vC=   22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b0000000010110000; // vC=  176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b0000000000100001; // vC=   33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111001; // iC= 1849 
vC = 14'b0000000010101100; // vC=  172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b0000000001010101; // vC=   85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111100; // iC= 1724 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011011; // iC= 1755 
vC = 14'b0000000011100111; // vC=  231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110010; // iC= 1778 
vC = 14'b0000000011001100; // vC=  204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b0000000010101110; // vC=  174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001100; // iC= 1740 
vC = 14'b0000000010101010; // vC=  170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100011; // iC= 1763 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001001; // iC= 1865 
vC = 14'b0000000011111000; // vC=  248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b0000000100010000; // vC=  272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000000100011010; // vC=  282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000000010011011; // vC=  155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b0000000100100000; // vC=  288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b0000000010101010; // vC=  170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111101; // iC= 1789 
vC = 14'b0000000100101010; // vC=  298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111101; // iC= 1853 
vC = 14'b0000000011010100; // vC=  212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b0000000100010001; // vC=  273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011101; // iC= 1693 
vC = 14'b0000000011111001; // vC=  249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b0000000101001011; // vC=  331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b0000000011111101; // vC=  253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b0000000100101111; // vC=  303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001100; // iC= 1740 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b0000000011100111; // vC=  231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b0000000101110000; // vC=  368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b0000000101010111; // vC=  343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b0000000100100110; // vC=  294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b0000000101111001; // vC=  377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101011; // iC= 1707 
vC = 14'b0000000100010110; // vC=  278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b0000000101111111; // vC=  383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b0000000100000011; // vC=  259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100001; // iC= 1697 
vC = 14'b0000000100100001; // vC=  289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b0000000100011101; // vC=  285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b0000000100001110; // vC=  270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b0000000101011100; // vC=  348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000001; // iC= 1665 
vC = 14'b0000000101001110; // vC=  334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000000101010001; // vC=  337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101100; // iC= 1772 
vC = 14'b0000000110010000; // vC=  400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b0000000110011110; // vC=  414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b0000000100111001; // vC=  313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b0000000110100111; // vC=  423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000101; // iC= 1669 
vC = 14'b0000000101010100; // vC=  340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b0000000101101101; // vC=  365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010100; // iC= 1748 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100100; // iC= 1764 
vC = 14'b0000000111110010; // vC=  498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b0000000111010011; // vC=  467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011000; // iC= 1752 
vC = 14'b0000000110100010; // vC=  418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101111; // iC= 1711 
vC = 14'b0000000111010001; // vC=  465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000010; // iC= 1730 
vC = 14'b0000000111101010; // vC=  490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110111; // iC= 1655 
vC = 14'b0000000101111100; // vC=  380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101001; // iC= 1705 
vC = 14'b0000000111001001; // vC=  457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100011; // iC= 1763 
vC = 14'b0000000111000000; // vC=  448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101100; // iC= 1644 
vC = 14'b0000000110111111; // vC=  447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b0000000111110100; // vC=  500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001011; // iC= 1675 
vC = 14'b0000001000000110; // vC=  518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010011; // iC= 1747 
vC = 14'b0000000111101100; // vC=  492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b0000001000101010; // vC=  554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000000111111000; // vC=  504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b0000000110101000; // vC=  424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100110; // iC= 1638 
vC = 14'b0000001001000001; // vC=  577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b0000000111010010; // vC=  466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011100; // iC= 1628 
vC = 14'b0000001000110000; // vC=  560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b0000000111000100; // vC=  452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b0000001001101000; // vC=  616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100110; // iC= 1638 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001110; // iC= 1678 
vC = 14'b0000001000110111; // vC=  567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111111; // iC= 1599 
vC = 14'b0000001000000101; // vC=  517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010011; // iC= 1619 
vC = 14'b0000001000000010; // vC=  514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b0000000111101000; // vC=  488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001001; // iC= 1609 
vC = 14'b0000001001011111; // vC=  607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001110; // iC= 1678 
vC = 14'b0000001001001010; // vC=  586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011010; // iC= 1562 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b0000001001000011; // vC=  579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111000; // iC= 1592 
vC = 14'b0000001001110100; // vC=  628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100001; // iC= 1697 
vC = 14'b0000001000011110; // vC=  542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b0000001000110110; // vC=  566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010100; // iC= 1556 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101111; // iC= 1583 
vC = 14'b0000001010011010; // vC=  666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110100; // iC= 1652 
vC = 14'b0000001010110111; // vC=  695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010111; // iC= 1559 
vC = 14'b0000001001010111; // vC=  599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110111; // iC= 1527 
vC = 14'b0000001001101000; // vC=  616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110100; // iC= 1652 
vC = 14'b0000001010001100; // vC=  652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001100; // iC= 1612 
vC = 14'b0000001010010101; // vC=  661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b0000001001111000; // vC=  632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110101; // iC= 1589 
vC = 14'b0000001001011110; // vC=  606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111000; // iC= 1528 
vC = 14'b0000001010100111; // vC=  679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000000; // iC= 1600 
vC = 14'b0000001010111100; // vC=  700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111101; // iC= 1533 
vC = 14'b0000001010001000; // vC=  648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110111; // iC= 1655 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101101; // iC= 1645 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110110; // iC= 1654 
vC = 14'b0000001010001111; // vC=  655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101111; // iC= 1583 
vC = 14'b0000001011010010; // vC=  722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b0000001011101101; // vC=  749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101001; // iC= 1641 
vC = 14'b0000001010001100; // vC=  652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100101; // iC= 1509 
vC = 14'b0000001010000001; // vC=  641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100101; // iC= 1637 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000111; // iC= 1543 
vC = 14'b0000001010101100; // vC=  684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b0000001011110100; // vC=  756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110110; // iC= 1526 
vC = 14'b0000001100000110; // vC=  774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111001; // iC= 1593 
vC = 14'b0000001011111100; // vC=  764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100010; // iC= 1506 
vC = 14'b0000001011101100; // vC=  748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000110; // iC= 1606 
vC = 14'b0000001011101010; // vC=  746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011001; // iC= 1561 
vC = 14'b0000001010011100; // vC=  668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110001; // iC= 1585 
vC = 14'b0000001011011001; // vC=  729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010001; // iC= 1553 
vC = 14'b0000001010111101; // vC=  701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001010; // iC= 1546 
vC = 14'b0000001100100010; // vC=  802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010011; // iC= 1555 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101011; // iC= 1515 
vC = 14'b0000001100011011; // vC=  795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011101; // iC= 1437 
vC = 14'b0000001100011110; // vC=  798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000100; // iC= 1476 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110100; // iC= 1524 
vC = 14'b0000001011010001; // vC=  721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110010; // iC= 1522 
vC = 14'b0000001101010101; // vC=  853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001111; // iC= 1551 
vC = 14'b0000001101100000; // vC=  864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111110; // iC= 1534 
vC = 14'b0000001100110101; // vC=  821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001101; // iC= 1421 
vC = 14'b0000001100010110; // vC=  790 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011100; // iC= 1500 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000101; // iC= 1413 
vC = 14'b0000001101000110; // vC=  838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111000; // iC= 1528 
vC = 14'b0000001101100011; // vC=  867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001101; // iC= 1485 
vC = 14'b0000001100010111; // vC=  791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011100; // iC= 1436 
vC = 14'b0000001110001011; // vC=  907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001010; // iC= 1546 
vC = 14'b0000001100000101; // vC=  773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111111; // iC= 1535 
vC = 14'b0000001110001001; // vC=  905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111110; // iC= 1406 
vC = 14'b0000001101101011; // vC=  875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011110; // iC= 1502 
vC = 14'b0000001101110101; // vC=  885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000111; // iC= 1479 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110010; // iC= 1458 
vC = 14'b0000001101000000; // vC=  832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001111; // iC= 1487 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001100; // iC= 1484 
vC = 14'b0000001110001110; // vC=  910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101111; // iC= 1391 
vC = 14'b0000001101110101; // vC=  885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111001; // iC= 1465 
vC = 14'b0000001101100000; // vC=  864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101100; // iC= 1452 
vC = 14'b0000001101110001; // vC=  881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000110; // iC= 1350 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011000; // iC= 1368 
vC = 14'b0000001101101010; // vC=  874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001110; // iC= 1422 
vC = 14'b0000001110001100; // vC=  908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001110; // iC= 1422 
vC = 14'b0000001101010000; // vC=  848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000000; // iC= 1408 
vC = 14'b0000001110100011; // vC=  931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101000; // iC= 1448 
vC = 14'b0000001111011100; // vC=  988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011001; // iC= 1369 
vC = 14'b0000001110110110; // vC=  950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111101; // iC= 1405 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011110; // iC= 1374 
vC = 14'b0000001111100001; // vC=  993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010101; // iC= 1429 
vC = 14'b0000001111010010; // vC=  978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b0000001111000100; // vC=  964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010111; // iC= 1303 
vC = 14'b0000001110011111; // vC=  927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110101; // iC= 1333 
vC = 14'b0000001111101101; // vC= 1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000010; // iC= 1346 
vC = 14'b0000001111100110; // vC=  998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101011; // iC= 1451 
vC = 14'b0000001110101010; // vC=  938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000100; // iC= 1348 
vC = 14'b0000001110100100; // vC=  932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010101; // iC= 1301 
vC = 14'b0000001111101110; // vC= 1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100101; // iC= 1317 
vC = 14'b0000001110000010; // vC=  898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111001; // iC= 1337 
vC = 14'b0000001110010001; // vC=  913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111010; // iC= 1402 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101011; // iC= 1387 
vC = 14'b0000001111100101; // vC=  997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010010; // iC= 1298 
vC = 14'b0000001111000101; // vC=  965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010001; // iC= 1361 
vC = 14'b0000001110101110; // vC=  942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100000; // iC= 1376 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111010; // iC= 1338 
vC = 14'b0000010000001101; // vC= 1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011111; // iC= 1247 
vC = 14'b0000001111110011; // vC= 1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010100; // iC= 1300 
vC = 14'b0000010000000101; // vC= 1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111111; // iC= 1343 
vC = 14'b0000001111001110; // vC=  974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101010; // iC= 1386 
vC = 14'b0000001110110100; // vC=  948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001111; // iC= 1295 
vC = 14'b0000001111111010; // vC= 1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000000; // iC= 1344 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100101; // iC= 1253 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000001; // iC= 1217 
vC = 14'b0000010000011010; // vC= 1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101101; // iC= 1261 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100100; // iC= 1316 
vC = 14'b0000010000000111; // vC= 1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110111; // iC= 1271 
vC = 14'b0000001111000110; // vC=  966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001110; // iC= 1294 
vC = 14'b0000010000001001; // vC= 1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001000; // iC= 1352 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011011; // iC= 1307 
vC = 14'b0000001111110011; // vC= 1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b0000010000111111; // vC= 1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010101; // iC= 1237 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110111; // iC= 1271 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110000; // iC= 1264 
vC = 14'b0000010000111001; // vC= 1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110010; // iC= 1266 
vC = 14'b0000010001110110; // vC= 1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110110; // iC= 1270 
vC = 14'b0000010000100001; // vC= 1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000100; // iC= 1220 
vC = 14'b0000010000000100; // vC= 1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000010; // iC= 1218 
vC = 14'b0000010000100001; // vC= 1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110101; // iC= 1205 
vC = 14'b0000010000100101; // vC= 1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000111; // iC= 1287 
vC = 14'b0000010001110000; // vC= 1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001111; // iC= 1167 
vC = 14'b0000001111110111; // vC= 1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011000; // iC= 1240 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110110; // iC= 1206 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001001; // iC= 1289 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111010; // iC= 1146 
vC = 14'b0000010010000000; // vC= 1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111110; // iC= 1278 
vC = 14'b0000010010000000; // vC= 1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111001; // iC= 1209 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010101; // iC= 1237 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100000; // iC= 1120 
vC = 14'b0000010010000101; // vC= 1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000010010110101; // vC= 1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001001; // iC= 1097 
vC = 14'b0000010010000000; // vC= 1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111110; // iC= 1150 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101010; // iC= 1194 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011010; // iC= 1114 
vC = 14'b0000010001101110; // vC= 1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011101; // iC= 1117 
vC = 14'b0000010010001111; // vC= 1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111011; // iC= 1211 
vC = 14'b0000010010101001; // vC= 1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001100; // iC= 1100 
vC = 14'b0000010010101011; // vC= 1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101110; // iC= 1070 
vC = 14'b0000010011010001; // vC= 1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011100; // iC= 1116 
vC = 14'b0000010010101101; // vC= 1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100110; // iC= 1062 
vC = 14'b0000010010101110; // vC= 1198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111100; // iC= 1212 
vC = 14'b0000010011000011; // vC= 1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010111; // iC= 1111 
vC = 14'b0000010011011010; // vC= 1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001101; // iC= 1101 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010100; // iC= 1044 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000110; // iC= 1094 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100000; // iC= 1120 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010101; // iC= 1173 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000110; // iC= 1094 
vC = 14'b0000010001111101; // vC= 1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100101; // iC= 1061 
vC = 14'b0000010011111001; // vC= 1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010100; // iC= 1108 
vC = 14'b0000010010110001; // vC= 1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100001; // iC= 1057 
vC = 14'b0000010001101110; // vC= 1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000011; // iC= 1091 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000000; // iC= 1088 
vC = 14'b0000010010101101; // vC= 1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000100; // iC= 1092 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101001; // iC= 1065 
vC = 14'b0000010010001001; // vC= 1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110010; // iC= 1138 
vC = 14'b0000010010101101; // vC= 1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000000; // iC= 1024 
vC = 14'b0000010010100011; // vC= 1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101101; // iC= 1005 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101101; // iC= 1069 
vC = 14'b0000010011110101; // vC= 1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100110; // iC= 1062 
vC = 14'b0000010010000000; // vC= 1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010000; // iC= 1040 
vC = 14'b0000010100011000; // vC= 1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110110; // iC= 1014 
vC = 14'b0000010100010000; // vC= 1296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010011; // iC= 1043 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010000; // iC= 1104 
vC = 14'b0000010100100000; // vC= 1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110100; // iC=  948 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111010; // iC=  954 
vC = 14'b0000010010011110; // vC= 1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000011; // iC= 1027 
vC = 14'b0000010011100000; // vC= 1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010101; // iC= 1045 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011000; // iC= 1048 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101100; // iC=  940 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000100; // iC= 1028 
vC = 14'b0000010011110011; // vC= 1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010111; // iC=  919 
vC = 14'b0000010010100100; // vC= 1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000111; // iC=  967 
vC = 14'b0000010010101111; // vC= 1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010000; // iC=  912 
vC = 14'b0000010100111011; // vC= 1339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010011; // iC=  915 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010001; // iC=  913 
vC = 14'b0000010100010011; // vC= 1299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111010; // iC= 1018 
vC = 14'b0000010100110100; // vC= 1332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110101; // iC=  885 
vC = 14'b0000010010110011; // vC= 1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000001; // iC=  897 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101000; // iC= 1000 
vC = 14'b0000010100010110; // vC= 1302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101011; // iC= 1003 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000111; // iC=  967 
vC = 14'b0000010101011100; // vC= 1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100011; // iC=  995 
vC = 14'b0000010011100011; // vC= 1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100111; // iC=  999 
vC = 14'b0000010100100001; // vC= 1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011011; // iC=  987 
vC = 14'b0000010101010001; // vC= 1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010100; // iC=  852 
vC = 14'b0000010011100000; // vC= 1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110001; // iC=  881 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110011; // iC=  883 
vC = 14'b0000010011001110; // vC= 1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110010; // iC=  818 
vC = 14'b0000010011101100; // vC= 1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001010; // iC=  906 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011001; // iC=  921 
vC = 14'b0000010100110000; // vC= 1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101101; // iC=  877 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101101; // iC=  941 
vC = 14'b0000010100011100; // vC= 1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010011; // iC=  915 
vC = 14'b0000010100100100; // vC= 1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101011; // iC=  875 
vC = 14'b0000010011100001; // vC= 1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110111; // iC=  823 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110111; // iC=  887 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010110; // iC=  854 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000110; // iC=  902 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011101; // iC=  861 
vC = 14'b0000010101000011; // vC= 1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011011; // iC=  795 
vC = 14'b0000010011111010; // vC= 1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111110; // iC=  830 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001000; // iC=  904 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110110; // iC=  758 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011111; // iC=  735 
vC = 14'b0000010101100100; // vC= 1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001010; // iC=  778 
vC = 14'b0000010100011000; // vC= 1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110001; // iC=  817 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100011; // iC=  739 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101001; // iC=  809 
vC = 14'b0000010100010110; // vC= 1302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010111; // iC=  791 
vC = 14'b0000010100001000; // vC= 1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110000; // iC=  816 
vC = 14'b0000010101110111; // vC= 1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110111; // iC=  759 
vC = 14'b0000010101001101; // vC= 1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000110; // iC=  838 
vC = 14'b0000010110000010; // vC= 1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011001; // iC=  729 
vC = 14'b0000010100111000; // vC= 1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100101; // iC=  805 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000011; // iC=  771 
vC = 14'b0000010101111000; // vC= 1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101010; // iC=  746 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101010; // iC=  746 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010001; // iC=  785 
vC = 14'b0000010101011010; // vC= 1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111001; // iC=  697 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100100; // iC=  676 
vC = 14'b0000010101100111; // vC= 1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100111; // iC=  679 
vC = 14'b0000010101100010; // vC= 1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010001; // iC=  785 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110110; // iC=  694 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000110; // iC=  710 
vC = 14'b0000010101111100; // vC= 1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111000; // iC=  696 
vC = 14'b0000010110010111; // vC= 1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111011; // iC=  635 
vC = 14'b0000010110010110; // vC= 1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010100; // iC=  724 
vC = 14'b0000010110111010; // vC= 1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101011; // iC=  619 
vC = 14'b0000010110101001; // vC= 1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011001; // iC=  665 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100010; // iC=  674 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101110; // iC=  750 
vC = 14'b0000010100111000; // vC= 1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000011; // iC=  707 
vC = 14'b0000010101010001; // vC= 1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010000; // iC=  592 
vC = 14'b0000010110111101; // vC= 1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100101; // iC=  741 
vC = 14'b0000010110101000; // vC= 1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000110; // iC=  582 
vC = 14'b0000010101000110; // vC= 1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100001; // iC=  609 
vC = 14'b0000010101101101; // vC= 1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000001; // iC=  641 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101010; // iC=  618 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000010; // iC=  642 
vC = 14'b0000010110110011; // vC= 1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101110; // iC=  622 
vC = 14'b0000010110010100; // vC= 1428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101101; // iC=  557 
vC = 14'b0000010101010111; // vC= 1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100101; // iC=  677 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001110; // iC=  654 
vC = 14'b0000010110110010; // vC= 1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111101; // iC=  573 
vC = 14'b0000010111100111; // vC= 1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110110; // iC=  566 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011100; // iC=  540 
vC = 14'b0000010101011110; // vC= 1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011011; // iC=  603 
vC = 14'b0000010111010011; // vC= 1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110010; // iC=  562 
vC = 14'b0000010110000100; // vC= 1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111001; // iC=  569 
vC = 14'b0000010110111111; // vC= 1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110011; // iC=  563 
vC = 14'b0000010111010010; // vC= 1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011101; // iC=  605 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000111; // iC=  519 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110011; // iC=  563 
vC = 14'b0000010110001000; // vC= 1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001100; // iC=  588 
vC = 14'b0000010111001111; // vC= 1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100110; // iC=  614 
vC = 14'b0000010110100001; // vC= 1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010110; // iC=  534 
vC = 14'b0000010111001111; // vC= 1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010110; // iC=  598 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010100; // iC=  468 
vC = 14'b0000010110011100; // vC= 1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100000; // iC=  544 
vC = 14'b0000010111011000; // vC= 1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011011; // iC=  475 
vC = 14'b0000010110111110; // vC= 1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111000; // iC=  504 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101000; // iC=  552 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111000; // iC=  440 
vC = 14'b0000010110000010; // vC= 1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110000; // iC=  560 
vC = 14'b0000010111101100; // vC= 1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100100; // iC=  420 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101111; // iC=  559 
vC = 14'b0000010111010000; // vC= 1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000000; // iC=  448 
vC = 14'b0000010110011111; // vC= 1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101100; // iC=  428 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100000; // iC=  480 
vC = 14'b0000010111001000; // vC= 1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000110; // iC=  390 
vC = 14'b0000010111011001; // vC= 1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000010; // iC=  514 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011100; // iC=  476 
vC = 14'b0000010101101010; // vC= 1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000111; // iC=  455 
vC = 14'b0000010110101000; // vC= 1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101100; // iC=  492 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101100; // iC=  364 
vC = 14'b0000010110101000; // vC= 1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001110; // iC=  398 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101010; // iC=  490 
vC = 14'b0000010101110111; // vC= 1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010100; // iC=  340 
vC = 14'b0000010101110010; // vC= 1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011110; // iC=  414 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010000; // iC=  336 
vC = 14'b0000010111110100; // vC= 1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001011; // iC=  395 
vC = 14'b0000010111110100; // vC= 1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000110; // iC=  390 
vC = 14'b0000010110010110; // vC= 1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111100; // iC=  380 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100010; // iC=  290 
vC = 14'b0000010111010010; // vC= 1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011000; // iC=  280 
vC = 14'b0000011000010010; // vC= 1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111011; // iC=  379 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000100; // iC=  260 
vC = 14'b0000010110110111; // vC= 1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010111; // iC=  343 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100011; // iC=  227 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001111; // iC=  207 
vC = 14'b0000010111011101; // vC= 1501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100101; // iC=  229 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010101; // iC=  213 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111100; // iC=  188 
vC = 14'b0000010111011100; // vC= 1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010110; // iC=  150 
vC = 14'b0000010111111011; // vC= 1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011110; // iC=  222 
vC = 14'b0000010111001110; // vC= 1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000101; // iC=  133 
vC = 14'b0000010110001010; // vC= 1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001000; // iC=  136 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110101; // iC=  117 
vC = 14'b0000010110110100; // vC= 1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001010; // iC=   74 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110011; // iC=  115 
vC = 14'b0000010110111010; // vC= 1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101111; // iC=   47 
vC = 14'b0000010110001110; // vC= 1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010100; // iC=   84 
vC = 14'b0000010110001110; // vC= 1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110100; // iC=  116 
vC = 14'b0000010110001100; // vC= 1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100001; // iC=   33 
vC = 14'b0000010111110010; // vC= 1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011001; // iC=   25 
vC = 14'b0000011000010011; // vC= 1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110101; // iC=  -11 
vC = 14'b0000010111110001; // vC= 1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110001; // iC=  -15 
vC = 14'b0000010111011011; // vC= 1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110011; // iC=   51 
vC = 14'b0000010111110100; // vC= 1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110010; // iC=  -14 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010110; // iC= -106 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001110; // iC=  -50 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110100; // iC=  -12 
vC = 14'b0000010111110001; // vC= 1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111110; // iC= -130 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010110; // iC= -106 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011100; // iC= -100 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111100; // iC=  -68 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010110; // iC= -106 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100011; // iC= -221 
vC = 14'b0000010110101101; // vC= 1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110010; // iC= -270 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011110; // iC= -290 
vC = 14'b0000010110111010; // vC= 1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011101; // iC= -291 
vC = 14'b0000010111100100; // vC= 1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000110; // iC= -314 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111111; // iC= -257 
vC = 14'b0000010111001001; // vC= 1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110001; // iC= -271 
vC = 14'b0000010101101111; // vC= 1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000100; // iC= -380 
vC = 14'b0000010110010001; // vC= 1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100000; // iC= -288 
vC = 14'b0000010101100101; // vC= 1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001101; // iC= -371 
vC = 14'b0000010110010111; // vC= 1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111001; // iC= -455 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000101; // iC= -443 
vC = 14'b0000010110011110; // vC= 1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101101; // iC= -403 
vC = 14'b0000010111010010; // vC= 1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100001; // iC= -479 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001110; // iC= -562 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001111; // iC= -561 
vC = 14'b0000010110101001; // vC= 1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110000; // iC= -592 
vC = 14'b0000010110111010; // vC= 1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000011; // iC= -573 
vC = 14'b0000010101010100; // vC= 1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010110; // iC= -554 
vC = 14'b0000010101111011; // vC= 1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110011; // iC= -589 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b0000010110000100; // vC= 1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111101; // iC= -579 
vC = 14'b0000010110001110; // vC= 1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011011; // iC= -613 
vC = 14'b0000010101111000; // vC= 1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101011; // iC= -725 
vC = 14'b0000010101011111; // vC= 1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000101; // iC= -635 
vC = 14'b0000010101001111; // vC= 1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100101; // iC= -667 
vC = 14'b0000010101010111; // vC= 1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010000; // iC= -688 
vC = 14'b0000010111000101; // vC= 1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001100; // iC= -820 
vC = 14'b0000010101010101; // vC= 1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010110; // iC= -810 
vC = 14'b0000010101100011; // vC= 1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111011; // iC= -837 
vC = 14'b0000010110000100; // vC= 1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010101; // iC= -811 
vC = 14'b0000010101110111; // vC= 1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111011; // iC= -773 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111111; // iC= -833 
vC = 14'b0000010101111100; // vC= 1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101100; // iC= -852 
vC = 14'b0000010100110100; // vC= 1332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111011; // iC= -901 
vC = 14'b0000010101111110; // vC= 1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001101; // iC= -883 
vC = 14'b0000010100011001; // vC= 1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010011; // iC= -941 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111000; // iC= -904 
vC = 14'b0000010101000100; // vC= 1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011101; // iC= -931 
vC = 14'b0000010100011101; // vC= 1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001011; // iC= -949 
vC = 14'b0000010101001100; // vC= 1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111111; // iC=-1025 
vC = 14'b0000010100101011; // vC= 1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000111; // iC= -953 
vC = 14'b0000010101110010; // vC= 1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011110; // iC=-1058 
vC = 14'b0000010011111011; // vC= 1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101011; // iC=-1109 
vC = 14'b0000010101100011; // vC= 1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010101; // iC=-1003 
vC = 14'b0000010100110011; // vC= 1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011000; // iC=-1064 
vC = 14'b0000010100111000; // vC= 1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101101; // iC=-1107 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101000; // iC=-1176 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110101; // iC=-1163 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111000; // iC=-1160 
vC = 14'b0000010100111111; // vC= 1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111000; // iC=-1096 
vC = 14'b0000010100000011; // vC= 1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001110; // iC=-1138 
vC = 14'b0000010101101101; // vC= 1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110100; // iC=-1228 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111111; // iC=-1153 
vC = 14'b0000010100100010; // vC= 1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111100; // iC=-1156 
vC = 14'b0000010100111110; // vC= 1342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000111; // iC=-1209 
vC = 14'b0000010100011100; // vC= 1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000111; // iC=-1209 
vC = 14'b0000010100100111; // vC= 1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000100; // iC=-1340 
vC = 14'b0000010101001100; // vC= 1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100101; // iC=-1307 
vC = 14'b0000010011000011; // vC= 1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101011; // iC=-1237 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100110; // iC=-1306 
vC = 14'b0000010100010100; // vC= 1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100010; // iC=-1246 
vC = 14'b0000010011101010; // vC= 1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000000; // iC=-1344 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110010; // iC=-1294 
vC = 14'b0000010100100001; // vC= 1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110110; // iC=-1354 
vC = 14'b0000010100011000; // vC= 1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001110; // iC=-1330 
vC = 14'b0000010011110011; // vC= 1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101000; // iC=-1304 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101100; // iC=-1428 
vC = 14'b0000010100001010; // vC= 1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110110; // iC=-1418 
vC = 14'b0000010010011010; // vC= 1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011111; // iC=-1377 
vC = 14'b0000010011110110; // vC= 1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101011; // iC=-1429 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b0000010011100101; // vC= 1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000011; // iC=-1469 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b0000010011010001; // vC= 1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110010; // iC=-1422 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011101; // iC=-1507 
vC = 14'b0000010010010110; // vC= 1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b0000010001010100; // vC= 1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b0000010010110101; // vC= 1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000010010110110; // vC= 1206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b0000010000111011; // vC= 1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101011; // iC=-1493 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001010; // iC=-1526 
vC = 14'b0000010010001111; // vC= 1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b0000010001011110; // vC= 1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b0000010000101100; // vC= 1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b0000010000100000; // vC= 1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011101; // iC=-1507 
vC = 14'b0000010000110001; // vC= 1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000001; // iC=-1599 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110001; // iC=-1615 
vC = 14'b0000010000000111; // vC= 1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b0000001111011101; // vC=  989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110101; // iC=-1611 
vC = 14'b0000010000000111; // vC= 1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110110; // iC=-1610 
vC = 14'b0000010000001100; // vC= 1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110111; // iC=-1545 
vC = 14'b0000001110011011; // vC=  923 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b0000001111100001; // vC=  993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b0000001111000100; // vC=  964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101100; // iC=-1556 
vC = 14'b0000001111000010; // vC=  962 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001010; // iC=-1654 
vC = 14'b0000001110010111; // vC=  919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b0000001110011101; // vC=  925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b0000001110111001; // vC=  953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b0000010000001100; // vC= 1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b0000001110101010; // vC=  938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100000; // iC=-1632 
vC = 14'b0000001110100000; // vC=  928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001000; // iC=-1656 
vC = 14'b0000001110001111; // vC=  911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b0000001111011101; // vC=  989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b0000001110010000; // vC=  912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b0000001110101000; // vC=  936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b0000001110101110; // vC=  942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b0000001110000011; // vC=  899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b0000001101011011; // vC=  859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b0000001110110000; // vC=  944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b0000001110000110; // vC=  902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110101; // iC=-1611 
vC = 14'b0000001110100100; // vC=  932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b0000001101111101; // vC=  893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b0000001100001000; // vC=  776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b0000001100111011; // vC=  827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000001100001001; // vC=  777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000001100101001; // vC=  809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b0000001100100011; // vC=  803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b0000001110000101; // vC=  901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000001011100000; // vC=  736 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b0000001101010010; // vC=  850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000001011010110; // vC=  726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011111; // iC=-1633 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b0000001011011100; // vC=  732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000001011110010; // vC=  754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b0000001011011010; // vC=  730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b0000001101000001; // vC=  833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000001011101100; // vC=  748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b0000001011000110; // vC=  710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000001010011010; // vC=  666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b0000001010011110; // vC=  670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000001010101100; // vC=  684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b0000001011101001; // vC=  745 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100011; // iC=-1693 
vC = 14'b0000001100010101; // vC=  789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101111; // iC=-1617 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b0000001010001001; // vC=  649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b0000001011011111; // vC=  735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b0000001011111011; // vC=  763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000001011011100; // vC=  732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000001010100111; // vC=  679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101101; // iC=-1683 
vC = 14'b0000001001110000; // vC=  624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b0000001010011001; // vC=  665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b0000001001101110; // vC=  622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000100; // iC=-1724 
vC = 14'b0000001001100010; // vC=  610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000001010010001; // vC=  657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b0000001010000101; // vC=  645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b0000001010100011; // vC=  675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b0000001000010010; // vC=  530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101010; // iC=-1686 
vC = 14'b0000001000011111; // vC=  543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000001000000001; // vC=  513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b0000001001110000; // vC=  624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b0000001000110100; // vC=  564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000001000001110; // vC=  526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b0000001000101101; // vC=  557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000001000110110; // vC=  566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b0000000111111001; // vC=  505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000001000111110; // vC=  574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000001001001001; // vC=  585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b0000001001010111; // vC=  599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000000110111111; // vC=  447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b0000001000110111; // vC=  567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001000; // iC=-1656 
vC = 14'b0000001000110100; // vC=  564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000000110101111; // vC=  431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100100; // iC=-1692 
vC = 14'b0000000111101010; // vC=  490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b0000000110011010; // vC=  410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b0000000111111100; // vC=  508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100101; // iC=-1627 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000000111001011; // vC=  459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b0000000111010110; // vC=  470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000001; // iC=-1663 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b0000000110000001; // vC=  385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000010; // iC=-1662 
vC = 14'b0000000110001111; // vC=  399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000000110010000; // vC=  400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b0000000111001000; // vC=  456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100000; // iC=-1632 
vC = 14'b0000000101010111; // vC=  343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b0000000110011110; // vC=  414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b0000000101011001; // vC=  345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b0000000110101111; // vC=  431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b0000000101101011; // vC=  363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000000110011100; // vC=  412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000000110000001; // vC=  385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b0000000101001110; // vC=  334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001010; // iC=-1654 
vC = 14'b0000000110100010; // vC=  418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000000110001000; // vC=  392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000000101111010; // vC=  378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b0000000100010111; // vC=  279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000000100010000; // vC=  272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b0000000100100010; // vC=  290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b0000000011100111; // vC=  231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b0000000011110011; // vC=  243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000000100001101; // vC=  269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b0000000101010011; // vC=  339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000000101100111; // vC=  359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b0000000101001100; // vC=  332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000000101010110; // vC=  342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b0000000011101000; // vC=  232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000000011000010; // vC=  194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000010; // iC=-1662 
vC = 14'b0000000100100111; // vC=  295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b0000000100101110; // vC=  302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110110; // iC=-1674 
vC = 14'b0000000011110111; // vC=  247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110000; // iC=-1680 
vC = 14'b0000000011100000; // vC=  224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000000011001000; // vC=  200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110100; // iC=-1612 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110000; // iC=-1680 
vC = 14'b0000000011100101; // vC=  229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000000010100111; // vC=  167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110110; // iC=-1610 
vC = 14'b0000000011101101; // vC=  237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b0000000010000011; // vC=  131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000000010110101; // vC=  181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b0000000011110000; // vC=  240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b0000000001011011; // vC=   91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000000001100000; // vC=   96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b0000000001000101; // vC=   69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100100; // iC=-1692 
vC = 14'b0000000010010011; // vC=  147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110101; // iC=-1611 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b0000000001011011; // vC=   91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011010; // iC=-1702 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b0000000000010110; // vC=   22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000000000001101; // vC=   13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010100; // iC=-1644 
vC = 14'b0000000001010011; // vC=   83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010100; // iC=-1644 
vC = 14'b0000000001011111; // vC=   95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b0000000010000011; // vC=  131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b0000000000000010; // vC=    2 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000000000100011; // vC=   35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000000000111101; // vC=   61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100101; // iC=-1627 
vC = 14'b1111111111011001; // vC=  -39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b1111111111001100; // vC=  -52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110111; // iC=-1673 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000000000100001; // vC=   33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100100; // iC=-1628 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110101; // iC=-1611 
vC = 14'b1111111111011101; // vC=  -35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010010; // iC=-1582 
vC = 14'b1111111111111111; // vC=   -1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b1111111111010000; // vC=  -48 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b0000000000000011; // vC=    3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b1111111111011000; // vC=  -40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b0000000000001011; // vC=   11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001000; // iC=-1656 
vC = 14'b1111111110101001; // vC=  -87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b1111111110100010; // vC=  -94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011101; // iC=-1699 
vC = 14'b1111111111000111; // vC=  -57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b0000000000001010; // vC=   10 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b1111111111110010; // vC=  -14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b1111111111110001; // vC=  -15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000111; // iC=-1657 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101001; // iC=-1623 
vC = 14'b1111111101010001; // vC= -175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100101; // iC=-1691 
vC = 14'b1111111111011000; // vC=  -40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b1111111101010001; // vC= -175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b1111111111000100; // vC=  -60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b1111111110001110; // vC= -114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b1111111110100000; // vC=  -96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100000; // iC=-1632 
vC = 14'b1111111100111010; // vC= -198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b1111111100111110; // vC= -194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101101; // iC=-1683 
vC = 14'b1111111110001000; // vC= -120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b1111111110100111; // vC=  -89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101011; // iC=-1557 
vC = 14'b1111111100111100; // vC= -196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110110; // iC=-1610 
vC = 14'b1111111101111100; // vC= -132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b1111111100110110; // vC= -202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b1111111101101011; // vC= -149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b1111111101111011; // vC= -133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b1111111110010011; // vC= -109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b1111111100001001; // vC= -247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b1111111100010100; // vC= -236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b1111111101001000; // vC= -184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b1111111101001011; // vC= -181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b1111111011101000; // vC= -280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b1111111101000110; // vC= -186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b1111111011010011; // vC= -301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111011; // iC=-1541 
vC = 14'b1111111100100000; // vC= -224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b1111111011110011; // vC= -269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b1111111100010010; // vC= -238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100011; // iC=-1565 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b1111111100111101; // vC= -195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001100; // iC=-1588 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b1111111011111100; // vC= -260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000111; // iC=-1529 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b1111111010100100; // vC= -348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b1111111100000101; // vC= -251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b1111111100001111; // vC= -241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b1111111010001001; // vC= -375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b1111111011001101; // vC= -307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010011; // iC=-1517 
vC = 14'b1111111011100110; // vC= -282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b1111111011010001; // vC= -303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000011; // iC=-1533 
vC = 14'b1111111011110001; // vC= -271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b1111111010001011; // vC= -373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111110; // iC=-1538 
vC = 14'b1111111001101001; // vC= -407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b1111111010010111; // vC= -361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110010; // iC=-1486 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b1111111011001111; // vC= -305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101001; // iC=-1623 
vC = 14'b1111111010111011; // vC= -325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100100; // iC=-1628 
vC = 14'b1111111001011111; // vC= -417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b1111111001111100; // vC= -388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b1111111011000001; // vC= -319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b1111111001101100; // vC= -404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110001; // iC=-1551 
vC = 14'b1111111010100011; // vC= -349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001010; // iC=-1462 
vC = 14'b1111111000101010; // vC= -470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110001; // iC=-1487 
vC = 14'b1111111001001011; // vC= -437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b1111111001111101; // vC= -387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b1111111000100011; // vC= -477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b1111111010100101; // vC= -347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001000; // iC=-1464 
vC = 14'b1111111000101010; // vC= -470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b1111111001010111; // vC= -425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b1111111000001100; // vC= -500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b1111111000111111; // vC= -449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110001; // iC=-1487 
vC = 14'b1111110111101110; // vC= -530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b1111111010000011; // vC= -381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100100; // iC=-1500 
vC = 14'b1111111010000100; // vC= -380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001011; // iC=-1461 
vC = 14'b1111111001010110; // vC= -426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b1111111001011111; // vC= -417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110010; // iC=-1422 
vC = 14'b1111111000111111; // vC= -449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011101; // iC=-1507 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b1111111001010010; // vC= -430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b1111110111011010; // vC= -550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b1111111001010110; // vC= -426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b1111110110111010; // vC= -582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b1111111001010000; // vC= -432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111111; // iC=-1537 
vC = 14'b1111110111101101; // vC= -531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b1111111000010010; // vC= -494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b1111110110111011; // vC= -581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b1111110110100001; // vC= -607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011011; // iC=-1381 
vC = 14'b1111110110111111; // vC= -577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b1111110110010111; // vC= -617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b1111110111100000; // vC= -544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110100; // iC=-1420 
vC = 14'b1111110110011000; // vC= -616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011001; // iC=-1383 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011011; // iC=-1381 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101011; // iC=-1493 
vC = 14'b1111110111000000; // vC= -576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110101; // iC=-1355 
vC = 14'b1111110111011000; // vC= -552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010111; // iC=-1385 
vC = 14'b1111110111111010; // vC= -518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010110; // iC=-1386 
vC = 14'b1111110110010110; // vC= -618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111111; // iC=-1473 
vC = 14'b1111110111110101; // vC= -523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b1111110111011000; // vC= -552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b1111110111000111; // vC= -569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b1111110110000000; // vC= -640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000111; // iC=-1337 
vC = 14'b1111110110000000; // vC= -640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110110; // iC=-1418 
vC = 14'b1111110110101101; // vC= -595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b1111110110101011; // vC= -597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101010; // iC=-1430 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010101; // iC=-1387 
vC = 14'b1111110110100000; // vC= -608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001110; // iC=-1330 
vC = 14'b1111110110100010; // vC= -606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111100; // iC=-1412 
vC = 14'b1111110110111000; // vC= -584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b1111110101100101; // vC= -667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100000; // iC=-1312 
vC = 14'b1111110101000000; // vC= -704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111001; // iC=-1351 
vC = 14'b1111110101100011; // vC= -669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010011; // iC=-1325 
vC = 14'b1111110110011110; // vC= -610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111010; // iC=-1414 
vC = 14'b1111110100101000; // vC= -728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001100; // iC=-1396 
vC = 14'b1111110110011010; // vC= -614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110100; // iC=-1420 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b1111110110001011; // vC= -629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110010; // iC=-1422 
vC = 14'b1111110011111000; // vC= -776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111111; // iC=-1281 
vC = 14'b1111110101110001; // vC= -655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100011; // iC=-1309 
vC = 14'b1111110011110111; // vC= -777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001101; // iC=-1395 
vC = 14'b1111110100011100; // vC= -740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b1111110100000101; // vC= -763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b1111110101110110; // vC= -650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100000; // iC=-1376 
vC = 14'b1111110011101011; // vC= -789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001010; // iC=-1398 
vC = 14'b1111110100101011; // vC= -725 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101000; // iC=-1304 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000100; // iC=-1404 
vC = 14'b1111110011010011; // vC= -813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001111; // iC=-1329 
vC = 14'b1111110100111110; // vC= -706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010001; // iC=-1327 
vC = 14'b1111110101001011; // vC= -693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001010; // iC=-1270 
vC = 14'b1111110100011000; // vC= -744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100011; // iC=-1245 
vC = 14'b1111110010110110; // vC= -842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001101; // iC=-1331 
vC = 14'b1111110100001011; // vC= -757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110101; // iC=-1291 
vC = 14'b1111110100010001; // vC= -751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110001; // iC=-1359 
vC = 14'b1111110011001110; // vC= -818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000100; // iC=-1212 
vC = 14'b1111110010100001; // vC= -863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111011; // iC=-1285 
vC = 14'b1111110010100101; // vC= -859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011011; // iC=-1317 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001100; // iC=-1204 
vC = 14'b1111110010110111; // vC= -841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b1111110010100000; // vC= -864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b1111110010001100; // vC= -884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101011; // iC=-1237 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011100; // iC=-1316 
vC = 14'b1111110100001011; // vC= -757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100100; // iC=-1308 
vC = 14'b1111110001111110; // vC= -898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110001; // iC=-1295 
vC = 14'b1111110011010110; // vC= -810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001011; // iC=-1205 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111011; // iC=-1285 
vC = 14'b1111110001101101; // vC= -915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010100; // iC=-1196 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101101; // iC=-1299 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111001; // iC=-1287 
vC = 14'b1111110011010011; // vC= -813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110110; // iC=-1290 
vC = 14'b1111110010001000; // vC= -888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010010; // iC=-1262 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b1111110010001100; // vC= -884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110001; // iC=-1231 
vC = 14'b1111110010000011; // vC= -893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000001; // iC=-1279 
vC = 14'b1111110010100110; // vC= -858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100000; // iC=-1184 
vC = 14'b1111110001000111; // vC= -953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001011; // iC=-1205 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001000; // iC=-1208 
vC = 14'b1111110010010101; // vC= -875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000011; // iC=-1149 
vC = 14'b1111110001110110; // vC= -906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100001; // iC=-1119 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111100; // iC=-1220 
vC = 14'b1111110010000100; // vC= -892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011100; // iC=-1124 
vC = 14'b1111110001111010; // vC= -902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111010; // iC=-1222 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001011; // iC=-1205 
vC = 14'b1111110000111001; // vC= -967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100110; // iC=-1114 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010110; // iC=-1194 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000000; // iC=-1088 
vC = 14'b1111110010101100; // vC= -852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111110; // iC=-1090 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101101; // iC=-1235 
vC = 14'b1111110000100001; // vC= -991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011101; // iC=-1187 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110010; // iC=-1102 
vC = 14'b1111110000110101; // vC= -971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110000; // iC=-1168 
vC = 14'b1111110010000001; // vC= -895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111011; // iC=-1157 
vC = 14'b1111110010010011; // vC= -877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000011; // iC=-1213 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010010; // iC=-1070 
vC = 14'b1111110001110101; // vC= -907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110100; // iC=-1100 
vC = 14'b1111101111101001; // vC=-1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010100; // iC=-1068 
vC = 14'b1111110000011110; // vC= -994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010010; // iC=-1198 
vC = 14'b1111110000010100; // vC=-1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000000; // iC=-1152 
vC = 14'b1111110000111011; // vC= -965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011110; // iC=-1186 
vC = 14'b1111101111100110; // vC=-1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011110; // iC=-1058 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011001; // iC=-1127 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110001; // iC=-1103 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011100; // iC=-1124 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001100; // iC=-1012 
vC = 14'b1111110001011001; // vC= -935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001111; // iC=-1073 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111011; // iC=-1157 
vC = 14'b1111110001010111; // vC= -937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100110; // iC=-1114 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111101; // iC=-1027 
vC = 14'b1111101111011100; // vC=-1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000111; // iC=-1081 
vC = 14'b1111101111110101; // vC=-1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010100; // iC=-1132 
vC = 14'b1111110001001111; // vC= -945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101110; // iC=-1106 
vC = 14'b1111101111010100; // vC=-1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111000; // iC=-1032 
vC = 14'b1111101110111000; // vC=-1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000101; // iC=-1083 
vC = 14'b1111101110101001; // vC=-1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011100; // iC=-1124 
vC = 14'b1111110000101000; // vC= -984 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011110; // iC=-1122 
vC = 14'b1111110000000111; // vC=-1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000001; // iC=-1087 
vC = 14'b1111101110100001; // vC=-1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110110; // iC=-1034 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111101; // iC=-1091 
vC = 14'b1111110000010011; // vC=-1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101010; // iC=-1046 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100111; // iC=-1049 
vC = 14'b1111101110111111; // vC=-1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110100; // iC= -972 
vC = 14'b1111101110001100; // vC=-1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101111; // iC= -977 
vC = 14'b1111101111111010; // vC=-1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011010; // iC= -998 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100111; // iC=-1049 
vC = 14'b1111101111111110; // vC=-1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110110; // iC=-1034 
vC = 14'b1111101111111110; // vC=-1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110011; // iC= -973 
vC = 14'b1111101110111010; // vC=-1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000011; // iC=-1021 
vC = 14'b1111101110110010; // vC=-1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010111; // iC=-1065 
vC = 14'b1111101110101101; // vC=-1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100111; // iC= -985 
vC = 14'b1111101110011001; // vC=-1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101011; // iC=-1045 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111010; // iC= -966 
vC = 14'b1111101111010011; // vC=-1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010001; // iC=-1007 
vC = 14'b1111101110101101; // vC=-1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000010; // iC= -958 
vC = 14'b1111101101100011; // vC=-1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110001; // iC= -975 
vC = 14'b1111101111010111; // vC=-1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101010; // iC= -918 
vC = 14'b1111101111000011; // vC=-1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110101; // iC= -971 
vC = 14'b1111101110010001; // vC=-1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111110; // iC= -898 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000000; // iC= -896 
vC = 14'b1111101110001101; // vC=-1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100001; // iC= -863 
vC = 14'b1111101101111010; // vC=-1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101111; // iC= -977 
vC = 14'b1111101101001100; // vC=-1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001101; // iC= -947 
vC = 14'b1111101111001110; // vC=-1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011011; // iC= -997 
vC = 14'b1111101100111110; // vC=-1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110010; // iC= -910 
vC = 14'b1111101111010001; // vC=-1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110101; // iC= -843 
vC = 14'b1111101110001101; // vC=-1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010100; // iC= -940 
vC = 14'b1111101110000111; // vC=-1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110000; // iC= -912 
vC = 14'b1111101110000011; // vC=-1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010011; // iC= -877 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001001; // iC= -887 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110000; // iC= -848 
vC = 14'b1111101110010100; // vC=-1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001011; // iC= -949 
vC = 14'b1111101101111000; // vC=-1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111101; // iC= -835 
vC = 14'b1111101100101100; // vC=-1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101001; // iC= -919 
vC = 14'b1111101101101010; // vC=-1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011100; // iC= -932 
vC = 14'b1111101101111010; // vC=-1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100011; // iC= -925 
vC = 14'b1111101110110100; // vC=-1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011100; // iC= -932 
vC = 14'b1111101110000110; // vC=-1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010000; // iC= -816 
vC = 14'b1111101100100100; // vC=-1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010010; // iC= -878 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111000; // iC= -904 
vC = 14'b1111101101001011; // vC=-1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110010; // iC= -910 
vC = 14'b1111101100010111; // vC=-1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011000; // iC= -872 
vC = 14'b1111101101111100; // vC=-1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010110; // iC= -874 
vC = 14'b1111101100110100; // vC=-1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110011; // iC= -781 
vC = 14'b1111101101000011; // vC=-1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010000; // iC= -880 
vC = 14'b1111101100100100; // vC=-1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110101; // iC= -843 
vC = 14'b1111101110011011; // vC=-1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001011; // iC= -757 
vC = 14'b1111101110010101; // vC=-1131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011000; // iC= -872 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100101; // iC= -859 
vC = 14'b1111101101010110; // vC=-1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100111; // iC= -793 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011001; // iC= -807 
vC = 14'b1111101011111011; // vC=-1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101010; // iC= -726 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011010; // iC= -806 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111100; // iC= -836 
vC = 14'b1111101100001101; // vC=-1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000001; // iC= -703 
vC = 14'b1111101011110110; // vC=-1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000000; // iC= -832 
vC = 14'b1111101101101010; // vC=-1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100101; // iC= -795 
vC = 14'b1111101011111100; // vC=-1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100000; // iC= -736 
vC = 14'b1111101101110110; // vC=-1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100100; // iC= -732 
vC = 14'b1111101011110001; // vC=-1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101110; // iC= -786 
vC = 14'b1111101101010000; // vC=-1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100110; // iC= -730 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110010; // iC= -718 
vC = 14'b1111101100111111; // vC=-1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100010; // iC= -670 
vC = 14'b1111101011001001; // vC=-1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100010; // iC= -798 
vC = 14'b1111101101001100; // vC=-1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011000; // iC= -680 
vC = 14'b1111101100100100; // vC=-1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010110; // iC= -746 
vC = 14'b1111101101001001; // vC=-1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100101; // iC= -731 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011101; // iC= -739 
vC = 14'b1111101011010010; // vC=-1326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111011; // iC= -709 
vC = 14'b1111101101000010; // vC=-1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000100; // iC= -700 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110100; // iC= -652 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001100; // iC= -756 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111010; // iC= -710 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011101; // iC= -675 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001101; // iC= -691 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100100; // iC= -604 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100111; // iC= -665 
vC = 14'b1111101011001101; // vC=-1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001110; // iC= -690 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100111; // iC= -601 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111101011010111; // vC=-1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011110; // iC= -610 
vC = 14'b1111101100100000; // vC=-1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000010; // iC= -702 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101000; // iC= -600 
vC = 14'b1111101010101100; // vC=-1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b1111101010110101; // vC=-1355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110010; // iC= -654 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011100; // iC= -612 
vC = 14'b1111101100101110; // vC=-1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001110; // iC= -562 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110101; // iC= -587 
vC = 14'b1111101100010011; // vC=-1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010101; // iC= -555 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100101; // iC= -539 
vC = 14'b1111101010101010; // vC=-1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111011; // iC= -581 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101111; // iC= -593 
vC = 14'b1111101011100011; // vC=-1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100110; // iC= -602 
vC = 14'b1111101011000011; // vC=-1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011101; // iC= -547 
vC = 14'b1111101011011110; // vC=-1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011110; // iC= -546 
vC = 14'b1111101011110011; // vC=-1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000100; // iC= -508 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110100; // iC= -588 
vC = 14'b1111101010001111; // vC=-1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010001; // iC= -559 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001000; // iC= -504 
vC = 14'b1111101011000010; // vC=-1342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100010; // iC= -478 
vC = 14'b1111101011001001; // vC=-1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001101; // iC= -499 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011010; // iC= -550 
vC = 14'b1111101011011100; // vC=-1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001100; // iC= -500 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110100; // iC= -524 
vC = 14'b1111101100010010; // vC=-1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100101; // iC= -475 
vC = 14'b1111101011010000; // vC=-1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111111; // iC= -513 
vC = 14'b1111101011111111; // vC=-1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100011; // iC= -541 
vC = 14'b1111101010000110; // vC=-1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010011; // iC= -493 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100101; // iC= -539 
vC = 14'b1111101010010010; // vC=-1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101010; // iC= -406 
vC = 14'b1111101001110011; // vC=-1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111010; // iC= -518 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001001; // iC= -439 
vC = 14'b1111101001110100; // vC=-1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100111; // iC= -473 
vC = 14'b1111101011110000; // vC=-1296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000111; // iC= -505 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101111; // iC= -465 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100011; // iC= -413 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011100; // iC= -420 
vC = 14'b1111101010001000; // vC=-1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001001; // iC= -375 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100100; // iC= -348 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111100; // iC= -388 
vC = 14'b1111101010011011; // vC=-1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010010; // iC= -494 
vC = 14'b1111101011010011; // vC=-1325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100111; // iC= -345 
vC = 14'b1111101010001000; // vC=-1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011000; // iC= -360 
vC = 14'b1111101011010101; // vC=-1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000000; // iC= -320 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111010; // iC= -390 
vC = 14'b1111101001111011; // vC=-1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101101; // iC= -403 
vC = 14'b1111101011001111; // vC=-1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101001; // iC= -343 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110001; // iC= -335 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000011; // iC= -445 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111111; // iC= -321 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111001; // iC= -391 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011110; // iC= -354 
vC = 14'b1111101001100100; // vC=-1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011001; // iC= -295 
vC = 14'b1111101010110011; // vC=-1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011000; // iC= -296 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101111; // iC= -337 
vC = 14'b1111101010000000; // vC=-1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110010; // iC= -270 
vC = 14'b1111101001001110; // vC=-1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010110; // iC= -298 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011110; // iC= -226 
vC = 14'b1111101001100111; // vC=-1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101110; // iC= -274 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000000; // iC= -256 
vC = 14'b1111101010111010; // vC=-1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111010; // iC= -198 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000001; // iC= -191 
vC = 14'b1111101001101000; // vC=-1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111001; // iC= -199 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010001; // iC= -239 
vC = 14'b1111101011001000; // vC=-1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111001; // iC= -199 
vC = 14'b1111101011010010; // vC=-1326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110101; // iC= -139 
vC = 14'b1111101001110001; // vC=-1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101100; // iC= -148 
vC = 14'b1111101011011100; // vC=-1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101011; // iC=  -85 
vC = 14'b1111101010101110; // vC=-1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111101; // iC= -195 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001111; // iC= -177 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000110; // iC=  -58 
vC = 14'b1111101010100010; // vC=-1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110111; // iC= -137 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111011; // iC= -133 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100010; // iC=  -30 
vC = 14'b1111101001110100; // vC=-1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001110; // iC=   14 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001110; // iC=  -50 
vC = 14'b1111101011001101; // vC=-1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000001; // iC=  -63 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100111; // iC=  -25 
vC = 14'b1111101011000001; // vC=-1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001101; // iC=   13 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011010; // iC=   26 
vC = 14'b1111101010011011; // vC=-1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011000; // iC=   88 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001001; // iC=   73 
vC = 14'b1111101010110011; // vC=-1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000010; // iC=   66 
vC = 14'b1111101011001110; // vC=-1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001101; // iC=   77 
vC = 14'b1111101011011011; // vC=-1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100011; // iC=  163 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101111; // iC=  111 
vC = 14'b1111101001100111; // vC=-1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101001; // iC=  169 
vC = 14'b1111101010101111; // vC=-1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110111; // iC=  311 
vC = 14'b1111101010110000; // vC=-1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010100; // iC=  276 
vC = 14'b1111101011001010; // vC=-1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010110; // iC=  278 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010111; // iC=  343 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110111; // iC=  375 
vC = 14'b1111101011010000; // vC=-1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100100; // iC=  292 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001001; // iC=  329 
vC = 14'b1111101001110000; // vC=-1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100001; // iC=  353 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110101; // iC=  373 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011010; // iC=  410 
vC = 14'b1111101001111101; // vC=-1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101011; // iC=  427 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110000; // iC=  560 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001011; // iC=  459 
vC = 14'b1111101011001110; // vC=-1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101000; // iC=  552 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111011; // iC=  571 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000110; // iC=  518 
vC = 14'b1111101001101100; // vC=-1428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000010; // iC=  642 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110001; // iC=  689 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101111; // iC=  687 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100101; // iC=  613 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010011; // iC=  723 
vC = 14'b1111101010100111; // vC=-1369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011001; // iC=  793 
vC = 14'b1111101001101110; // vC=-1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011101; // iC=  733 
vC = 14'b1111101001101010; // vC=-1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101011; // iC=  811 
vC = 14'b1111101010011011; // vC=-1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110101; // iC=  821 
vC = 14'b1111101011100111; // vC=-1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011101; // iC=  861 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011001; // iC=  793 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110100; // iC=  820 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111001; // iC=  825 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101100; // iC=  876 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000101; // iC=  965 
vC = 14'b1111101010000010; // vC=-1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110001; // iC= 1009 
vC = 14'b1111101011111001; // vC=-1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011101; // iC=  925 
vC = 14'b1111101011000001; // vC=-1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010100; // iC=  916 
vC = 14'b1111101010101111; // vC=-1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101111; // iC= 1071 
vC = 14'b1111101100000111; // vC=-1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111000; // iC= 1016 
vC = 14'b1111101100010010; // vC=-1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101011; // iC= 1131 
vC = 14'b1111101010100010; // vC=-1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000010; // iC= 1154 
vC = 14'b1111101011110100; // vC=-1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111010; // iC= 1082 
vC = 14'b1111101010100100; // vC=-1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100101; // iC= 1061 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100000; // iC= 1120 
vC = 14'b1111101100010100; // vC=-1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011010; // iC= 1114 
vC = 14'b1111101011001010; // vC=-1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011111; // iC= 1183 
vC = 14'b1111101011010000; // vC=-1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010010; // iC= 1170 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011101; // iC= 1245 
vC = 14'b1111101011101110; // vC=-1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001000; // iC= 1224 
vC = 14'b1111101011011110; // vC=-1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101100; // iC= 1260 
vC = 14'b1111101100110101; // vC=-1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111011; // iC= 1211 
vC = 14'b1111101011011001; // vC=-1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111100; // iC= 1340 
vC = 14'b1111101100011000; // vC=-1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110101; // iC= 1333 
vC = 14'b1111101100111110; // vC=-1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111110; // iC= 1278 
vC = 14'b1111101011111101; // vC=-1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100110; // iC= 1382 
vC = 14'b1111101100111100; // vC=-1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101000; // iC= 1320 
vC = 14'b1111101101010001; // vC=-1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100110; // iC= 1446 
vC = 14'b1111101100001100; // vC=-1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111111; // iC= 1343 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000110; // iC= 1478 
vC = 14'b1111101100101111; // vC=-1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001101; // iC= 1421 
vC = 14'b1111101100011001; // vC=-1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101100; // iC= 1388 
vC = 14'b1111101101011100; // vC=-1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010111; // iC= 1495 
vC = 14'b1111101101111001; // vC=-1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110110; // iC= 1398 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110110; // iC= 1526 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000010; // iC= 1538 
vC = 14'b1111101100100101; // vC=-1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101011; // iC= 1515 
vC = 14'b1111101101101110; // vC=-1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111011; // iC= 1595 
vC = 14'b1111101110001110; // vC=-1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110111; // iC= 1591 
vC = 14'b1111101101101001; // vC=-1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000111; // iC= 1479 
vC = 14'b1111101101011101; // vC=-1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b1111101101101000; // vC=-1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111011; // iC= 1531 
vC = 14'b1111101110000011; // vC=-1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101111; // iC= 1583 
vC = 14'b1111101101100110; // vC=-1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011010; // iC= 1626 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001011; // iC= 1675 
vC = 14'b1111101110101110; // vC=-1106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b1111101111001010; // vC=-1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100100; // iC= 1636 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b1111101110001001; // vC=-1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b1111101110011111; // vC=-1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000001; // iC= 1729 
vC = 14'b1111101101101100; // vC=-1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011010; // iC= 1626 
vC = 14'b1111101111101001; // vC=-1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b1111101111111100; // vC=-1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011100; // iC= 1628 
vC = 14'b1111101110011100; // vC=-1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100111; // iC= 1639 
vC = 14'b1111101111101001; // vC=-1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101001; // iC= 1705 
vC = 14'b1111101110110010; // vC=-1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010101; // iC= 1749 
vC = 14'b1111101111111011; // vC=-1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001000; // iC= 1672 
vC = 14'b1111101111010110; // vC=-1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110001; // iC= 1777 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b1111110000100101; // vC= -987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110101; // iC= 1781 
vC = 14'b1111101110100101; // vC=-1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101101; // iC= 1709 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100100; // iC= 1764 
vC = 14'b1111101110101111; // vC=-1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b1111110000000001; // vC=-1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000111; // iC= 1799 
vC = 14'b1111110000110001; // vC= -975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001010; // iC= 1738 
vC = 14'b1111110000001101; // vC=-1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b1111101111101111; // vC=-1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110001; // iC= 1777 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101101; // iC= 1837 
vC = 14'b1111101111110110; // vC=-1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001011; // iC= 1739 
vC = 14'b1111110001100000; // vC= -928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111101111111110; // vC=-1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b1111110001010101; // vC= -939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011110; // iC= 1886 
vC = 14'b1111110001110110; // vC= -906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b1111110010000001; // vC= -895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101100; // iC= 1772 
vC = 14'b1111110010000101; // vC= -891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001001; // iC= 1865 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011111; // iC= 1759 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011000; // iC= 1880 
vC = 14'b1111110000000011; // vC=-1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b1111110000101010; // vC= -982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b1111110001110110; // vC= -906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111110001011111; // vC= -929 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b1111110000111110; // vC= -962 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b1111110010000101; // vC= -891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b1111110011001110; // vC= -818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b1111110011010011; // vC= -813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100110; // iC= 1830 
vC = 14'b1111110001101111; // vC= -913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111110010111010; // vC= -838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b1111110010101101; // vC= -851 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b1111110011011111; // vC= -801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111110011100111; // vC= -793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011100; // iC= 1820 
vC = 14'b1111110011110101; // vC= -779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b1111110100101010; // vC= -726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111110011010001; // vC= -815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010011; // iC= 1811 
vC = 14'b1111110100011011; // vC= -741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011000; // iC= 1880 
vC = 14'b1111110011001001; // vC= -823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b1111110011101000; // vC= -792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b1111110101010000; // vC= -688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111110100001000; // vC= -760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101101; // iC= 1837 
vC = 14'b1111110100000001; // vC= -767 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111110100100011; // vC= -733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111110011111010; // vC= -774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111110101001001; // vC= -695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110100111001; // vC= -711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111110101010010; // vC= -686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111110100100011; // vC= -733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b1111110101001000; // vC= -696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001000; // iC= 1864 
vC = 14'b1111110100100011; // vC= -733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111110101100010; // vC= -670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100110; // iC= 1830 
vC = 14'b1111110101101010; // vC= -662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b1111110110011011; // vC= -613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111110110110001; // vC= -591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110100111110; // vC= -706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b1111110101111011; // vC= -645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110110010001; // vC= -623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b1111110110111011; // vC= -581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000101; // iC= 1861 
vC = 14'b1111110111010101; // vC= -555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b1111110110111011; // vC= -581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111110101100001; // vC= -671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000100; // iC= 1860 
vC = 14'b1111110111101101; // vC= -531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101010; // iC= 1898 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b1111110110111000; // vC= -584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001001; // iC= 1865 
vC = 14'b1111110110011100; // vC= -612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b1111110111100111; // vC= -537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111110111101011; // vC= -533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b1111110110010011; // vC= -621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111110110011001; // vC= -615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111110110001011; // vC= -629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111110110101111; // vC= -593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011100; // iC= 1884 
vC = 14'b1111110110101101; // vC= -595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b1111110111101110; // vC= -530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b1111110111101110; // vC= -530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b1111110111000011; // vC= -573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b1111111000111010; // vC= -454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110110110101; // vC= -587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111111000000000; // vC= -512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111101; // iC= 1853 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111111001100011; // vC= -413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111111001011110; // vC= -418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010010; // iC= 1874 
vC = 14'b1111111001111000; // vC= -392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b1111110111110111; // vC= -521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b1111111000100011; // vC= -477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111011; // iC= 1851 
vC = 14'b1111110111110000; // vC= -528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111110111110010; // vC= -526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111111001100100; // vC= -412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111111000011100; // vC= -484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b1111111000100000; // vC= -480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111111001001111; // vC= -433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b1111111000110000; // vC= -464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111111010100010; // vC= -350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111010110001; // vC= -335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111111010100110; // vC= -346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111111011001011; // vC= -309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b1111111010111100; // vC= -324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b1111111001101111; // vC= -401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111111010110111; // vC= -329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000101; // iC= 1861 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111111001101100; // vC= -404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111111010001100; // vC= -372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111111011011111; // vC= -289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111010101001; // vC= -343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b1111111010111110; // vC= -322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b1111111010101000; // vC= -344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001101; // iC= 1869 
vC = 14'b1111111100001100; // vC= -244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b1111111011100001; // vC= -287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001010; // iC= 1866 
vC = 14'b1111111011101011; // vC= -277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001101; // iC= 1869 
vC = 14'b1111111100010001; // vC= -239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111100010011; // vC= -237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b1111111100111000; // vC= -200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b1111111100111011; // vC= -197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b1111111100111000; // vC= -200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b1111111011000010; // vC= -318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b1111111101010001; // vC= -175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111111100000100; // vC= -252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b1111111100101111; // vC= -209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110110; // iC= 1846 
vC = 14'b1111111101100010; // vC= -158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111111101001111; // vC= -177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b1111111101101001; // vC= -151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011000; // iC= 1880 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111111100110000; // vC= -208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b1111111101011001; // vC= -167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111111100111011; // vC= -197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111100101010; // vC= -214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111001; // iC= 1849 
vC = 14'b1111111110000001; // vC= -127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b1111111110110000; // vC=  -80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b1111111110001110; // vC= -114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b1111111110011110; // vC=  -98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111111101000011; // vC= -189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b1111111111001110; // vC=  -50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b1111111101011000; // vC= -168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b1111111111100111; // vC=  -25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b1111111101010100; // vC= -172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b1111111101101000; // vC= -152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b1111111110110100; // vC=  -76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111111111100011; // vC=  -29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111111111011011; // vC=  -37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010001; // iC= 1873 
vC = 14'b1111111110001111; // vC= -113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111111110101011; // vC=  -85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b1111111110111001; // vC=  -71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b1111111110110110; // vC=  -74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111111111011010; // vC=  -38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b1111111111001110; // vC=  -50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b0000000000001011; // vC=   11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111111111011101; // vC=  -35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b0000000000011101; // vC=   29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b0000000000100000; // vC=   32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b0000000000101011; // vC=   43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b0000000001011101; // vC=   93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b1111111111001100; // vC=  -52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b0000000001101100; // vC=  108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111001; // iC= 1849 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111111111110001; // vC=  -15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b0000000001100111; // vC=  103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b0000000000010011; // vC=   19 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b0000000000001001; // vC=    9 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b0000000000100000; // vC=   32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101111; // iC= 1839 
vC = 14'b0000000000110100; // vC=   52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100011; // iC= 1827 
vC = 14'b0000000000100001; // vC=   33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010000; // iC= 1808 
vC = 14'b0000000000100011; // vC=   35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b0000000010001011; // vC=  139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101001; // iC= 1833 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011001; // iC= 1881 
vC = 14'b0000000010001010; // vC=  138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b0000000010101010; // vC=  170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b0000000001111001; // vC=  121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000100; // iC= 1796 
vC = 14'b0000000010000001; // vC=  129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101001; // iC= 1833 
vC = 14'b0000000001100111; // vC=  103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110111; // iC= 1783 
vC = 14'b0000000010111110; // vC=  190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b0000000011111100; // vC=  252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b0000000011001111; // vC=  207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b0000000011010011; // vC=  211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111110; // iC= 1790 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b0000000100100010; // vC=  290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b0000000100010001; // vC=  273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b0000000101001101; // vC=  333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b0000000100111011; // vC=  315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b0000000100010010; // vC=  274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b0000000101001011; // vC=  331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000000; // iC= 1792 
vC = 14'b0000000101100000; // vC=  352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b0000000101000001; // vC=  321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011100; // iC= 1884 
vC = 14'b0000000011101101; // vC=  237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b0000000110000001; // vC=  385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001000; // iC= 1864 
vC = 14'b0000000101101010; // vC=  362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010111; // iC= 1751 
vC = 14'b0000000100111111; // vC=  319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b0000000100010100; // vC=  276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111101; // iC= 1853 
vC = 14'b0000000100110101; // vC=  309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111101; // iC= 1853 
vC = 14'b0000000100011100; // vC=  284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b0000000101100001; // vC=  353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b0000000100100110; // vC=  294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110010; // iC= 1778 
vC = 14'b0000000100111001; // vC=  313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b0000000101101100; // vC=  364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001011; // iC= 1739 
vC = 14'b0000000100101001; // vC=  297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100011; // iC= 1763 
vC = 14'b0000000101101100; // vC=  364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b0000000111010100; // vC=  468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100010; // iC= 1826 
vC = 14'b0000000110101101; // vC=  429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b0000000101000011; // vC=  323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b0000000101101010; // vC=  362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101111; // iC= 1839 
vC = 14'b0000000110100011; // vC=  419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b0000000110011010; // vC=  410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000000101101101; // vC=  365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101101; // iC= 1709 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b0000000110101000; // vC=  424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b0000000110101001; // vC=  425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101011; // iC= 1707 
vC = 14'b0000000111011111; // vC=  479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101101; // iC= 1837 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011111; // iC= 1759 
vC = 14'b0000001000000111; // vC=  519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b0000000110111000; // vC=  440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000011; // iC= 1795 
vC = 14'b0000000110011000; // vC=  408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b0000000111001000; // vC=  456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010011; // iC= 1811 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100000; // iC= 1824 
vC = 14'b0000000111111110; // vC=  510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b0000000111101011; // vC=  491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000001000110100; // vC=  564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001001; // iC= 1737 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b0000001000011101; // vC=  541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b0000000111010000; // vC=  464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000001001010101; // vC=  597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b0000001001010001; // vC=  593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011101; // iC= 1693 
vC = 14'b0000000111010001; // vC=  465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000100; // iC= 1668 
vC = 14'b0000000111011111; // vC=  479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b0000001001001110; // vC=  590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110010; // iC= 1650 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b0000001001011111; // vC=  607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b0000001000100001; // vC=  545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b0000001000000111; // vC=  519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001101; // iC= 1677 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010101; // iC= 1685 
vC = 14'b0000001000010011; // vC=  531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001011; // iC= 1675 
vC = 14'b0000001000111011; // vC=  571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011000; // iC= 1688 
vC = 14'b0000001001011101; // vC=  605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b0000001000111100; // vC=  572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010100; // iC= 1620 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100010; // iC= 1634 
vC = 14'b0000001001111101; // vC=  637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b0000001010011011; // vC=  667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001111; // iC= 1615 
vC = 14'b0000001001001110; // vC=  590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b0000001000111100; // vC=  572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100011; // iC= 1699 
vC = 14'b0000001010000111; // vC=  647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001001; // iC= 1609 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b0000001001110010; // vC=  626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001110; // iC= 1742 
vC = 14'b0000001001011011; // vC=  603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110000; // iC= 1584 
vC = 14'b0000001001101100; // vC=  620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011000; // iC= 1688 
vC = 14'b0000001011011111; // vC=  735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b0000001001101110; // vC=  622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010010; // iC= 1682 
vC = 14'b0000001010001110; // vC=  654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100100; // iC= 1636 
vC = 14'b0000001100000011; // vC=  771 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011011; // iC= 1563 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b0000001010011100; // vC=  668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100001; // iC= 1697 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101011; // iC= 1643 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101101; // iC= 1645 
vC = 14'b0000001010110001; // vC=  689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100001; // iC= 1697 
vC = 14'b0000001011011101; // vC=  733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000100; // iC= 1668 
vC = 14'b0000001010100111; // vC=  679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011101; // iC= 1629 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b0000001011100111; // vC=  743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100110; // iC= 1638 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110001; // iC= 1649 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001111; // iC= 1551 
vC = 14'b0000001100110010; // vC=  818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101001; // iC= 1641 
vC = 14'b0000001100110111; // vC=  823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010001; // iC= 1553 
vC = 14'b0000001011100101; // vC=  741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011010; // iC= 1626 
vC = 14'b0000001011100011; // vC=  739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001000; // iC= 1544 
vC = 14'b0000001101000001; // vC=  833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101110; // iC= 1582 
vC = 14'b0000001011011000; // vC=  728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100100; // iC= 1636 
vC = 14'b0000001011101101; // vC=  749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010110; // iC= 1558 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010100; // iC= 1556 
vC = 14'b0000001101110010; // vC=  882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011011; // iC= 1499 
vC = 14'b0000001101011001; // vC=  857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101000; // iC= 1512 
vC = 14'b0000001101100111; // vC=  871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100011; // iC= 1507 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110110; // iC= 1526 
vC = 14'b0000001100110101; // vC=  821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110101; // iC= 1589 
vC = 14'b0000001100001010; // vC=  778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010100; // iC= 1492 
vC = 14'b0000001101011011; // vC=  859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111011; // iC= 1531 
vC = 14'b0000001100011111; // vC=  799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010111; // iC= 1559 
vC = 14'b0000001101101111; // vC=  879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001100; // iC= 1484 
vC = 14'b0000001101101010; // vC=  874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111101; // iC= 1597 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001111; // iC= 1551 
vC = 14'b0000001100110001; // vC=  817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001011; // iC= 1611 
vC = 14'b0000001101010001; // vC=  849 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011000; // iC= 1496 
vC = 14'b0000001110111011; // vC=  955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010100; // iC= 1492 
vC = 14'b0000001110101100; // vC=  940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100010; // iC= 1506 
vC = 14'b0000001110100110; // vC=  934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b0000001101010000; // vC=  848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b0000001110101110; // vC=  942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110010; // iC= 1458 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011010; // iC= 1434 
vC = 14'b0000001101110011; // vC=  883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100111; // iC= 1447 
vC = 14'b0000001101000110; // vC=  838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010000; // iC= 1488 
vC = 14'b0000001101100101; // vC=  869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011110; // iC= 1502 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111010; // iC= 1530 
vC = 14'b0000001110101011; // vC=  939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101010; // iC= 1514 
vC = 14'b0000001101101101; // vC=  877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110111; // iC= 1527 
vC = 14'b0000001110101111; // vC=  943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000110; // iC= 1542 
vC = 14'b0000001101110001; // vC=  881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111010; // iC= 1466 
vC = 14'b0000001111100100; // vC=  996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101001; // iC= 1449 
vC = 14'b0000001101110111; // vC=  887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b0000001110010011; // vC=  915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000101; // iC= 1477 
vC = 14'b0000001111101110; // vC= 1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011101; // iC= 1437 
vC = 14'b0000001111100011; // vC=  995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011001; // iC= 1497 
vC = 14'b0000001111100010; // vC=  994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110010; // iC= 1458 
vC = 14'b0000001110001010; // vC=  906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011001; // iC= 1497 
vC = 14'b0000001110111011; // vC=  955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011100; // iC= 1436 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011101; // iC= 1437 
vC = 14'b0000001111010101; // vC=  981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010110; // iC= 1430 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000101; // iC= 1413 
vC = 14'b0000010000100011; // vC= 1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001001; // iC= 1353 
vC = 14'b0000001110110001; // vC=  945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000010; // iC= 1410 
vC = 14'b0000010000100110; // vC= 1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001100; // iC= 1420 
vC = 14'b0000001110111011; // vC=  955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101011; // iC= 1387 
vC = 14'b0000010000110111; // vC= 1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101001; // iC= 1385 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101001; // iC= 1449 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010001; // iC= 1425 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101100; // iC= 1388 
vC = 14'b0000010001011010; // vC= 1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001000; // iC= 1352 
vC = 14'b0000010000101110; // vC= 1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100110; // iC= 1318 
vC = 14'b0000001111001100; // vC=  972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101110; // iC= 1454 
vC = 14'b0000010000110100; // vC= 1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110010; // iC= 1394 
vC = 14'b0000010000100011; // vC= 1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000111; // iC= 1415 
vC = 14'b0000001111111001; // vC= 1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010011; // iC= 1299 
vC = 14'b0000010000000111; // vC= 1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011111; // iC= 1311 
vC = 14'b0000010001100001; // vC= 1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011011; // iC= 1371 
vC = 14'b0000010000101110; // vC= 1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011010; // iC= 1370 
vC = 14'b0000001111101000; // vC= 1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101100; // iC= 1388 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010010; // iC= 1362 
vC = 14'b0000001111101110; // vC= 1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000001; // iC= 1345 
vC = 14'b0000001111111100; // vC= 1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111010; // iC= 1274 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101101; // iC= 1389 
vC = 14'b0000010001000101; // vC= 1093 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000011; // iC= 1411 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101001; // iC= 1257 
vC = 14'b0000010001010011; // vC= 1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100101; // iC= 1317 
vC = 14'b0000010001011010; // vC= 1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101111; // iC= 1327 
vC = 14'b0000010000001010; // vC= 1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110011; // iC= 1267 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101000; // iC= 1384 
vC = 14'b0000010001000001; // vC= 1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010101; // iC= 1365 
vC = 14'b0000010001101001; // vC= 1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010010; // iC= 1298 
vC = 14'b0000010001111001; // vC= 1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000100; // iC= 1284 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011011; // iC= 1243 
vC = 14'b0000010001111010; // vC= 1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100100; // iC= 1252 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000100; // iC= 1284 
vC = 14'b0000010001000000; // vC= 1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001110; // iC= 1230 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101110; // iC= 1326 
vC = 14'b0000010010010110; // vC= 1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100101; // iC= 1253 
vC = 14'b0000010001000101; // vC= 1093 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111000; // iC= 1208 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000001; // iC= 1281 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101010; // iC= 1322 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011101; // iC= 1245 
vC = 14'b0000010001010110; // vC= 1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010110; // iC= 1174 
vC = 14'b0000010010101100; // vC= 1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001101; // iC= 1229 
vC = 14'b0000010011101001; // vC= 1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110010; // iC= 1202 
vC = 14'b0000010010000001; // vC= 1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100000; // iC= 1184 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111101; // iC= 1149 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000000; // iC= 1280 
vC = 14'b0000010010011110; // vC= 1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011011; // iC= 1179 
vC = 14'b0000010001111011; // vC= 1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111111; // iC= 1279 
vC = 14'b0000010001101011; // vC= 1131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000100; // iC= 1284 
vC = 14'b0000010100001000; // vC= 1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011101; // iC= 1245 
vC = 14'b0000010011001011; // vC= 1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111011; // iC= 1275 
vC = 14'b0000010010100101; // vC= 1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100101; // iC= 1189 
vC = 14'b0000010100001111; // vC= 1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110011; // iC= 1203 
vC = 14'b0000010100000101; // vC= 1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001010; // iC= 1162 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001110; // iC= 1230 
vC = 14'b0000010010001001; // vC= 1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001100; // iC= 1164 
vC = 14'b0000010010001111; // vC= 1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011101; // iC= 1245 
vC = 14'b0000010011111000; // vC= 1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000011; // iC= 1091 
vC = 14'b0000010100000111; // vC= 1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010111; // iC= 1239 
vC = 14'b0000010100000101; // vC= 1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010100; // iC= 1108 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101011; // iC= 1131 
vC = 14'b0000010010010100; // vC= 1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111101; // iC= 1149 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b0000010011111100; // vC= 1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101111; // iC= 1071 
vC = 14'b0000010010100101; // vC= 1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b0000010011010000; // vC= 1232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010011; // iC= 1107 
vC = 14'b0000010010110001; // vC= 1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011001; // iC= 1049 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001100; // iC= 1100 
vC = 14'b0000010011000001; // vC= 1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111011; // iC= 1147 
vC = 14'b0000010011000010; // vC= 1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101010; // iC= 1130 
vC = 14'b0000010011111011; // vC= 1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001010; // iC= 1098 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000101; // iC= 1029 
vC = 14'b0000010011100100; // vC= 1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101000; // iC= 1064 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111011; // iC= 1083 
vC = 14'b0000010011001110; // vC= 1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011101; // iC= 1053 
vC = 14'b0000010011001001; // vC= 1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000000; // iC= 1024 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101110; // iC= 1006 
vC = 14'b0000010101001010; // vC= 1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101100; // iC= 1068 
vC = 14'b0000010011110111; // vC= 1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110010; // iC= 1074 
vC = 14'b0000010101000111; // vC= 1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111001; // iC= 1081 
vC = 14'b0000010100110011; // vC= 1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100011; // iC= 1059 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101000; // iC= 1000 
vC = 14'b0000010100000001; // vC= 1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101000; // iC= 1000 
vC = 14'b0000010100001010; // vC= 1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110111; // iC= 1015 
vC = 14'b0000010100011001; // vC= 1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001100; // iC= 1100 
vC = 14'b0000010101100000; // vC= 1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000001; // iC=  961 
vC = 14'b0000010100011000; // vC= 1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001111; // iC= 1103 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111101; // iC= 1085 
vC = 14'b0000010100111110; // vC= 1342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110000; // iC= 1008 
vC = 14'b0000010101101011; // vC= 1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001101; // iC=  973 
vC = 14'b0000010101010110; // vC= 1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011011; // iC=  987 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101110; // iC=  942 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101110; // iC= 1006 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110111; // iC=  951 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100011; // iC= 1059 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001000; // iC= 1032 
vC = 14'b0000010110100000; // vC= 1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111011; // iC= 1019 
vC = 14'b0000010110001110; // vC= 1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110111; // iC= 1015 
vC = 14'b0000010100011100; // vC= 1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111111; // iC= 1023 
vC = 14'b0000010110010001; // vC= 1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100001; // iC=  929 
vC = 14'b0000010110011000; // vC= 1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101100; // iC=  876 
vC = 14'b0000010100110001; // vC= 1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100110; // iC=  870 
vC = 14'b0000010110110011; // vC= 1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011011; // iC=  987 
vC = 14'b0000010101101111; // vC= 1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011100; // iC=  860 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001000; // iC=  968 
vC = 14'b0000010100110001; // vC= 1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111010; // iC=  890 
vC = 14'b0000010110111111; // vC= 1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000110; // iC=  966 
vC = 14'b0000010111000100; // vC= 1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101101; // iC=  877 
vC = 14'b0000010110010110; // vC= 1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111011; // iC=  891 
vC = 14'b0000010101110001; // vC= 1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000101; // iC=  901 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111011; // iC=  827 
vC = 14'b0000010111010000; // vC= 1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101000; // iC=  936 
vC = 14'b0000010110001100; // vC= 1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101011; // iC=  811 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110011; // iC=  819 
vC = 14'b0000010110000001; // vC= 1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110011; // iC=  819 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110110; // iC=  886 
vC = 14'b0000010110110100; // vC= 1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101100; // iC=  940 
vC = 14'b0000010110010101; // vC= 1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101001; // iC=  937 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100000; // iC=  800 
vC = 14'b0000010101001011; // vC= 1355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100000; // iC=  864 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011001; // iC=  793 
vC = 14'b0000010110000010; // vC= 1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001011; // iC=  779 
vC = 14'b0000010111001011; // vC= 1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110010; // iC=  882 
vC = 14'b0000010101100111; // vC= 1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001010; // iC=  778 
vC = 14'b0000010111001010; // vC= 1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000001; // iC=  897 
vC = 14'b0000010101100010; // vC= 1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101001; // iC=  809 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010010; // iC=  850 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001111; // iC=  783 
vC = 14'b0000010110110111; // vC= 1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011010; // iC=  858 
vC = 14'b0000010110101101; // vC= 1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000011; // iC=  771 
vC = 14'b0000010101111101; // vC= 1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010100; // iC=  724 
vC = 14'b0000010110000101; // vC= 1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110010; // iC=  818 
vC = 14'b0000010110110100; // vC= 1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110010; // iC=  818 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111000; // iC=  824 
vC = 14'b0000010110110111; // vC= 1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001010; // iC=  778 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001010; // iC=  842 
vC = 14'b0000010111110010; // vC= 1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001011; // iC=  779 
vC = 14'b0000010110010100; // vC= 1428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110111; // iC=  823 
vC = 14'b0000010110101001; // vC= 1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011110; // iC=  734 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101011; // iC=  811 
vC = 14'b0000011000010011; // vC= 1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000101; // iC=  773 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100111; // iC=  679 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011110; // iC=  798 
vC = 14'b0000010110101001; // vC= 1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101111; // iC=  687 
vC = 14'b0000010110110000; // vC= 1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001000; // iC=  712 
vC = 14'b0000010111101100; // vC= 1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b0000010110110010; // vC= 1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111111; // iC=  767 
vC = 14'b0000010110111001; // vC= 1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101011; // iC=  747 
vC = 14'b0000010111000100; // vC= 1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101100; // iC=  684 
vC = 14'b0000010111111001; // vC= 1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110000; // iC=  752 
vC = 14'b0000010110011111; // vC= 1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010010; // iC=  722 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101111; // iC=  751 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010101; // iC=  725 
vC = 14'b0000010111000010; // vC= 1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001110; // iC=  590 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101100; // iC=  620 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110010; // iC=  690 
vC = 14'b0000010111111111; // vC= 1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010000; // iC=  592 
vC = 14'b0000010111111110; // vC= 1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011011; // iC=  667 
vC = 14'b0000011000011001; // vC= 1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011011; // iC=  603 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100111; // iC=  615 
vC = 14'b0000010111011100; // vC= 1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100001; // iC=  673 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111011; // iC=  699 
vC = 14'b0000010111011011; // vC= 1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101100; // iC=  620 
vC = 14'b0000010110101101; // vC= 1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011111; // iC=  543 
vC = 14'b0000010110101001; // vC= 1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100000; // iC=  672 
vC = 14'b0000010111000100; // vC= 1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110001; // iC=  561 
vC = 14'b0000010110100000; // vC= 1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101000; // iC=  616 
vC = 14'b0000011000001001; // vC= 1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111111; // iC=  639 
vC = 14'b0000010110110110; // vC= 1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011011; // iC=  603 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000100; // iC=  516 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101000; // iC=  616 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101100; // iC=  556 
vC = 14'b0000010111010111; // vC= 1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111010; // iC=  634 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110100; // iC=  628 
vC = 14'b0000010111110111; // vC= 1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110110; // iC=  630 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101101; // iC=  493 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000111; // iC=  583 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001111; // iC=  591 
vC = 14'b0000010111100100; // vC= 1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011010; // iC=  602 
vC = 14'b0000011000101101; // vC= 1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111010; // iC=  570 
vC = 14'b0000011001010101; // vC= 1621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010010; // iC=  594 
vC = 14'b0000010111011100; // vC= 1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010111; // iC=  535 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101010; // iC=  426 
vC = 14'b0000010111110010; // vC= 1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110111; // iC=  567 
vC = 14'b0000011000111110; // vC= 1598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000011; // iC=  451 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010111; // iC=  471 
vC = 14'b0000010111000000; // vC= 1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000011; // iC=  451 
vC = 14'b0000010111011000; // vC= 1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111100; // iC=  508 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000010; // iC=  386 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000110; // iC=  518 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010011; // iC=  467 
vC = 14'b0000011000001001; // vC= 1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010101; // iC=  405 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011110; // iC=  414 
vC = 14'b0000010111100011; // vC= 1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100101; // iC=  421 
vC = 14'b0000010111111111; // vC= 1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011110; // iC=  350 
vC = 14'b0000010111011110; // vC= 1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010010; // iC=  466 
vC = 14'b0000010111011100; // vC= 1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111110; // iC=  318 
vC = 14'b0000010111110010; // vC= 1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011011; // iC=  347 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100000; // iC=  352 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000010; // iC=  322 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101110; // iC=  366 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000000; // iC=  384 
vC = 14'b0000011001001110; // vC= 1614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101001; // iC=  233 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100010; // iC=  290 
vC = 14'b0000011001100110; // vC= 1638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110110; // iC=  246 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100001; // iC=  289 
vC = 14'b0000011001011001; // vC= 1625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111100; // iC=  316 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111001; // iC=  185 
vC = 14'b0000011001100101; // vC= 1637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010010; // iC=  274 
vC = 14'b0000010111110001; // vC= 1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001101; // iC=  141 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111001; // iC=  121 
vC = 14'b0000010111011101; // vC= 1501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000000; // iC=  128 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111001; // iC=  121 
vC = 14'b0000011001011000; // vC= 1624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100100; // iC=  164 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000001; // iC=  193 
vC = 14'b0000010111111111; // vC= 1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010111; // iC=  151 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010010; // iC=   82 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000101; // iC=    5 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001000; // iC=  136 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011011; // iC=   27 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010101; // iC=   85 
vC = 14'b0000010111110101; // vC= 1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010111; // iC=   23 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100010; // iC=   34 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110011; // iC=  -77 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001000; // iC= -120 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010100; // iC=  -44 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111010; // iC=   -6 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101000; // iC=  -24 
vC = 14'b0000011000101010; // vC= 1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001100; // iC= -180 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111100; // iC= -132 
vC = 14'b0000011001010001; // vC= 1617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010010; // iC= -238 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111111; // iC= -193 
vC = 14'b0000011001000001; // vC= 1601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111110; // iC= -130 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000100; // iC= -252 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110010; // iC= -334 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100000; // iC= -352 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111111; // iC= -321 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011111; // iC= -353 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011100; // iC= -356 
vC = 14'b0000010111101001; // vC= 1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101101; // iC= -339 
vC = 14'b0000011000010010; // vC= 1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110110; // iC= -394 
vC = 14'b0000011001001100; // vC= 1612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010000; // iC= -432 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101010; // iC= -406 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110000; // iC= -464 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010011; // iC= -429 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000011; // iC= -509 
vC = 14'b0000010111010011; // vC= 1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110101; // iC= -523 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100110; // iC= -602 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011001; // iC= -487 
vC = 14'b0000010111110011; // vC= 1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000010; // iC= -574 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011010; // iC= -550 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111100; // iC= -644 
vC = 14'b0000010111010000; // vC= 1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001010; // iC= -630 
vC = 14'b0000011000110001; // vC= 1585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111010; // iC= -646 
vC = 14'b0000010111011001; // vC= 1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000000; // iC= -768 
vC = 14'b0000011000101101; // vC= 1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111101; // iC= -707 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001100; // iC= -756 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110010; // iC= -718 
vC = 14'b0000010111101100; // vC= 1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001101; // iC= -755 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001011; // iC= -821 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011110; // iC= -866 
vC = 14'b0000010110011100; // vC= 1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100111; // iC= -793 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010011; // iC= -813 
vC = 14'b0000010110010011; // vC= 1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010010; // iC= -942 
vC = 14'b0000010111110101; // vC= 1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001010; // iC= -886 
vC = 14'b0000010110111001; // vC= 1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001100; // iC= -884 
vC = 14'b0000010110010101; // vC= 1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001011; // iC= -949 
vC = 14'b0000010111110100; // vC= 1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110011; // iC= -973 
vC = 14'b0000010110010000; // vC= 1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000100; // iC=-1020 
vC = 14'b0000010111111011; // vC= 1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110100; // iC= -972 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011000; // iC=-1000 
vC = 14'b0000010111101011; // vC= 1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001100; // iC=-1076 
vC = 14'b0000010111010110; // vC= 1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111101; // iC= -963 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000010; // iC=-1022 
vC = 14'b0000010101010001; // vC= 1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101110; // iC=-1042 
vC = 14'b0000010111010010; // vC= 1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111010; // iC=-1094 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000011; // iC=-1085 
vC = 14'b0000010101111010; // vC= 1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010110; // iC=-1066 
vC = 14'b0000010101000000; // vC= 1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001001; // iC=-1207 
vC = 14'b0000010100110001; // vC= 1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100011; // iC=-1117 
vC = 14'b0000010101110010; // vC= 1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011101; // iC=-1251 
vC = 14'b0000010100110001; // vC= 1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100100; // iC=-1116 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100111; // iC=-1177 
vC = 14'b0000010110000100; // vC= 1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010111; // iC=-1193 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011110; // iC=-1314 
vC = 14'b0000010100110100; // vC= 1332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001010; // iC=-1334 
vC = 14'b0000010101000111; // vC= 1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011000; // iC=-1320 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101000; // iC=-1304 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111101; // iC=-1283 
vC = 14'b0000010101100001; // vC= 1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100001; // iC=-1375 
vC = 14'b0000010101100101; // vC= 1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100101; // iC=-1371 
vC = 14'b0000010100110111; // vC= 1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000111; // iC=-1401 
vC = 14'b0000010011101101; // vC= 1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b0000010100000111; // vC= 1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101110; // iC=-1362 
vC = 14'b0000010101101011; // vC= 1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111110; // iC=-1346 
vC = 14'b0000010101111001; // vC= 1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100000; // iC=-1312 
vC = 14'b0000010100101001; // vC= 1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b0000010011100000; // vC= 1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010000; // iC=-1392 
vC = 14'b0000010100011101; // vC= 1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000010011110111; // vC= 1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b0000010011011100; // vC= 1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b0000010100000011; // vC= 1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001111; // iC=-1457 
vC = 14'b0000010010110101; // vC= 1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b0000010100010101; // vC= 1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100010; // iC=-1502 
vC = 14'b0000010011100111; // vC= 1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010010; // iC=-1518 
vC = 14'b0000010011110010; // vC= 1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b0000010011100000; // vC= 1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000010010001111; // vC= 1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000010100001111; // vC= 1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011000; // iC=-1512 
vC = 14'b0000010010110111; // vC= 1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000010011111111; // vC= 1279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b0000010011001101; // vC= 1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b0000010001110111; // vC= 1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110100; // iC=-1548 
vC = 14'b0000010011100100; // vC= 1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000010010010011; // vC= 1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b0000010010110111; // vC= 1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b0000010001001000; // vC= 1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000010; // iC=-1534 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000010010010101; // vC= 1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b0000010010011011; // vC= 1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b0000010010110001; // vC= 1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111001; // iC=-1607 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b0000010000101111; // vC= 1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110001; // iC=-1679 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101101; // iC=-1683 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b0000010001000011; // vC= 1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100011; // iC=-1629 
vC = 14'b0000010001100000; // vC= 1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b0000010000100100; // vC= 1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b0000010001110111; // vC= 1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b0000010000110001; // vC= 1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b0000010000100001; // vC= 1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b0000010000011101; // vC= 1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b0000010000110000; // vC= 1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b0000001111010110; // vC=  982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b0000010000100001; // vC= 1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b0000010000100011; // vC= 1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111101; // iC=-1603 
vC = 14'b0000001111010111; // vC=  983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000001111100100; // vC=  996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000001110101011; // vC=  939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b0000010000101010; // vC= 1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000010000010000; // vC= 1040 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000010000100100; // vC= 1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b0000001111111010; // vC= 1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b0000001110111111; // vC=  959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b0000001111001111; // vC=  975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000010; // iC=-1662 
vC = 14'b0000001110100000; // vC=  928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b0000001110001010; // vC=  906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101010; // iC=-1750 
vC = 14'b0000001111101000; // vC= 1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000001101100110; // vC=  870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000001101011011; // vC=  859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b0000001110100111; // vC=  935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b0000001111010100; // vC=  980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000001101110111; // vC=  887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000001101010010; // vC=  850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000001110101101; // vC=  941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001100110111; // vC=  823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000001110110100; // vC=  948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b0000001110100111; // vC=  935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000001110111000; // vC=  952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b0000001100101111; // vC=  815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000001101000011; // vC=  835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000001110011101; // vC=  925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b0000001100000001; // vC=  769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000001110000111; // vC=  903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000001101010100; // vC=  852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000001011111000; // vC=  760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000001011100111; // vC=  743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b0000001101110111; // vC=  887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011000; // iC=-1704 
vC = 14'b0000001100110110; // vC=  822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001011001010; // vC=  714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000001011011010; // vC=  730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000001100011101; // vC=  797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110111; // iC=-1673 
vC = 14'b0000001100111000; // vC=  824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000001011101100; // vC=  748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000001010111111; // vC=  703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b0000001011011001; // vC=  729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101010; // iC=-1750 
vC = 14'b0000001010111110; // vC=  702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000001011011001; // vC=  729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000001011011000; // vC=  728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b0000001011001111; // vC=  719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000001011010101; // vC=  725 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000001010101000; // vC=  680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b0000001010000001; // vC=  641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000001011000011; // vC=  707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000001001011100; // vC=  604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000001010110010; // vC=  690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000001001001010; // vC=  586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000001010100100; // vC=  676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b0000001001110000; // vC=  624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000001010001100; // vC=  652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101010; // iC=-1750 
vC = 14'b0000001000111110; // vC=  574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b0000001010010011; // vC=  659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b0000001001111010; // vC=  634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001010001101; // vC=  653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000001001111010; // vC=  634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010100; // iC=-1836 
vC = 14'b0000001001100010; // vC=  610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000001000101000; // vC=  552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001110; // iC=-1842 
vC = 14'b0000000111110000; // vC=  496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000001000000011; // vC=  515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000001000101100; // vC=  556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000001001100110; // vC=  614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000001001001001; // vC=  585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000001000100000; // vC=  544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000001000010001; // vC=  529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000000110110000; // vC=  432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101001; // iC=-1815 
vC = 14'b0000001000110100; // vC=  564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001100; // iC=-1844 
vC = 14'b0000001000011001; // vC=  537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b0000000111110100; // vC=  500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b0000000110111001; // vC=  441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000001000011001; // vC=  537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000001000000011; // vC=  515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b0000000111100011; // vC=  483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000000101111111; // vC=  383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000000111110101; // vC=  501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000000111111011; // vC=  507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001110; // iC=-1842 
vC = 14'b0000000111000001; // vC=  449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b0000000110111101; // vC=  445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000101110000; // vC=  368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000101000010; // vC=  322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000000101011111; // vC=  351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b0000000110101100; // vC=  428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000000110001100; // vC=  396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000000100110010; // vC=  306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000000110100101; // vC=  421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000000101010100; // vC=  340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000000100111011; // vC=  315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000000100101110; // vC=  302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000000011111111; // vC=  255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000000101100100; // vC=  356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000000101100110; // vC=  358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b0000000101010111; // vC=  343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000000101100100; // vC=  356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000000011010110; // vC=  214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000000100111101; // vC=  317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000000010111101; // vC=  189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111010; // iC=-1798 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000000100001001; // vC=  265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001111; // iC=-1841 
vC = 14'b0000000010101111; // vC=  175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b0000000011011001; // vC=  217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000000100010001; // vC=  273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000000100011100; // vC=  284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000000100001001; // vC=  265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000000011010010; // vC=  210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000000011110100; // vC=  244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000000010001100; // vC=  140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000000100000011; // vC=  259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000000010111000; // vC=  184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000000001110110; // vC=  118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b0000000010011011; // vC=  155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b0000000001011110; // vC=   94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b0000000011000110; // vC=  198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b0000000011001001; // vC=  201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100011; // iC=-1693 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110110; // iC=-1674 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b0000000010101110; // vC=  174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b0000000010001100; // vC=  140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b0000000010001011; // vC=  139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000000000101101; // vC=   45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011101; // iC=-1699 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b0000000001100101; // vC=  101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b0000000010001011; // vC=  139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b0000000000000111; // vC=    7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b0000000000110100; // vC=   52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111111; // iC=-1665 
vC = 14'b0000000000101100; // vC=   44 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000000001001110; // vC=   78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b1111111111111100; // vC=   -4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b0000000000011000; // vC=   24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b1111111111011011; // vC=  -37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b0000000000011101; // vC=   29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b0000000000101111; // vC=   47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b1111111110101100; // vC=  -84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010010; // iC=-1646 
vC = 14'b1111111111010101; // vC=  -43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b1111111111100001; // vC=  -31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000000000000010; // vC=    2 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000001; // iC=-1663 
vC = 14'b0000000000001110; // vC=   14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110111; // iC=-1673 
vC = 14'b1111111110101001; // vC=  -87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b1111111110010101; // vC= -107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100011; // iC=-1693 
vC = 14'b0000000000000100; // vC=    4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b1111111110110101; // vC=  -75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b1111111110011010; // vC= -102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011111; // iC=-1633 
vC = 14'b1111111110100111; // vC=  -89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b1111111110000010; // vC= -126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b1111111101011111; // vC= -161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b1111111101111001; // vC= -135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b1111111111010001; // vC=  -47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010010; // iC=-1646 
vC = 14'b1111111101110001; // vC= -143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b1111111111000011; // vC=  -61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b1111111101110010; // vC= -142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b1111111110001010; // vC= -118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b1111111110000000; // vC= -128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b1111111100111001; // vC= -199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100011; // iC=-1693 
vC = 14'b1111111100111100; // vC= -196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101001; // iC=-1623 
vC = 14'b1111111100111010; // vC= -198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b1111111101111111; // vC= -129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b1111111101111111; // vC= -129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b1111111101011011; // vC= -165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b1111111011111010; // vC= -262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b1111111100100101; // vC= -219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b1111111011011000; // vC= -296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b1111111101011011; // vC= -165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010111; // iC=-1641 
vC = 14'b1111111011100011; // vC= -285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011001; // iC=-1639 
vC = 14'b1111111100110111; // vC= -201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100101; // iC=-1627 
vC = 14'b1111111011001010; // vC= -310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101101; // iC=-1683 
vC = 14'b1111111101011001; // vC= -167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000001; // iC=-1663 
vC = 14'b1111111101000000; // vC= -192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b1111111010111101; // vC= -323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b1111111100110000; // vC= -208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b1111111101000010; // vC= -190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010001; // iC=-1583 
vC = 14'b1111111010100100; // vC= -348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b1111111100000101; // vC= -251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011110; // iC=-1634 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b1111111010111100; // vC= -324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110100; // iC=-1612 
vC = 14'b1111111100100101; // vC= -219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b1111111010011011; // vC= -357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b1111111011111010; // vC= -262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b1111111010010101; // vC= -363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b1111111011101111; // vC= -273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b1111111010111001; // vC= -327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110111; // iC=-1673 
vC = 14'b1111111011000011; // vC= -317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b1111111011111010; // vC= -262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b1111111010000001; // vC= -383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011111; // iC=-1633 
vC = 14'b1111111010110000; // vC= -336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111111; // iC=-1665 
vC = 14'b1111111011000000; // vC= -320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b1111111001010001; // vC= -431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b1111111001010000; // vC= -432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b1111111001111001; // vC= -391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010100; // iC=-1580 
vC = 14'b1111111010111011; // vC= -325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b1111111010111110; // vC= -322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b1111111001110010; // vC= -398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b1111111001100001; // vC= -415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b1111111001110100; // vC= -396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b1111111000101110; // vC= -466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b1111111000111101; // vC= -451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b1111111000011000; // vC= -488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001110; // iC=-1586 
vC = 14'b1111110111110111; // vC= -521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b1111111001101000; // vC= -408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b1111110111110110; // vC= -522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b1111110111101000; // vC= -536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010111; // iC=-1513 
vC = 14'b1111110111111010; // vC= -518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101100; // iC=-1556 
vC = 14'b1111110111111000; // vC= -520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100111; // iC=-1497 
vC = 14'b1111111000000011; // vC= -509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b1111110111101000; // vC= -536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110101; // iC=-1611 
vC = 14'b1111111001000111; // vC= -441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b1111110111000010; // vC= -574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101110; // iC=-1618 
vC = 14'b1111110110111110; // vC= -578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b1111111000010110; // vC= -490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b1111111000110110; // vC= -458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100110; // iC=-1562 
vC = 14'b1111110110100001; // vC= -607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b1111110111100011; // vC= -541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110001; // iC=-1487 
vC = 14'b1111110110011000; // vC= -616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101011; // iC=-1493 
vC = 14'b1111110111110100; // vC= -524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b1111110111010101; // vC= -555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b1111110111010100; // vC= -556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101101; // iC=-1491 
vC = 14'b1111110110000000; // vC= -640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b1111110111011110; // vC= -546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b1111110110001101; // vC= -627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000011; // iC=-1533 
vC = 14'b1111110111010111; // vC= -553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b1111110110001100; // vC= -628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b1111110110010001; // vC= -623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001110; // iC=-1458 
vC = 14'b1111110111010111; // vC= -553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100100; // iC=-1436 
vC = 14'b1111110110111000; // vC= -584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b1111110111000000; // vC= -576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b1111110110111011; // vC= -581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001010; // iC=-1526 
vC = 14'b1111110111010001; // vC= -559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100011; // iC=-1501 
vC = 14'b1111110110010100; // vC= -620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b1111110110101111; // vC= -593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001101; // iC=-1459 
vC = 14'b1111110111001010; // vC= -566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b1111110100100111; // vC= -729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001010; // iC=-1398 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001001; // iC=-1399 
vC = 14'b1111110101000000; // vC= -704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b1111110110111001; // vC= -583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001111; // iC=-1457 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100010; // iC=-1502 
vC = 14'b1111110110000011; // vC= -637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b1111110110100000; // vC= -608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b1111110100110010; // vC= -718 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011110; // iC=-1378 
vC = 14'b1111110100111101; // vC= -707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111110100000101; // vC= -763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001110; // iC=-1458 
vC = 14'b1111110100010100; // vC= -748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b1111110100001001; // vC= -759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100010; // iC=-1374 
vC = 14'b1111110011110000; // vC= -784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111010; // iC=-1478 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b1111110100000110; // vC= -762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110010; // iC=-1422 
vC = 14'b1111110100000110; // vC= -762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001101; // iC=-1395 
vC = 14'b1111110100110110; // vC= -714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111110011111100; // vC= -772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000100; // iC=-1404 
vC = 14'b1111110101001011; // vC= -693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111110011110011; // vC= -781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011000; // iC=-1384 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111001; // iC=-1351 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111101; // iC=-1347 
vC = 14'b1111110100011111; // vC= -737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b1111110100011110; // vC= -738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011101; // iC=-1443 
vC = 14'b1111110100101111; // vC= -721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110010; // iC=-1422 
vC = 14'b1111110100111110; // vC= -706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b1111110100001100; // vC= -756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110110; // iC=-1418 
vC = 14'b1111110011011101; // vC= -803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100101; // iC=-1435 
vC = 14'b1111110100000100; // vC= -764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111100; // iC=-1284 
vC = 14'b1111110010011101; // vC= -867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100100; // iC=-1436 
vC = 14'b1111110100000101; // vC= -763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011011; // iC=-1381 
vC = 14'b1111110011111000; // vC= -776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110000; // iC=-1296 
vC = 14'b1111110011101000; // vC= -792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111101; // iC=-1411 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101100; // iC=-1300 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100010; // iC=-1310 
vC = 14'b1111110010010101; // vC= -875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111000; // iC=-1352 
vC = 14'b1111110001110111; // vC= -905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111110010001111; // vC= -881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000010; // iC=-1342 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100001; // iC=-1247 
vC = 14'b1111110001010100; // vC= -940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101010; // iC=-1302 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110111; // iC=-1289 
vC = 14'b1111110010111010; // vC= -838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100011; // iC=-1373 
vC = 14'b1111110001111010; // vC= -902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100110; // iC=-1370 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100111; // iC=-1369 
vC = 14'b1111110010010110; // vC= -874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000001; // iC=-1279 
vC = 14'b1111110001100000; // vC= -928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110011; // iC=-1357 
vC = 14'b1111110000111100; // vC= -964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110010; // iC=-1294 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001011; // iC=-1269 
vC = 14'b1111110010100011; // vC= -861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000001; // iC=-1279 
vC = 14'b1111110011000000; // vC= -832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010101; // iC=-1195 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111001; // iC=-1223 
vC = 14'b1111110010100111; // vC= -857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001000; // iC=-1208 
vC = 14'b1111110000011011; // vC= -997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100000; // iC=-1184 
vC = 14'b1111110001110101; // vC= -907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110000; // iC=-1296 
vC = 14'b1111110001110011; // vC= -909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101100; // iC=-1300 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111100; // iC=-1284 
vC = 14'b1111110001001101; // vC= -947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b1111110001001000; // vC= -952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b1111110001000011; // vC= -957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101000; // iC=-1176 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110000; // iC=-1296 
vC = 14'b1111110001010100; // vC= -940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b1111101111110100; // vC=-1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110001; // iC=-1231 
vC = 14'b1111101111110111; // vC=-1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111101; // iC=-1283 
vC = 14'b1111110000001000; // vC=-1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000111; // iC=-1209 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001010; // iC=-1142 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110111; // iC=-1161 
vC = 14'b1111110000101000; // vC= -984 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011011; // iC=-1189 
vC = 14'b1111110000000010; // vC=-1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010100; // iC=-1132 
vC = 14'b1111101111011101; // vC=-1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010100; // iC=-1132 
vC = 14'b1111110000000001; // vC=-1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010000; // iC=-1264 
vC = 14'b1111101111111010; // vC=-1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111001; // iC=-1223 
vC = 14'b1111110000011010; // vC= -998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010100; // iC=-1260 
vC = 14'b1111110000010111; // vC=-1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b1111110001001100; // vC= -948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b1111110000111001; // vC= -967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111111; // iC=-1153 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010001; // iC=-1199 
vC = 14'b1111101111111001; // vC=-1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001101; // iC=-1139 
vC = 14'b1111101111001100; // vC=-1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010001; // iC=-1071 
vC = 14'b1111101111000010; // vC=-1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010111; // iC=-1129 
vC = 14'b1111101111000101; // vC=-1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110100; // iC=-1164 
vC = 14'b1111101111101100; // vC=-1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010001; // iC=-1135 
vC = 14'b1111101111011101; // vC=-1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011011; // iC=-1189 
vC = 14'b1111101111001010; // vC=-1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000010; // iC=-1150 
vC = 14'b1111101110101000; // vC=-1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101001; // iC=-1175 
vC = 14'b1111101111010001; // vC=-1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001100; // iC=-1140 
vC = 14'b1111101111001111; // vC=-1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101100; // iC=-1172 
vC = 14'b1111110000000011; // vC=-1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110010; // iC=-1038 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000011; // iC=-1085 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010011; // iC=-1133 
vC = 14'b1111101110000111; // vC=-1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101100; // iC=-1108 
vC = 14'b1111101111011000; // vC=-1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000010; // iC=-1086 
vC = 14'b1111101101101100; // vC=-1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000111; // iC=-1017 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001001; // iC=-1079 
vC = 14'b1111101111010110; // vC=-1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010100; // iC=-1004 
vC = 14'b1111101111100111; // vC=-1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011101; // iC= -995 
vC = 14'b1111101111101101; // vC=-1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100010; // iC= -990 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011101; // iC= -995 
vC = 14'b1111101101011111; // vC=-1185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100010; // iC=-1054 
vC = 14'b1111101111000010; // vC=-1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000000; // iC=-1024 
vC = 14'b1111101110101001; // vC=-1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011010; // iC= -998 
vC = 14'b1111101101101111; // vC=-1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111100; // iC= -964 
vC = 14'b1111101101110111; // vC=-1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010101; // iC=-1067 
vC = 14'b1111101101011010; // vC=-1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010100; // iC=-1004 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111101; // iC=-1091 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101100; // iC=-1044 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111011; // iC=-1093 
vC = 14'b1111101110001010; // vC=-1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011110; // iC=-1058 
vC = 14'b1111101110110001; // vC=-1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010010; // iC= -942 
vC = 14'b1111101101101110; // vC=-1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001100; // iC= -948 
vC = 14'b1111101110100001; // vC=-1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000011; // iC=-1021 
vC = 14'b1111101100110111; // vC=-1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101010; // iC= -918 
vC = 14'b1111101101101011; // vC=-1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101101; // iC=-1043 
vC = 14'b1111101100100100; // vC=-1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010001; // iC=-1007 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100110; // iC= -922 
vC = 14'b1111101101001101; // vC=-1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110111; // iC= -969 
vC = 14'b1111101100100111; // vC=-1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101011; // iC=-1045 
vC = 14'b1111101100011001; // vC=-1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100101; // iC= -923 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111001; // iC=-1031 
vC = 14'b1111101110000110; // vC=-1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001111; // iC=-1009 
vC = 14'b1111101100010011; // vC=-1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010010; // iC=-1006 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001001; // iC= -951 
vC = 14'b1111101101110100; // vC=-1164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010110; // iC= -874 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111001; // iC= -903 
vC = 14'b1111101101100111; // vC=-1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010111; // iC= -937 
vC = 14'b1111101100111011; // vC=-1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001101; // iC= -947 
vC = 14'b1111101101001000; // vC=-1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001000; // iC= -888 
vC = 14'b1111101100011000; // vC=-1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010100; // iC= -876 
vC = 14'b1111101101000110; // vC=-1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b1111101101101100; // vC=-1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000100; // iC= -956 
vC = 14'b1111101011111111; // vC=-1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001001; // iC= -823 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010011; // iC= -877 
vC = 14'b1111101100001010; // vC=-1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100011; // iC= -861 
vC = 14'b1111101011111100; // vC=-1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000010; // iC= -894 
vC = 14'b1111101100011011; // vC=-1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011011; // iC= -869 
vC = 14'b1111101101010010; // vC=-1198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111111; // iC= -897 
vC = 14'b1111101011100100; // vC=-1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001000; // iC= -824 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010110; // iC= -810 
vC = 14'b1111101011111010; // vC=-1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011111; // iC= -865 
vC = 14'b1111101011111011; // vC=-1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101100; // iC= -852 
vC = 14'b1111101100001100; // vC=-1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101011; // iC= -853 
vC = 14'b1111101100101000; // vC=-1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111000; // iC= -776 
vC = 14'b1111101101001000; // vC=-1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111011; // iC= -901 
vC = 14'b1111101011010110; // vC=-1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110101; // iC= -907 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001000; // iC= -888 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110101; // iC= -779 
vC = 14'b1111101100101000; // vC=-1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010110; // iC= -746 
vC = 14'b1111101101000110; // vC=-1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001011; // iC= -757 
vC = 14'b1111101101001011; // vC=-1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010000; // iC= -816 
vC = 14'b1111101011110011; // vC=-1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010011; // iC= -877 
vC = 14'b1111101100011111; // vC=-1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100001; // iC= -799 
vC = 14'b1111101011101001; // vC=-1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110101; // iC= -843 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101001; // iC= -855 
vC = 14'b1111101100111011; // vC=-1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011001; // iC= -807 
vC = 14'b1111101010110100; // vC=-1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011100; // iC= -740 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111001; // iC= -711 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101001; // iC= -791 
vC = 14'b1111101011000011; // vC=-1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000100; // iC= -764 
vC = 14'b1111101011100010; // vC=-1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111100; // iC= -708 
vC = 14'b1111101100001001; // vC=-1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010011; // iC= -749 
vC = 14'b1111101011111110; // vC=-1282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000101; // iC= -699 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001111; // iC= -817 
vC = 14'b1111101010110011; // vC=-1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101101; // iC= -787 
vC = 14'b1111101010110100; // vC=-1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100000; // iC= -672 
vC = 14'b1111101100001000; // vC=-1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100110; // iC= -794 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100100; // iC= -668 
vC = 14'b1111101010110111; // vC=-1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110111; // iC= -777 
vC = 14'b1111101011110100; // vC=-1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100010; // iC= -734 
vC = 14'b1111101001111100; // vC=-1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110110; // iC= -650 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001100; // iC= -756 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001001; // iC= -695 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011001; // iC= -679 
vC = 14'b1111101010011000; // vC=-1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010001; // iC= -623 
vC = 14'b1111101001111110; // vC=-1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110000; // iC= -720 
vC = 14'b1111101011011001; // vC=-1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101110; // iC= -594 
vC = 14'b1111101011010001; // vC=-1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111101; // iC= -643 
vC = 14'b1111101010101110; // vC=-1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100001; // iC= -671 
vC = 14'b1111101011010000; // vC=-1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011010; // iC= -678 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011011; // iC= -613 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011111; // iC= -673 
vC = 14'b1111101011100111; // vC=-1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001001; // iC= -631 
vC = 14'b1111101010001011; // vC=-1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001101; // iC= -563 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000001; // iC= -575 
vC = 14'b1111101010000010; // vC=-1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111001; // iC= -583 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000011; // iC= -573 
vC = 14'b1111101010011101; // vC=-1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111000; // iC= -584 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110110; // iC= -650 
vC = 14'b1111101001101110; // vC=-1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011010; // iC= -550 
vC = 14'b1111101001110000; // vC=-1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010000; // iC= -560 
vC = 14'b1111101001011110; // vC=-1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111110; // iC= -578 
vC = 14'b1111101010010010; // vC=-1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101100; // iC= -596 
vC = 14'b1111101001110011; // vC=-1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111101; // iC= -515 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001110; // iC= -498 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110100; // iC= -524 
vC = 14'b1111101010011010; // vC=-1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001111; // iC= -561 
vC = 14'b1111101011011011; // vC=-1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100010; // iC= -606 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110111; // iC= -585 
vC = 14'b1111101000110111; // vC=-1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011000; // iC= -552 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110101; // iC= -459 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000111; // iC= -505 
vC = 14'b1111101010011100; // vC=-1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111011; // iC= -517 
vC = 14'b1111101000110101; // vC=-1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101001; // iC= -535 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000111; // iC= -569 
vC = 14'b1111101001101110; // vC=-1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111111; // iC= -513 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100100; // iC= -540 
vC = 14'b1111101000101111; // vC=-1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001101; // iC= -435 
vC = 14'b1111101010100001; // vC=-1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101100; // iC= -468 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100000; // iC= -416 
vC = 14'b1111101001111110; // vC=-1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100111; // iC= -473 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011001; // iC= -551 
vC = 14'b1111101010101110; // vC=-1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000010; // iC= -510 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010100; // iC= -492 
vC = 14'b1111101001111110; // vC=-1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111101; // iC= -451 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001110; // iC= -498 
vC = 14'b1111101001101101; // vC=-1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011000; // iC= -488 
vC = 14'b1111101000111001; // vC=-1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011100; // iC= -420 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100010; // iC= -350 
vC = 14'b1111101000110100; // vC=-1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110000; // iC= -464 
vC = 14'b1111101001100001; // vC=-1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000011; // iC= -445 
vC = 14'b1111101000011100; // vC=-1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110110; // iC= -458 
vC = 14'b1111101010001000; // vC=-1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001011; // iC= -309 
vC = 14'b1111101001001000; // vC=-1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100011; // iC= -349 
vC = 14'b1111101000110101; // vC=-1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010001; // iC= -303 
vC = 14'b1111101000001100; // vC=-1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100111; // iC= -345 
vC = 14'b1111101010010000; // vC=-1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011001; // iC= -295 
vC = 14'b1111101010010110; // vC=-1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000100; // iC= -252 
vC = 14'b1111101010001001; // vC=-1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001010; // iC= -374 
vC = 14'b1111101001110100; // vC=-1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011110; // iC= -226 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110001; // iC= -335 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100001; // iC= -223 
vC = 14'b1111101000100010; // vC=-1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101001; // iC= -279 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011001; // iC= -295 
vC = 14'b1111101010011100; // vC=-1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011010; // iC= -166 
vC = 14'b1111101001110001; // vC=-1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101111; // iC= -273 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100011; // iC= -285 
vC = 14'b1111101001011000; // vC=-1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110110; // iC= -266 
vC = 14'b1111101001110101; // vC=-1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101110; // iC= -146 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000111; // iC= -121 
vC = 14'b1111101000101100; // vC=-1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101101; // iC=  -83 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111000; // iC= -200 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010000; // iC= -176 
vC = 14'b1111101000100010; // vC=-1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001000; // iC=  -56 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110110; // iC=  -10 
vC = 14'b1111101000010101; // vC=-1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010010; // iC=  -46 
vC = 14'b1111101000110110; // vC=-1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110111; // iC=  -73 
vC = 14'b1111101000010011; // vC=-1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100001; // iC=  -31 
vC = 14'b1111101010001011; // vC=-1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111011; // iC=  -69 
vC = 14'b1111101001010001; // vC=-1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000001; // iC=   65 
vC = 14'b1111101000001000; // vC=-1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101110; // iC=   46 
vC = 14'b1111101010010111; // vC=-1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101100; // iC=   44 
vC = 14'b1111101001010001; // vC=-1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010000; // iC=   80 
vC = 14'b1111101001100101; // vC=-1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101001; // iC=  105 
vC = 14'b1111101000111100; // vC=-1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100000; // iC=   32 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111000; // iC=  120 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011011; // iC=   91 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110010; // iC=  114 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011010; // iC=  218 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101111; // iC=  239 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110000; // iC=  176 
vC = 14'b1111101000111011; // vC=-1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100010; // iC=  290 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010010; // iC=  338 
vC = 14'b1111101000101111; // vC=-1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111001; // iC=  313 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000100; // iC=  388 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100100; // iC=  292 
vC = 14'b1111101000011111; // vC=-1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111110; // iC=  382 
vC = 14'b1111101001100001; // vC=-1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101111; // iC=  431 
vC = 14'b1111101000011010; // vC=-1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110111; // iC=  375 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101110; // iC=  366 
vC = 14'b1111101001111011; // vC=-1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001010; // iC=  458 
vC = 14'b1111101000110101; // vC=-1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001111; // iC=  527 
vC = 14'b1111101001010001; // vC=-1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000111; // iC=  455 
vC = 14'b1111101010010001; // vC=-1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100101; // iC=  613 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111111; // iC=  575 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001000; // iC=  520 
vC = 14'b1111101000110000; // vC=-1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000011; // iC=  579 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100011; // iC=  547 
vC = 14'b1111101010001111; // vC=-1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001011; // iC=  715 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110110; // iC=  630 
vC = 14'b1111101000111011; // vC=-1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001010; // iC=  714 
vC = 14'b1111101000100100; // vC=-1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011010; // iC=  666 
vC = 14'b1111101001110001; // vC=-1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100011; // iC=  803 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000001; // iC=  769 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b1111101000101111; // vC=-1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100110; // iC=  806 
vC = 14'b1111101011000001; // vC=-1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011000; // iC=  792 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010001; // iC=  849 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001101; // iC=  845 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000000; // iC=  896 
vC = 14'b1111101010111110; // vC=-1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110000; // iC=  944 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110101; // iC= 1013 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101001; // iC= 1001 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100100; // iC= 1060 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101011; // iC=  939 
vC = 14'b1111101011010010; // vC=-1326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101011; // iC= 1003 
vC = 14'b1111101010010100; // vC=-1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010100; // iC= 1108 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101010; // iC= 1002 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110001; // iC= 1073 
vC = 14'b1111101010001110; // vC=-1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000001; // iC= 1153 
vC = 14'b1111101011100111; // vC=-1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000001; // iC= 1089 
vC = 14'b1111101011101001; // vC=-1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000000; // iC= 1216 
vC = 14'b1111101011110001; // vC=-1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001100; // iC= 1164 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010100; // iC= 1172 
vC = 14'b1111101010001001; // vC=-1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011000; // iC= 1176 
vC = 14'b1111101100010100; // vC=-1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000010; // iC= 1282 
vC = 14'b1111101100000100; // vC=-1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101001; // iC= 1257 
vC = 14'b1111101010001000; // vC=-1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010111; // iC= 1239 
vC = 14'b1111101011111001; // vC=-1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110100; // iC= 1268 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111110; // iC= 1342 
vC = 14'b1111101011110100; // vC=-1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000000; // iC= 1280 
vC = 14'b1111101100010111; // vC=-1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000001; // iC= 1409 
vC = 14'b1111101010101010; // vC=-1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101011; // iC= 1451 
vC = 14'b1111101100101011; // vC=-1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111010; // iC= 1338 
vC = 14'b1111101100110111; // vC=-1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001101; // iC= 1421 
vC = 14'b1111101010111010; // vC=-1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110011; // iC= 1395 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100000; // iC= 1376 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101001; // iC= 1449 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001111; // iC= 1423 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101011; // iC= 1451 
vC = 14'b1111101011111111; // vC=-1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101110; // iC= 1582 
vC = 14'b1111101101010001; // vC=-1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111111; // iC= 1471 
vC = 14'b1111101100001001; // vC=-1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010001; // iC= 1617 
vC = 14'b1111101011110011; // vC=-1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b1111101101101001; // vC=-1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110100; // iC= 1652 
vC = 14'b1111101101001011; // vC=-1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100001; // iC= 1633 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011010; // iC= 1626 
vC = 14'b1111101100101001; // vC=-1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100100; // iC= 1572 
vC = 14'b1111101101000001; // vC=-1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011110; // iC= 1630 
vC = 14'b1111101110100001; // vC=-1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011110; // iC= 1630 
vC = 14'b1111101110011011; // vC=-1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110001; // iC= 1713 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b1111101100111110; // vC=-1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b1111101110101100; // vC=-1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110000; // iC= 1648 
vC = 14'b1111101101110100; // vC=-1164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b1111101110101010; // vC=-1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000110; // iC= 1734 
vC = 14'b1111101101111000; // vC=-1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110110; // iC= 1654 
vC = 14'b1111101111000101; // vC=-1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b1111101101101000; // vC=-1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b1111101110111111; // vC=-1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b1111101110101100; // vC=-1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b1111101110011001; // vC=-1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010111; // iC= 1751 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b1111101111101000; // vC=-1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110101; // iC= 1845 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b1111101110101111; // vC=-1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b1111101101111100; // vC=-1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111101110100100; // vC=-1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b1111101110111111; // vC=-1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b1111101110010110; // vC=-1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b1111101111001101; // vC=-1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110000; // iC= 1840 
vC = 14'b1111110000000010; // vC=-1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111101111011000; // vC=-1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000111; // iC= 1863 
vC = 14'b1111101111001111; // vC=-1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111110000001100; // vC=-1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111110001001010; // vC= -950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b1111110000001100; // vC=-1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b1111101111111111; // vC=-1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b1111110000001110; // vC=-1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b1111110001100000; // vC= -928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111110000011101; // vC= -995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001101; // iC= 1869 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b1111110001100011; // vC= -925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b1111110000110010; // vC= -974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111101111111100; // vC=-1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b1111110000011101; // vC= -995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101011; // iC= 1835 
vC = 14'b1111110001111001; // vC= -903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101100; // iC= 1964 
vC = 14'b1111110001110100; // vC= -908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111110001100001; // vC= -927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110001111111; // vC= -897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b1111110001111011; // vC= -901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b1111110010010011; // vC= -877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110010000010; // vC= -894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111110011000011; // vC= -829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111110001101000; // vC= -920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111110011110100; // vC= -780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001010; // iC= 1866 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b1111110010000000; // vC= -896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111101; // iC= 1853 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111110011110011; // vC= -781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b1111110011111110; // vC= -770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011101; // iC= 2013 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001001; // iC= 1865 
vC = 14'b1111110011100110; // vC= -794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110101001011; // vC= -693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110011010100; // vC= -812 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b1111110100011000; // vC= -744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110101100010; // vC= -670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111110100101110; // vC= -722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111110011110001; // vC= -783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b1111110100011111; // vC= -737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b1111110100111011; // vC= -709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111110110000111; // vC= -633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111110100011000; // vC= -744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b1111110110100001; // vC= -607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101011; // iC= 2027 
vC = 14'b1111110101000000; // vC= -704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010100; // iC= 2004 
vC = 14'b1111110101111000; // vC= -648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111110110100010; // vC= -606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111110110101110; // vC= -594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b1111110101010011; // vC= -685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b1111110101110111; // vC= -649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111110110111001; // vC= -583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b1111110111000111; // vC= -569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011110; // iC= 1886 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111110111001000; // vC= -568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011101; // iC= 2013 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b1111110111101100; // vC= -532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b1111110111110100; // vC= -524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b1111110101111111; // vC= -641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111111000000111; // vC= -505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b1111111000010111; // vC= -489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111110111101100; // vC= -532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111110111000001; // vC= -575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b1111110110011110; // vC= -610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b1111111000010010; // vC= -494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111110110110011; // vC= -589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111110111000000; // vC= -576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b1111111001001101; // vC= -435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b1111111000000001; // vC= -511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111111000000111; // vC= -505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111110111110010; // vC= -526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000100; // iC= 1924 
vC = 14'b1111110111111100; // vC= -516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111110111111011; // vC= -517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111111001111010; // vC= -390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b1111111010000000; // vC= -384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111110111111110; // vC= -514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111111000101011; // vC= -469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b1111111000000100; // vC= -508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b1111111000000111; // vC= -505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111111010011010; // vC= -358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111111001101001; // vC= -407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111111000100011; // vC= -477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111110; // iC= 1982 
vC = 14'b1111111001000101; // vC= -443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b1111111010001000; // vC= -376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111111011000110; // vC= -314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b1111111010100100; // vC= -348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111111010100110; // vC= -346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110010; // iC= 2034 
vC = 14'b1111111010011011; // vC= -357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111111001101110; // vC= -402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001100; // iC= 2060 
vC = 14'b1111111010100111; // vC= -345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b1111111011101011; // vC= -277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001101; // iC= 2061 
vC = 14'b1111111001111010; // vC= -390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111111001110011; // vC= -397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111111011000001; // vC= -319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b1111111010111111; // vC= -321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111111011110100; // vC= -268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111111010000001; // vC= -383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b1111111010101100; // vC= -340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111110; // iC= 1982 
vC = 14'b1111111100101101; // vC= -211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111111011111101; // vC= -259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b1111111010100000; // vC= -352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111111100011101; // vC= -227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b1111111100101011; // vC= -213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b1111111011010001; // vC= -303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111111101010010; // vC= -174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b1111111100000001; // vC= -255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111111011111111; // vC= -257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111111011111011; // vC= -261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111100001111; // vC= -241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111111101010101; // vC= -171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111101100100; // vC= -156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b1111111011111111; // vC= -257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101011; // iC= 2027 
vC = 14'b1111111100111100; // vC= -196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111111101101011; // vC= -149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100010; // iC= 2018 
vC = 14'b1111111110000001; // vC= -127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b1111111110011111; // vC=  -97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000111; // iC= 1991 
vC = 14'b1111111101001111; // vC= -177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111111100111110; // vC= -194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b1111111110110011; // vC=  -77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000000; // iC= 1984 
vC = 14'b1111111101100011; // vC= -157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011011; // iC= 2011 
vC = 14'b1111111100111100; // vC= -196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101010; // iC= 1898 
vC = 14'b1111111111011010; // vC=  -38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b1111111110110110; // vC=  -74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111111111001110; // vC=  -50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100011; // iC= 2019 
vC = 14'b1111111111001101; // vC=  -51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b1111111111000011; // vC=  -61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111111101100110; // vC= -154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111111111001010; // vC=  -54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b0000000000001000; // vC=    8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111111110101011; // vC=  -85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111111110101111; // vC=  -81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111111111000111; // vC=  -57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111111110111111; // vC=  -65 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111111111000100; // vC=  -60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111111010010; // vC=  -46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b1111111111000101; // vC=  -59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b1111111111111000; // vC=   -8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011001; // iC= 1881 
vC = 14'b0000000000111000; // vC=   56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011100; // iC= 1948 
vC = 14'b1111111111101001; // vC=  -23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111111111001000; // vC=  -56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001111; // iC= 1871 
vC = 14'b0000000000000110; // vC=    6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b0000000001110001; // vC=  113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b1111111111111111; // vC=   -1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b0000000001011101; // vC=   93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111111111101011; // vC=  -21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b0000000000010010; // vC=   18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b0000000000010100; // vC=   20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010100; // iC= 2004 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b0000000001000101; // vC=   69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110010; // iC= 1906 
vC = 14'b0000000001110101; // vC=  117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011100; // iC= 1948 
vC = 14'b0000000001101011; // vC=  107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b0000000010111000; // vC=  184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b0000000001110010; // vC=  114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b0000000010010110; // vC=  150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b0000000010011101; // vC=  157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b0000000010001101; // vC=  141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b0000000010111101; // vC=  189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b0000000010001001; // vC=  137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b0000000001010111; // vC=   87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b0000000010001010; // vC=  138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b0000000010000100; // vC=  132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b0000000010000110; // vC=  134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b0000000011000010; // vC=  194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111101; // iC= 1853 
vC = 14'b0000000010010010; // vC=  146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b0000000010011001; // vC=  153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b0000000011111110; // vC=  254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b0000000011100001; // vC=  225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b0000000100011000; // vC=  280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001000; // iC= 1864 
vC = 14'b0000000100010101; // vC=  277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b0000000010110010; // vC=  178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b0000000100100010; // vC=  290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b0000000100001001; // vC=  265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b0000000101001010; // vC=  330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b0000000100100000; // vC=  288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b0000000100010011; // vC=  275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b0000000011101110; // vC=  238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b0000000011101110; // vC=  238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b0000000011101101; // vC=  237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b0000000101001101; // vC=  333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001001; // iC= 1865 
vC = 14'b0000000101100010; // vC=  354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b0000000101110010; // vC=  370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b0000000100100001; // vC=  289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b0000000100010111; // vC=  279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110001; // iC= 1841 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001010; // iC= 1866 
vC = 14'b0000000100011000; // vC=  280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b0000000100111101; // vC=  317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010011; // iC= 1811 
vC = 14'b0000000101111001; // vC=  377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b0000000110010111; // vC=  407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b0000000101010010; // vC=  338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011100; // iC= 1820 
vC = 14'b0000000111000101; // vC=  453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000000101000101; // vC=  325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b0000000101111101; // vC=  381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000000110111011; // vC=  443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b0000000110111011; // vC=  443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b0000000110101100; // vC=  428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b0000000101111100; // vC=  380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011011; // iC= 1755 
vC = 14'b0000000111101111; // vC=  495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b0000000101101111; // vC=  367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b0000000101110000; // vC=  368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b0000000110011010; // vC=  410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110001; // iC= 1777 
vC = 14'b0000000101111110; // vC=  382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b0000000110101000; // vC=  424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111001; // iC= 1785 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b0000001000101100; // vC=  556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000001000110110; // vC=  566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010010; // iC= 1874 
vC = 14'b0000000111001110; // vC=  462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b0000000111001100; // vC=  460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b0000001000000010; // vC=  514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111000; // iC= 1720 
vC = 14'b0000000111101011; // vC=  491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b0000000111101101; // vC=  493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101100; // iC= 1772 
vC = 14'b0000001001101001; // vC=  617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b0000001001101011; // vC=  619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b0000001001110011; // vC=  627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b0000001000011010; // vC=  538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b0000001001000001; // vC=  577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101011; // iC= 1707 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101011; // iC= 1707 
vC = 14'b0000001001100010; // vC=  610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010100; // iC= 1748 
vC = 14'b0000001001010110; // vC=  598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000111; // iC= 1799 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b0000001001010000; // vC=  592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101111; // iC= 1711 
vC = 14'b0000001001100011; // vC=  611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000001000101000; // vC=  552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000011; // iC= 1795 
vC = 14'b0000001010011000; // vC=  664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b0000001000110000; // vC=  560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110001; // iC= 1777 
vC = 14'b0000001000100111; // vC=  551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b0000001011000011; // vC=  707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001110; // iC= 1742 
vC = 14'b0000001001101100; // vC=  620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000010; // iC= 1794 
vC = 14'b0000001011010111; // vC=  727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101001; // iC= 1705 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000001011001010; // vC=  714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b0000001010110011; // vC=  691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000001010000110; // vC=  646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b0000001001011001; // vC=  601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b0000001010001010; // vC=  650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b0000001001111010; // vC=  634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100001; // iC= 1633 
vC = 14'b0000001010010011; // vC=  659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111011; // iC= 1659 
vC = 14'b0000001001111101; // vC=  637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b0000001011110011; // vC=  755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000001010000011; // vC=  643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b0000001100100111; // vC=  807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001110; // iC= 1678 
vC = 14'b0000001100010101; // vC=  789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b0000001010011010; // vC=  666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001110; // iC= 1678 
vC = 14'b0000001100011101; // vC=  797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b0000001011101010; // vC=  746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010101; // iC= 1749 
vC = 14'b0000001100111111; // vC=  831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000001100010100; // vC=  788 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101111; // iC= 1711 
vC = 14'b0000001011100011; // vC=  739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101000; // iC= 1640 
vC = 14'b0000001100100010; // vC=  802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b0000001011100001; // vC=  737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001001; // iC= 1737 
vC = 14'b0000001100101001; // vC=  809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b0000001011111110; // vC=  766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101011; // iC= 1579 
vC = 14'b0000001101100100; // vC=  868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b0000001101001101; // vC=  845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101111; // iC= 1583 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000111; // iC= 1671 
vC = 14'b0000001101010011; // vC=  851 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b0000001011101101; // vC=  749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100110; // iC= 1574 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110001; // iC= 1649 
vC = 14'b0000001100011011; // vC=  795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000101; // iC= 1669 
vC = 14'b0000001100111110; // vC=  830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111001; // iC= 1593 
vC = 14'b0000001101101100; // vC=  876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011111; // iC= 1695 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000101; // iC= 1541 
vC = 14'b0000001110000111; // vC=  903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011001; // iC= 1625 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110101; // iC= 1525 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b0000001110000111; // vC=  903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b0000001101000111; // vC=  839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b0000001110000110; // vC=  902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101101; // iC= 1645 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110101; // iC= 1589 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110100; // iC= 1524 
vC = 14'b0000001110100110; // vC=  934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001001; // iC= 1609 
vC = 14'b0000001101101000; // vC=  872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101111; // iC= 1519 
vC = 14'b0000001110011101; // vC=  925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010010; // iC= 1554 
vC = 14'b0000001110101111; // vC=  943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110111; // iC= 1527 
vC = 14'b0000001101101011; // vC=  875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100111; // iC= 1511 
vC = 14'b0000001101101100; // vC=  876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001101; // iC= 1549 
vC = 14'b0000001111010001; // vC=  977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111111; // iC= 1599 
vC = 14'b0000001111000001; // vC=  961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b0000001101110101; // vC=  885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111011; // iC= 1595 
vC = 14'b0000001111100101; // vC=  997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010010; // iC= 1490 
vC = 14'b0000001110011101; // vC=  925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101010; // iC= 1578 
vC = 14'b0000001111000101; // vC=  965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010111; // iC= 1559 
vC = 14'b0000001101110011; // vC=  883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000101; // iC= 1477 
vC = 14'b0000001110010101; // vC=  917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101000; // iC= 1576 
vC = 14'b0000001111010001; // vC=  977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011010; // iC= 1498 
vC = 14'b0000001110111111; // vC=  959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001011; // iC= 1547 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b0000001111111100; // vC= 1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101001; // iC= 1449 
vC = 14'b0000001110011001; // vC=  921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011101; // iC= 1501 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000010; // iC= 1474 
vC = 14'b0000010000110000; // vC= 1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100101; // iC= 1509 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001000; // iC= 1416 
vC = 14'b0000010000111100; // vC= 1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001010; // iC= 1546 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001101; // iC= 1549 
vC = 14'b0000001111110111; // vC= 1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001011; // iC= 1419 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b0000001111011100; // vC=  988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001100; // iC= 1484 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000111; // iC= 1543 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110000; // iC= 1392 
vC = 14'b0000010000111001; // vC= 1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011000; // iC= 1496 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010111; // iC= 1431 
vC = 14'b0000010000111011; // vC= 1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101101; // iC= 1453 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110111; // iC= 1463 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110011; // iC= 1523 
vC = 14'b0000001111100000; // vC=  992 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110000; // iC= 1392 
vC = 14'b0000001111101000; // vC= 1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011100; // iC= 1372 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101000; // iC= 1384 
vC = 14'b0000010000010101; // vC= 1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001000; // iC= 1480 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010001; // iC= 1489 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111111; // iC= 1407 
vC = 14'b0000001111111000; // vC= 1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111011; // iC= 1339 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001011; // iC= 1355 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111010; // iC= 1466 
vC = 14'b0000010000001010; // vC= 1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101000; // iC= 1320 
vC = 14'b0000010001000101; // vC= 1093 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011001; // iC= 1433 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110100; // iC= 1396 
vC = 14'b0000010010010111; // vC= 1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010100; // iC= 1428 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011000; // iC= 1432 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010011; // iC= 1427 
vC = 14'b0000010001110011; // vC= 1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010001; // iC= 1297 
vC = 14'b0000010010000001; // vC= 1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101110; // iC= 1326 
vC = 14'b0000010010001001; // vC= 1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011101; // iC= 1437 
vC = 14'b0000010010110101; // vC= 1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000011; // iC= 1283 
vC = 14'b0000010001110000; // vC= 1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000101; // iC= 1285 
vC = 14'b0000010001111001; // vC= 1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010101; // iC= 1429 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111110; // iC= 1406 
vC = 14'b0000010001110011; // vC= 1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011001; // iC= 1369 
vC = 14'b0000010001101111; // vC= 1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000110; // iC= 1350 
vC = 14'b0000010011000010; // vC= 1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111111; // iC= 1279 
vC = 14'b0000010001000111; // vC= 1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011100; // iC= 1244 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000010; // iC= 1346 
vC = 14'b0000010001010010; // vC= 1106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110011; // iC= 1331 
vC = 14'b0000010010101101; // vC= 1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001110; // iC= 1358 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101101; // iC= 1261 
vC = 14'b0000010001100000; // vC= 1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001100; // iC= 1292 
vC = 14'b0000010010110101; // vC= 1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010001; // iC= 1361 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011101; // iC= 1245 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010101; // iC= 1301 
vC = 14'b0000010011000010; // vC= 1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001111; // iC= 1295 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000100; // iC= 1220 
vC = 14'b0000010011011000; // vC= 1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110110; // iC= 1270 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000010100010110; // vC= 1302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010011; // iC= 1299 
vC = 14'b0000010010001101; // vC= 1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011110; // iC= 1246 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100101; // iC= 1253 
vC = 14'b0000010011010001; // vC= 1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001011; // iC= 1291 
vC = 14'b0000010010010011; // vC= 1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111010; // iC= 1274 
vC = 14'b0000010100010100; // vC= 1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001101; // iC= 1229 
vC = 14'b0000010011110100; // vC= 1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010111; // iC= 1175 
vC = 14'b0000010010101000; // vC= 1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100000; // iC= 1184 
vC = 14'b0000010011101010; // vC= 1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000000; // iC= 1280 
vC = 14'b0000010011011010; // vC= 1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001001; // iC= 1161 
vC = 14'b0000010011001100; // vC= 1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111001; // iC= 1209 
vC = 14'b0000010010100101; // vC= 1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010001; // iC= 1233 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100100; // iC= 1188 
vC = 14'b0000010100011110; // vC= 1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101100; // iC= 1132 
vC = 14'b0000010011110111; // vC= 1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011010; // iC= 1178 
vC = 14'b0000010100110110; // vC= 1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110000; // iC= 1200 
vC = 14'b0000010011100001; // vC= 1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000011; // iC= 1219 
vC = 14'b0000010011000100; // vC= 1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100001; // iC= 1249 
vC = 14'b0000010011001111; // vC= 1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101100; // iC= 1132 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111010; // iC= 1210 
vC = 14'b0000010100000111; // vC= 1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011011; // iC= 1243 
vC = 14'b0000010011001001; // vC= 1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101110; // iC= 1198 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110111; // iC= 1079 
vC = 14'b0000010100000000; // vC= 1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000011; // iC= 1155 
vC = 14'b0000010011101100; // vC= 1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101100; // iC= 1196 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000111; // iC= 1223 
vC = 14'b0000010100001000; // vC= 1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010111; // iC= 1111 
vC = 14'b0000010011101000; // vC= 1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010001; // iC= 1169 
vC = 14'b0000010100110000; // vC= 1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011111; // iC= 1055 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110000; // iC= 1136 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001000; // iC= 1096 
vC = 14'b0000010100011001; // vC= 1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010010; // iC= 1106 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100101; // iC= 1125 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011011; // iC= 1051 
vC = 14'b0000010110000100; // vC= 1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010100; // iC= 1044 
vC = 14'b0000010101110000; // vC= 1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011100; // iC= 1116 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010010; // iC= 1106 
vC = 14'b0000010100111001; // vC= 1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101011; // iC= 1067 
vC = 14'b0000010101010100; // vC= 1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001011; // iC= 1099 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011100; // iC= 1116 
vC = 14'b0000010100110010; // vC= 1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110001; // iC= 1137 
vC = 14'b0000010101010110; // vC= 1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101110; // iC= 1134 
vC = 14'b0000010110011110; // vC= 1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011110; // iC= 1054 
vC = 14'b0000010100010101; // vC= 1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110100; // iC= 1076 
vC = 14'b0000010110111000; // vC= 1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100001; // iC=  993 
vC = 14'b0000010101001110; // vC= 1358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101010; // iC= 1066 
vC = 14'b0000010100110011; // vC= 1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001111; // iC= 1103 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011000; // iC= 1048 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101110; // iC=  942 
vC = 14'b0000010110110010; // vC= 1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000010; // iC=  962 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101011; // iC=  939 
vC = 14'b0000010100110111; // vC= 1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110110; // iC=  950 
vC = 14'b0000010101011001; // vC= 1369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001000; // iC=  968 
vC = 14'b0000010101011100; // vC= 1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010111; // iC=  919 
vC = 14'b0000010101101011; // vC= 1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111110; // iC= 1022 
vC = 14'b0000010111000100; // vC= 1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100111; // iC=  999 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111111; // iC= 1023 
vC = 14'b0000010101011111; // vC= 1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110000; // iC=  944 
vC = 14'b0000010111001001; // vC= 1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101111; // iC= 1007 
vC = 14'b0000010110011010; // vC= 1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110000; // iC=  944 
vC = 14'b0000010111100010; // vC= 1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010111; // iC=  919 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110111; // iC=  887 
vC = 14'b0000010110001100; // vC= 1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010110; // iC=  982 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001000; // iC=  904 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110001; // iC=  945 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101010; // iC=  938 
vC = 14'b0000010101011110; // vC= 1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011001; // iC=  857 
vC = 14'b0000010111110111; // vC= 1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110000; // iC=  880 
vC = 14'b0000010111001000; // vC= 1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110100; // iC=  884 
vC = 14'b0000010110001000; // vC= 1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011101; // iC=  925 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010100; // iC=  916 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000011; // iC=  963 
vC = 14'b0000010110110000; // vC= 1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111101; // iC=  829 
vC = 14'b0000010101111110; // vC= 1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011000; // iC=  920 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001100; // iC=  908 
vC = 14'b0000010110100001; // vC= 1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101110; // iC=  878 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111111; // iC=  895 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101111; // iC=  815 
vC = 14'b0000010110010000; // vC= 1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011101; // iC=  925 
vC = 14'b0000010111100100; // vC= 1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b0000010110010111; // vC= 1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101100; // iC=  812 
vC = 14'b0000010110111110; // vC= 1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010010; // iC=  850 
vC = 14'b0000010111110010; // vC= 1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111000; // iC=  824 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010000; // iC=  784 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011100; // iC=  796 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100111; // iC=  743 
vC = 14'b0000010110110110; // vC= 1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000000; // iC=  896 
vC = 14'b0000010111001101; // vC= 1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000101; // iC=  837 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100001; // iC=  801 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100000; // iC=  800 
vC = 14'b0000010110110110; // vC= 1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100101; // iC=  805 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001110; // iC=  846 
vC = 14'b0000010110101000; // vC= 1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101110; // iC=  750 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001010; // iC=  714 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b0000010110100010; // vC= 1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111011; // iC=  699 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001010; // iC=  778 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110101; // iC=  757 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110110; // iC=  758 
vC = 14'b0000010111100001; // vC= 1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101000; // iC=  680 
vC = 14'b0000010111000101; // vC= 1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001001; // iC=  713 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101011; // iC=  683 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001110; // iC=  782 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110111; // iC=  759 
vC = 14'b0000010111010111; // vC= 1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011000; // iC=  664 
vC = 14'b0000010111000011; // vC= 1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111101; // iC=  701 
vC = 14'b0000010111110001; // vC= 1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110001; // iC=  753 
vC = 14'b0000010111010101; // vC= 1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110010; // iC=  690 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010111; // iC=  663 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100011; // iC=  739 
vC = 14'b0000010111011000; // vC= 1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110010; // iC=  626 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110110; // iC=  630 
vC = 14'b0000010111101100; // vC= 1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010111; // iC=  599 
vC = 14'b0000010111100111; // vC= 1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010010; // iC=  594 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101101; // iC=  685 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001010; // iC=  714 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100111; // iC=  615 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000011; // iC=  579 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011001; // iC=  601 
vC = 14'b0000011001011101; // vC= 1629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111110; // iC=  574 
vC = 14'b0000011001010010; // vC= 1618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101000; // iC=  616 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110010; // iC=  626 
vC = 14'b0000011000111000; // vC= 1592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010101; // iC=  597 
vC = 14'b0000011001010101; // vC= 1621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101001; // iC=  681 
vC = 14'b0000011001101100; // vC= 1644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001101; // iC=  589 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000110; // iC=  518 
vC = 14'b0000010111111000; // vC= 1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000100; // iC=  516 
vC = 14'b0000011001100100; // vC= 1636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000000; // iC=  512 
vC = 14'b0000011000001101; // vC= 1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001100; // iC=  588 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111110; // iC=  510 
vC = 14'b0000011000010111; // vC= 1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111111; // iC=  639 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000010; // iC=  514 
vC = 14'b0000010111101010; // vC= 1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100101; // iC=  549 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101100; // iC=  556 
vC = 14'b0000011000110100; // vC= 1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011100; // iC=  540 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000110; // iC=  518 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100101; // iC=  549 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111010; // iC=  506 
vC = 14'b0000011000110100; // vC= 1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010100; // iC=  596 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100101; // iC=  549 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000111; // iC=  455 
vC = 14'b0000011000101000; // vC= 1576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101011; // iC=  555 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010001; // iC=  529 
vC = 14'b0000010111110011; // vC= 1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001110; // iC=  526 
vC = 14'b0000010111111000; // vC= 1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010010; // iC=  530 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000110; // iC=  454 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010001; // iC=  465 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111110; // iC=  382 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111100; // iC=  508 
vC = 14'b0000010111110101; // vC= 1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100011; // iC=  355 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010000; // iC=  464 
vC = 14'b0000011010001011; // vC= 1675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110010; // iC=  370 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111101; // iC=  445 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000110; // iC=  390 
vC = 14'b0000011001100111; // vC= 1639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111100; // iC=  444 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001101; // iC=  269 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111110; // iC=  382 
vC = 14'b0000011010000000; // vC= 1664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010001; // iC=  337 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010101; // iC=  277 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000010; // iC=  322 
vC = 14'b0000011000110101; // vC= 1589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110010; // iC=  242 
vC = 14'b0000011000101100; // vC= 1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011011; // iC=  219 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000110; // iC=  198 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110010; // iC=  178 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100001; // iC=  225 
vC = 14'b0000011001111010; // vC= 1658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010000; // iC=  144 
vC = 14'b0000011000011001; // vC= 1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000011; // iC=  259 
vC = 14'b0000011001010100; // vC= 1620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100100; // iC=  228 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110101; // iC=  245 
vC = 14'b0000011010000110; // vC= 1670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001011; // iC=  203 
vC = 14'b0000011001100101; // vC= 1637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010000; // iC=  144 
vC = 14'b0000011001101100; // vC= 1644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000101; // iC=  133 
vC = 14'b0000011001011011; // vC= 1627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011000; // iC=  152 
vC = 14'b0000011000001101; // vC= 1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111100; // iC=  124 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011000; // iC=   24 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000111; // iC=   71 
vC = 14'b0000011001111001; // vC= 1657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111101; // iC=   61 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010110; // iC=   86 
vC = 14'b0000011010010010; // vC= 1682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111110; // iC=   -2 
vC = 14'b0000011001010111; // vC= 1623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111000; // iC=   56 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100111; // iC=  -25 
vC = 14'b0000011000101010; // vC= 1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110101; // iC=  -75 
vC = 14'b0000011000101011; // vC= 1579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101011; // iC=  -85 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100011; // iC= -157 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100001; // iC=  -31 
vC = 14'b0000011001100011; // vC= 1635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101100; // iC= -148 
vC = 14'b0000011000101010; // vC= 1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011111; // iC= -161 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001101; // iC= -243 
vC = 14'b0000011010001101; // vC= 1677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000100; // iC= -124 
vC = 14'b0000011001010110; // vC= 1622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011101; // iC= -227 
vC = 14'b0000011001100110; // vC= 1638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000100; // iC= -188 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011001; // iC= -295 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010001; // iC= -239 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000110; // iC= -378 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110010; // iC= -398 
vC = 14'b0000011001011001; // vC= 1625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111101; // iC= -323 
vC = 14'b0000011010000110; // vC= 1670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100001; // iC= -287 
vC = 14'b0000011001110010; // vC= 1650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001011; // iC= -309 
vC = 14'b0000011001110010; // vC= 1650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101000; // iC= -344 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000110; // iC= -506 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000010; // iC= -446 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100101; // iC= -475 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001011; // iC= -565 
vC = 14'b0000010111111111; // vC= 1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100010; // iC= -478 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001100; // iC= -564 
vC = 14'b0000011001101001; // vC= 1641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110000; // iC= -528 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110100; // iC= -524 
vC = 14'b0000010111011100; // vC= 1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101000; // iC= -600 
vC = 14'b0000010111110011; // vC= 1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011100; // iC= -612 
vC = 14'b0000011001100011; // vC= 1635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011110; // iC= -674 
vC = 14'b0000010111101001; // vC= 1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010111; // iC= -745 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010110; // iC= -618 
vC = 14'b0000010111011110; // vC= 1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110000; // iC= -720 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110010; // iC= -718 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110111; // iC= -713 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111010; // iC= -838 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000001; // iC= -767 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000000; // iC= -768 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100001; // iC= -863 
vC = 14'b0000011000010010; // vC= 1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000110; // iC= -826 
vC = 14'b0000011000011101; // vC= 1565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101000; // iC= -856 
vC = 14'b0000010111000010; // vC= 1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111001; // iC= -903 
vC = 14'b0000010111100011; // vC= 1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111100; // iC= -900 
vC = 14'b0000010111111111; // vC= 1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111000; // iC= -968 
vC = 14'b0000010110111111; // vC= 1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010000; // iC= -944 
vC = 14'b0000010111000101; // vC= 1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011101; // iC= -995 
vC = 14'b0000010111001011; // vC= 1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111011; // iC= -965 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011111; // iC= -929 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011101; // iC= -995 
vC = 14'b0000010101111111; // vC= 1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100100; // iC=-1116 
vC = 14'b0000010111110101; // vC= 1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010011; // iC=-1133 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000010; // iC=-1150 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110110; // iC=-1162 
vC = 14'b0000010111011100; // vC= 1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101100; // iC=-1044 
vC = 14'b0000010110110100; // vC= 1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011110; // iC=-1186 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110011; // iC=-1101 
vC = 14'b0000011000000001; // vC= 1537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000010; // iC=-1214 
vC = 14'b0000010101101100; // vC= 1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010000; // iC=-1136 
vC = 14'b0000010110010010; // vC= 1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110110; // iC=-1226 
vC = 14'b0000010110100000; // vC= 1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110001; // iC=-1167 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101011; // iC=-1173 
vC = 14'b0000010110010111; // vC= 1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b0000010101110111; // vC= 1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111111; // iC=-1217 
vC = 14'b0000010110111010; // vC= 1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100000; // iC=-1312 
vC = 14'b0000010101010101; // vC= 1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010110; // iC=-1322 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110101; // iC=-1291 
vC = 14'b0000010110010010; // vC= 1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b0000010111001001; // vC= 1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000000; // iC=-1344 
vC = 14'b0000010110100000; // vC= 1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000111; // iC=-1337 
vC = 14'b0000010100111001; // vC= 1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b0000010100010111; // vC= 1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111000; // iC=-1352 
vC = 14'b0000010101111110; // vC= 1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001111; // iC=-1393 
vC = 14'b0000010100010100; // vC= 1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b0000010101000000; // vC= 1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001110; // iC=-1394 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001110; // iC=-1394 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b0000010100101110; // vC= 1326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010111; // iC=-1449 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011000; // iC=-1512 
vC = 14'b0000010100000111; // vC= 1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b0000010101101110; // vC= 1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b0000010011111000; // vC= 1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b0000010100100111; // vC= 1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010111; // iC=-1449 
vC = 14'b0000010011001111; // vC= 1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b0000010011111001; // vC= 1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b0000010011101111; // vC= 1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b0000010011010001; // vC= 1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b0000010011110100; // vC= 1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b0000010100101001; // vC= 1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010010; // iC=-1518 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110111; // iC=-1545 
vC = 14'b0000010100111101; // vC= 1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001101; // iC=-1587 
vC = 14'b0000010011010011; // vC= 1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b0000010011000100; // vC= 1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000010011011010; // vC= 1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b0000010011001001; // vC= 1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b0000010001111100; // vC= 1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100011; // iC=-1565 
vC = 14'b0000010011111011; // vC= 1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000010011010001; // vC= 1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b0000010010100111; // vC= 1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b0000010011000010; // vC= 1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000010011010101; // vC= 1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100000; // iC=-1632 
vC = 14'b0000010011011000; // vC= 1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b0000010001101000; // vC= 1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b0000010001110010; // vC= 1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b0000010001101100; // vC= 1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b0000010011011100; // vC= 1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000010010110010; // vC= 1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b0000010001101100; // vC= 1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000111; // iC=-1657 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000010000111011; // vC= 1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000101; // iC=-1595 
vC = 14'b0000010000110110; // vC= 1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b0000010000100100; // vC= 1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011010; // iC=-1702 
vC = 14'b0000010000101110; // vC= 1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b0000010010000000; // vC= 1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b0000010000110001; // vC= 1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001111100101; // vC=  997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b0000010000111101; // vC= 1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b0000001111111111; // vC= 1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000010000010111; // vC= 1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b0000010001001000; // vC= 1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000001111010011; // vC=  979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000001111111110; // vC= 1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b0000001111111101; // vC= 1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000001110010011; // vC=  915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b0000001111111011; // vC= 1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b0000001110011001; // vC=  921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011101; // iC=-1699 
vC = 14'b0000001101111100; // vC=  892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000010000001010; // vC= 1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000001110101101; // vC=  941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000001110011100; // vC=  924 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000001111100001; // vC=  993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b0000001101010011; // vC=  851 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b0000001111100101; // vC=  997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001101110111; // vC=  887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000001101000001; // vC=  833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b0000001111000000; // vC=  960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101010; // iC=-1750 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111011; // iC=-1797 
vC = 14'b0000001101111011; // vC=  891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000001101111010; // vC=  890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000001101010100; // vC=  852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b0000001110001110; // vC=  910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000001101110100; // vC=  884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b0000001100100111; // vC=  807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000001100101001; // vC=  809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000001101101011; // vC=  875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000001101101010; // vC=  874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000001101000101; // vC=  837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000001101101101; // vC=  877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010000; // iC=-1840 
vC = 14'b0000001011110000; // vC=  752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000001101011110; // vC=  862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000001011110100; // vC=  756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000001100100101; // vC=  805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000001101000111; // vC=  839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000001100000010; // vC=  770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000001100110111; // vC=  823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000001011100011; // vC=  739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010000; // iC=-1840 
vC = 14'b0000001011101101; // vC=  749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000001100101000; // vC=  808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101001; // iC=-1815 
vC = 14'b0000001100000101; // vC=  773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b0000001100001111; // vC=  783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001010; // iC=-1846 
vC = 14'b0000001100011010; // vC=  794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111100; // iC=-1860 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b0000001010010101; // vC=  661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b0000001011010000; // vC=  720 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000001011010001; // vC=  721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b0000001001101000; // vC=  616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000001011000011; // vC=  707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111011; // iC=-1797 
vC = 14'b0000001001011111; // vC=  607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b0000001011001110; // vC=  718 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000001001111111; // vC=  639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000001011010000; // vC=  720 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000001001101100; // vC=  620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b0000001010100000; // vC=  672 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b0000001001011011; // vC=  603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000001000010001; // vC=  529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101010; // iC=-1750 
vC = 14'b0000001010011000; // vC=  664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000001001111110; // vC=  638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000001000001000; // vC=  520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001000101011; // vC=  555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010100; // iC=-1836 
vC = 14'b0000001000111010; // vC=  570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000001001000011; // vC=  579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000000111101111; // vC=  495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111111; // iC=-1857 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000001000111001; // vC=  569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000001000101001; // vC=  553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000000111011111; // vC=  479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110100; // iC=-1868 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000001000100001; // vC=  545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b0000001000101010; // vC=  554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000000111101001; // vC=  489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000001000110101; // vC=  565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101000; // iC=-1880 
vC = 14'b0000000111100001; // vC=  481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b0000000110011111; // vC=  415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010011; // iC=-1837 
vC = 14'b0000000110101011; // vC=  427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001111; // iC=-1841 
vC = 14'b0000000110011111; // vC=  415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000001000001001; // vC=  521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000000110011101; // vC=  413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000000111001001; // vC=  457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110000; // iC=-1872 
vC = 14'b0000000110011000; // vC=  408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000000101111111; // vC=  383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000000101011110; // vC=  350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b0000000110110011; // vC=  435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000000111100000; // vC=  480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111010; // iC=-1798 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000000110001101; // vC=  397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000000111001100; // vC=  460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000000101111011; // vC=  379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000101100001; // vC=  353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000110101001; // vC=  425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000110100111; // vC=  423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000110110000; // vC=  432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000000100101011; // vC=  299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000000101111100; // vC=  380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101111; // iC=-1873 
vC = 14'b0000000101011001; // vC=  345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111100; // iC=-1860 
vC = 14'b0000000100101010; // vC=  298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000000100011111; // vC=  287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000000100101000; // vC=  296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000000011100000; // vC=  224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000000100100001; // vC=  289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101001; // iC=-1815 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000000100110101; // vC=  309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000000100011101; // vC=  285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b0000000011101101; // vC=  237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b0000000010101111; // vC=  175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000000010111111; // vC=  191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b0000000011001111; // vC=  207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000000100100000; // vC=  288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111100; // iC=-1860 
vC = 14'b0000000010001111; // vC=  143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000000100010101; // vC=  277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000000011101000; // vC=  232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000000011100101; // vC=  229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110010; // iC=-1870 
vC = 14'b0000000011010110; // vC=  214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110110; // iC=-1866 
vC = 14'b0000000010011110; // vC=  158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000000010100011; // vC=  163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111010; // iC=-1798 
vC = 14'b0000000001010101; // vC=   85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000000000110011; // vC=   51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000000000111001; // vC=   57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000001101101; // vC=  109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b0000000010101011; // vC=  171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000000000010101; // vC=   21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000010; // iC=-1854 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000000000111011; // vC=   59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b1111111111111000; // vC=   -8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b0000000001101001; // vC=  105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b0000000000100011; // vC=   35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b1111111111100000; // vC=  -32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b0000000000111111; // vC=   63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b1111111111110000; // vC=  -16 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011010; // iC=-1830 
vC = 14'b0000000000011100; // vC=   28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011010; // iC=-1830 
vC = 14'b0000000000111111; // vC=   63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b1111111111111010; // vC=   -6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000000000101101; // vC=   45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000000000011001; // vC=   25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b1111111111010110; // vC=  -42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000000000110101; // vC=   53 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b1111111110011101; // vC=  -99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b1111111111110001; // vC=  -15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b1111111110100001; // vC=  -95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b1111111110000101; // vC= -123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b1111111111010100; // vC=  -44 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b1111111110100000; // vC=  -96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b1111111110100011; // vC=  -93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b1111111101100001; // vC= -159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b1111111111110010; // vC=  -14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b1111111111101110; // vC=  -18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b1111111101011101; // vC= -163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011110; // iC=-1698 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b1111111101000011; // vC= -189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b1111111101110111; // vC= -137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b1111111111000010; // vC=  -62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b1111111101110111; // vC= -137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b1111111101010000; // vC= -176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b1111111101011001; // vC= -167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b1111111101101100; // vC= -148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b1111111110100110; // vC=  -90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b1111111101100100; // vC= -156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b1111111100011000; // vC= -232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b1111111100101001; // vC= -215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b1111111011111000; // vC= -264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b1111111101010101; // vC= -171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b1111111101001110; // vC= -178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b1111111101010111; // vC= -169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b1111111101011111; // vC= -161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b1111111100000011; // vC= -253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111010; // iC=-1670 
vC = 14'b1111111011110001; // vC= -271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b1111111011100111; // vC= -281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001000; // iC=-1656 
vC = 14'b1111111100100010; // vC= -222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110000; // iC=-1680 
vC = 14'b1111111100010111; // vC= -233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101011; // iC=-1621 
vC = 14'b1111111100000100; // vC= -252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b1111111100000101; // vC= -251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b1111111011110011; // vC= -269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b1111111011110010; // vC= -270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b1111111010101111; // vC= -337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b1111111010101001; // vC= -343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b1111111011100110; // vC= -282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b1111111011111001; // vC= -263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000001; // iC=-1599 
vC = 14'b1111111010011010; // vC= -358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101000; // iC=-1688 
vC = 14'b1111111010100010; // vC= -350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b1111111010010111; // vC= -361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001101; // iC=-1651 
vC = 14'b1111111011111010; // vC= -262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001101; // iC=-1587 
vC = 14'b1111111011110100; // vC= -268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101101; // iC=-1619 
vC = 14'b1111111011110001; // vC= -271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b1111111001010101; // vC= -427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b1111111010010110; // vC= -362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100011; // iC=-1693 
vC = 14'b1111111010001100; // vC= -372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b1111111001100000; // vC= -416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b1111111001110011; // vC= -397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b1111111001100100; // vC= -412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b1111111010011001; // vC= -359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b1111111000100000; // vC= -480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b1111111001110001; // vC= -399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b1111111001011001; // vC= -423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b1111111000001111; // vC= -497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b1111111010011000; // vC= -360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b1111111000010010; // vC= -494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b1111111010001100; // vC= -372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001100; // iC=-1588 
vC = 14'b1111111001111101; // vC= -387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b1111111000100010; // vC= -478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100011; // iC=-1693 
vC = 14'b1111111001010001; // vC= -431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b1111111001111001; // vC= -391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100110; // iC=-1562 
vC = 14'b1111111001010010; // vC= -430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111111; // iC=-1537 
vC = 14'b1111111001001111; // vC= -433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010100; // iC=-1644 
vC = 14'b1111111000111101; // vC= -451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b1111110111000111; // vC= -569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b1111110111111110; // vC= -514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b1111110111110101; // vC= -523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b1111111000101011; // vC= -469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b1111110111001100; // vC= -564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011000; // iC=-1512 
vC = 14'b1111111000000000; // vC= -512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100011; // iC=-1565 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101111; // iC=-1553 
vC = 14'b1111110111001011; // vC= -565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100110; // iC=-1562 
vC = 14'b1111110111011011; // vC= -549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011101; // iC=-1571 
vC = 14'b1111110111000111; // vC= -569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b1111111000011011; // vC= -485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b1111111000001001; // vC= -503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100011; // iC=-1629 
vC = 14'b1111110111001111; // vC= -561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b1111110110000010; // vC= -638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b1111110111101100; // vC= -532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b1111110111010111; // vC= -553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b1111110111011010; // vC= -550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111001; // iC=-1607 
vC = 14'b1111110111110101; // vC= -523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b1111110111101101; // vC= -531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011101; // iC=-1507 
vC = 14'b1111110111100011; // vC= -541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b1111110101100010; // vC= -670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b1111110111000101; // vC= -571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b1111110101001001; // vC= -695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b1111110110111001; // vC= -583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b1111110110100110; // vC= -602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101111; // iC=-1553 
vC = 14'b1111110110001100; // vC= -628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010111; // iC=-1449 
vC = 14'b1111110110010111; // vC= -617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110111; // iC=-1481 
vC = 14'b1111110101010111; // vC= -681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b1111110100110010; // vC= -718 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000110; // iC=-1466 
vC = 14'b1111110100010100; // vC= -748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b1111110101110000; // vC= -656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b1111110101110000; // vC= -656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b1111110100010101; // vC= -747 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100011; // iC=-1437 
vC = 14'b1111110101111010; // vC= -646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100111; // iC=-1497 
vC = 14'b1111110110010001; // vC= -623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b1111110011110110; // vC= -778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b1111110110001001; // vC= -631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000011; // iC=-1533 
vC = 14'b1111110100001101; // vC= -755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b1111110011110011; // vC= -781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b1111110100110011; // vC= -717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100011; // iC=-1501 
vC = 14'b1111110101011000; // vC= -680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b1111110100101101; // vC= -723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010111; // iC=-1513 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b1111110100110110; // vC= -714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000100; // iC=-1468 
vC = 14'b1111110100001101; // vC= -755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b1111110100110100; // vC= -716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b1111110100100101; // vC= -731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111010; // iC=-1414 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010010; // iC=-1518 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011111; // iC=-1441 
vC = 14'b1111110011011110; // vC= -802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100110; // iC=-1370 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100011; // iC=-1373 
vC = 14'b1111110100110001; // vC= -719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b1111110100100011; // vC= -733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100110; // iC=-1434 
vC = 14'b1111110100000011; // vC= -765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100001; // iC=-1375 
vC = 14'b1111110100001001; // vC= -759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111110011001011; // vC= -821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100100; // iC=-1436 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110000; // iC=-1360 
vC = 14'b1111110010000011; // vC= -893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010111; // iC=-1321 
vC = 14'b1111110011100110; // vC= -794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101000; // iC=-1368 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100101; // iC=-1371 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b1111110010010101; // vC= -875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011011; // iC=-1317 
vC = 14'b1111110010011110; // vC= -866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011111; // iC=-1313 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100011; // iC=-1373 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011001; // iC=-1319 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001100; // iC=-1332 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011100; // iC=-1316 
vC = 14'b1111110001010001; // vC= -943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110111; // iC=-1353 
vC = 14'b1111110011010001; // vC= -815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b1111110011001100; // vC= -820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110010; // iC=-1422 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010101; // iC=-1323 
vC = 14'b1111110000110111; // vC= -969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001110; // iC=-1330 
vC = 14'b1111110011001100; // vC= -820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111110; // iC=-1346 
vC = 14'b1111110001101101; // vC= -915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101000; // iC=-1304 
vC = 14'b1111110000101100; // vC= -980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010101; // iC=-1387 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101101; // iC=-1363 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110110; // iC=-1290 
vC = 14'b1111110000011010; // vC= -998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011001; // iC=-1383 
vC = 14'b1111110001110101; // vC= -907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001111; // iC=-1393 
vC = 14'b1111110000111101; // vC= -963 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010010; // iC=-1326 
vC = 14'b1111110001001100; // vC= -948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101101; // iC=-1235 
vC = 14'b1111110001100100; // vC= -924 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010010; // iC=-1262 
vC = 14'b1111110010000011; // vC= -893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b1111110000100111; // vC= -985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100110; // iC=-1306 
vC = 14'b1111110001101000; // vC= -920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111101; // iC=-1347 
vC = 14'b1111110001001110; // vC= -946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101011; // iC=-1301 
vC = 14'b1111110000110100; // vC= -972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110000; // iC=-1232 
vC = 14'b1111110001110111; // vC= -905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111010; // iC=-1350 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000100; // iC=-1212 
vC = 14'b1111101111011101; // vC=-1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011110; // iC=-1250 
vC = 14'b1111110000010001; // vC=-1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000101; // iC=-1339 
vC = 14'b1111110000010111; // vC=-1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011111; // iC=-1249 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011110; // iC=-1314 
vC = 14'b1111110001011111; // vC= -929 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101100; // iC=-1172 
vC = 14'b1111110000000010; // vC=-1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b1111110001001000; // vC= -952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000100; // iC=-1276 
vC = 14'b1111101110111101; // vC=-1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111110; // iC=-1282 
vC = 14'b1111101111010100; // vC=-1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110110; // iC=-1290 
vC = 14'b1111101111010101; // vC=-1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000111; // iC=-1209 
vC = 14'b1111101111111111; // vC=-1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b1111110001001101; // vC= -947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000010; // iC=-1150 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000000; // iC=-1280 
vC = 14'b1111101111111101; // vC=-1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b1111110000011111; // vC= -993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001100; // iC=-1204 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111100; // iC=-1156 
vC = 14'b1111101110100001; // vC=-1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110011; // iC=-1229 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101000; // iC=-1240 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001100; // iC=-1140 
vC = 14'b1111101110010000; // vC=-1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b1111101110100100; // vC=-1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111100; // iC=-1156 
vC = 14'b1111101111000010; // vC=-1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b1111101111101110; // vC=-1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100110; // iC=-1178 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100011; // iC=-1181 
vC = 14'b1111101111100001; // vC=-1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110100; // iC=-1100 
vC = 14'b1111101110100111; // vC=-1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001001; // iC=-1207 
vC = 14'b1111101110111101; // vC=-1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010010; // iC=-1198 
vC = 14'b1111101110010011; // vC=-1133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001111; // iC=-1201 
vC = 14'b1111101101101011; // vC=-1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110010; // iC=-1166 
vC = 14'b1111101111000001; // vC=-1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010100; // iC=-1196 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100000; // iC=-1184 
vC = 14'b1111101111010101; // vC=-1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101011; // iC=-1109 
vC = 14'b1111101110111011; // vC=-1093 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010110; // iC=-1194 
vC = 14'b1111101110110010; // vC=-1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101100; // iC=-1172 
vC = 14'b1111101110100110; // vC=-1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110011; // iC=-1165 
vC = 14'b1111101111000010; // vC=-1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110001; // iC=-1103 
vC = 14'b1111101101100100; // vC=-1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000111; // iC=-1145 
vC = 14'b1111101110010000; // vC=-1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100110; // iC=-1050 
vC = 14'b1111101110010100; // vC=-1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010100; // iC=-1132 
vC = 14'b1111101101100101; // vC=-1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101001; // iC=-1047 
vC = 14'b1111101101010111; // vC=-1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110110; // iC=-1162 
vC = 14'b1111101101110010; // vC=-1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100111; // iC=-1113 
vC = 14'b1111101111000000; // vC=-1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100010; // iC=-1118 
vC = 14'b1111101110100000; // vC=-1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001111; // iC=-1073 
vC = 14'b1111101101111010; // vC=-1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000000; // iC=-1024 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111101110111001; // vC=-1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011111; // iC=-1121 
vC = 14'b1111101101101111; // vC=-1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010111; // iC=-1129 
vC = 14'b1111101100100100; // vC=-1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110100; // iC= -972 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110001; // iC= -975 
vC = 14'b1111101101000010; // vC=-1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010001; // iC=-1071 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101001; // iC= -983 
vC = 14'b1111101110100000; // vC=-1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011111; // iC= -993 
vC = 14'b1111101101110101; // vC=-1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100111; // iC= -985 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000111; // iC=-1017 
vC = 14'b1111101110011001; // vC=-1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011111; // iC= -993 
vC = 14'b1111101101000101; // vC=-1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001000; // iC=-1080 
vC = 14'b1111101101111110; // vC=-1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001000; // iC=-1080 
vC = 14'b1111101101000010; // vC=-1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100100; // iC=-1052 
vC = 14'b1111101100111000; // vC=-1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001000; // iC=-1016 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110000; // iC= -912 
vC = 14'b1111101100001010; // vC=-1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b1111101011110010; // vC=-1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101101; // iC= -979 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010001; // iC=-1007 
vC = 14'b1111101101000110; // vC=-1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000111; // iC=-1017 
vC = 14'b1111101100000011; // vC=-1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000110; // iC= -954 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110110; // iC=-1034 
vC = 14'b1111101100110000; // vC=-1232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011001; // iC= -935 
vC = 14'b1111101100110001; // vC=-1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110011; // iC= -973 
vC = 14'b1111101101010011; // vC=-1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010000; // iC=-1008 
vC = 14'b1111101100000101; // vC=-1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101011; // iC= -981 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110110; // iC= -906 
vC = 14'b1111101011100010; // vC=-1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110100; // iC= -908 
vC = 14'b1111101011011001; // vC=-1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110010; // iC= -910 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001011; // iC= -885 
vC = 14'b1111101101001100; // vC=-1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011101; // iC= -867 
vC = 14'b1111101100000101; // vC=-1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000011; // iC= -893 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000001; // iC= -959 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111000; // iC= -840 
vC = 14'b1111101010110011; // vC=-1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001011; // iC= -949 
vC = 14'b1111101100111010; // vC=-1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011100; // iC= -868 
vC = 14'b1111101011100011; // vC=-1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110000; // iC= -848 
vC = 14'b1111101100011111; // vC=-1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100011; // iC= -925 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101011; // iC= -789 
vC = 14'b1111101100101001; // vC=-1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111100; // iC= -900 
vC = 14'b1111101010111101; // vC=-1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101010; // iC= -854 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100010; // iC= -862 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110011; // iC= -845 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000010; // iC= -830 
vC = 14'b1111101100011001; // vC=-1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100111; // iC= -857 
vC = 14'b1111101010001110; // vC=-1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001000; // iC= -760 
vC = 14'b1111101011111111; // vC=-1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101110; // iC= -786 
vC = 14'b1111101011110101; // vC=-1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011010; // iC= -870 
vC = 14'b1111101100010010; // vC=-1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001101; // iC= -755 
vC = 14'b1111101010010101; // vC=-1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010010; // iC= -878 
vC = 14'b1111101010000110; // vC=-1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010111; // iC= -809 
vC = 14'b1111101100010001; // vC=-1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010101; // iC= -811 
vC = 14'b1111101010010100; // vC=-1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111101011111010; // vC=-1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100101; // iC= -795 
vC = 14'b1111101010100100; // vC=-1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111001; // iC= -775 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001011; // iC= -757 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111010; // iC= -710 
vC = 14'b1111101011001001; // vC=-1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110010; // iC= -846 
vC = 14'b1111101011010001; // vC=-1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101110; // iC= -722 
vC = 14'b1111101011100101; // vC=-1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110010; // iC= -782 
vC = 14'b1111101011011000; // vC=-1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111100; // iC= -708 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010010; // iC= -686 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100001; // iC= -671 
vC = 14'b1111101001110011; // vC=-1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011000; // iC= -744 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110000; // iC= -720 
vC = 14'b1111101010011100; // vC=-1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001000; // iC= -760 
vC = 14'b1111101010111100; // vC=-1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101000; // iC= -728 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101011; // iC= -725 
vC = 14'b1111101010110001; // vC=-1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110110; // iC= -650 
vC = 14'b1111101001101111; // vC=-1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010010; // iC= -686 
vC = 14'b1111101011011011; // vC=-1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100011; // iC= -669 
vC = 14'b1111101010001011; // vC=-1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100000; // iC= -608 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000100; // iC= -700 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101111; // iC= -657 
vC = 14'b1111101011010011; // vC=-1325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100011; // iC= -733 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010101; // iC= -619 
vC = 14'b1111101010010010; // vC=-1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000001; // iC= -703 
vC = 14'b1111101000110110; // vC=-1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100011; // iC= -605 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110000; // iC= -656 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010110; // iC= -618 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011100; // iC= -612 
vC = 14'b1111101011001011; // vC=-1333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111100; // iC= -708 
vC = 14'b1111101010110010; // vC=-1358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000111; // iC= -633 
vC = 14'b1111101011000010; // vC=-1342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100100; // iC= -604 
vC = 14'b1111101010110100; // vC=-1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011110; // iC= -546 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011011; // iC= -613 
vC = 14'b1111101001101001; // vC=-1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001101; // iC= -563 
vC = 14'b1111101000110110; // vC=-1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110100; // iC= -524 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100010; // iC= -670 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001010; // iC= -566 
vC = 14'b1111101000110110; // vC=-1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101011; // iC= -661 
vC = 14'b1111101001001101; // vC=-1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110000; // iC= -656 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111111; // iC= -641 
vC = 14'b1111101001010001; // vC=-1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011100; // iC= -484 
vC = 14'b1111101000110000; // vC=-1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110101; // iC= -587 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110001; // iC= -527 
vC = 14'b1111101000011011; // vC=-1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010100; // iC= -492 
vC = 14'b1111101001111011; // vC=-1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100100; // iC= -476 
vC = 14'b1111101010100111; // vC=-1369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100110; // iC= -602 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100100; // iC= -540 
vC = 14'b1111101010011100; // vC=-1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000010; // iC= -510 
vC = 14'b1111101001110110; // vC=-1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111101; // iC= -451 
vC = 14'b1111101010000010; // vC=-1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010001; // iC= -495 
vC = 14'b1111101001001101; // vC=-1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101110; // iC= -530 
vC = 14'b1111101010000011; // vC=-1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001010; // iC= -438 
vC = 14'b1111101010010001; // vC=-1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110100; // iC= -460 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100101; // iC= -475 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011110; // iC= -418 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000110; // iC= -506 
vC = 14'b1111101001000100; // vC=-1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100011; // iC= -477 
vC = 14'b1111101001101100; // vC=-1428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100001; // iC= -415 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101011; // iC= -405 
vC = 14'b1111101000011111; // vC=-1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001110; // iC= -370 
vC = 14'b1111101001000110; // vC=-1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001101; // iC= -435 
vC = 14'b1111101000000000; // vC=-1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101011; // iC= -405 
vC = 14'b1111100111110000; // vC=-1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010100; // iC= -428 
vC = 14'b1111101001011110; // vC=-1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001010; // iC= -438 
vC = 14'b1111101000011100; // vC=-1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001111; // iC= -433 
vC = 14'b1111100111101011; // vC=-1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010001; // iC= -303 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100111; // iC= -409 
vC = 14'b1111100111110110; // vC=-1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000110; // iC= -314 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001001; // iC= -311 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000001; // iC= -319 
vC = 14'b1111101000001000; // vC=-1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001100; // iC= -308 
vC = 14'b1111101000101111; // vC=-1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001100; // iC= -244 
vC = 14'b1111100111101001; // vC=-1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010001; // iC= -303 
vC = 14'b1111101000001010; // vC=-1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111000; // iC= -328 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111001; // iC= -199 
vC = 14'b1111101000010100; // vC=-1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110010; // iC= -206 
vC = 14'b1111101000011010; // vC=-1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001111; // iC= -305 
vC = 14'b1111101001110110; // vC=-1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011100; // iC= -228 
vC = 14'b1111101001010100; // vC=-1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100011; // iC= -157 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010101; // iC= -235 
vC = 14'b1111100111110110; // vC=-1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111010; // iC= -134 
vC = 14'b1111101000001001; // vC=-1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011111; // iC= -161 
vC = 14'b1111100111111000; // vC=-1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110001; // iC= -143 
vC = 14'b1111100111111011; // vC=-1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000101; // iC= -187 
vC = 14'b1111100111100111; // vC=-1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111001; // iC=  -71 
vC = 14'b1111100111101001; // vC=-1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110011; // iC= -141 
vC = 14'b1111101001011110; // vC=-1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100010; // iC=  -30 
vC = 14'b1111101001101111; // vC=-1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010100; // iC=  -44 
vC = 14'b1111101000110101; // vC=-1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011001; // iC=   25 
vC = 14'b1111101001011000; // vC=-1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110111; // iC=   -9 
vC = 14'b1111100111111001; // vC=-1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100001; // iC=  -95 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111001; // iC=   -7 
vC = 14'b1111101000111011; // vC=-1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010110; // iC=   22 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101100; // iC=   44 
vC = 14'b1111100111110000; // vC=-1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101001; // iC=  105 
vC = 14'b1111101001101111; // vC=-1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111001; // iC=  121 
vC = 14'b1111101001110101; // vC=-1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011100; // iC=  156 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111101; // iC=   61 
vC = 14'b1111101000011010; // vC=-1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101110; // iC=  174 
vC = 14'b1111100111110110; // vC=-1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010010; // iC=  210 
vC = 14'b1111101000000011; // vC=-1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101001; // iC=  233 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001110; // iC=  206 
vC = 14'b1111101000111011; // vC=-1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100010; // iC=  290 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001100; // iC=  204 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101101; // iC=  237 
vC = 14'b1111100111011110; // vC=-1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011110; // iC=  286 
vC = 14'b1111101000100111; // vC=-1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011000; // iC=  280 
vC = 14'b1111101000011100; // vC=-1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110111; // iC=  375 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100011; // iC=  419 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101000; // iC=  360 
vC = 14'b1111101000010001; // vC=-1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101101; // iC=  429 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010110; // iC=  406 
vC = 14'b1111100111111000; // vC=-1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010011; // iC=  531 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101001; // iC=  489 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010101; // iC=  597 
vC = 14'b1111101000011010; // vC=-1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010111; // iC=  471 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100011; // iC=  611 
vC = 14'b1111101000000010; // vC=-1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111110; // iC=  510 
vC = 14'b1111101001110110; // vC=-1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101111; // iC=  623 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000011; // iC=  579 
vC = 14'b1111101010000000; // vC=-1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100111; // iC=  615 
vC = 14'b1111101000011001; // vC=-1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100110; // iC=  614 
vC = 14'b1111101010001101; // vC=-1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000001; // iC=  705 
vC = 14'b1111101010010010; // vC=-1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101011; // iC=  747 
vC = 14'b1111101010011101; // vC=-1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100100; // iC=  740 
vC = 14'b1111101000100111; // vC=-1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011001; // iC=  729 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001011; // iC=  843 
vC = 14'b1111101001001111; // vC=-1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110101; // iC=  821 
vC = 14'b1111101001111110; // vC=-1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100010; // iC=  802 
vC = 14'b1111101000010010; // vC=-1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010111; // iC=  919 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101000; // iC=  808 
vC = 14'b1111101001110100; // vC=-1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100101; // iC=  933 
vC = 14'b1111101010010110; // vC=-1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011110; // iC=  990 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010001; // iC=  977 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100110; // iC=  998 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110101; // iC=  949 
vC = 14'b1111101010000000; // vC=-1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100110; // iC=  998 
vC = 14'b1111101010110100; // vC=-1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101101; // iC= 1005 
vC = 14'b1111101010001101; // vC=-1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011001; // iC= 1049 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100000; // iC= 1056 
vC = 14'b1111101000111111; // vC=-1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111001; // iC= 1017 
vC = 14'b1111101011010011; // vC=-1325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101111; // iC= 1199 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000111; // iC= 1095 
vC = 14'b1111101010110101; // vC=-1355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000010; // iC= 1218 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101101; // iC= 1133 
vC = 14'b1111101001110101; // vC=-1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101001; // iC= 1129 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101000; // iC= 1192 
vC = 14'b1111101010111011; // vC=-1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110110; // iC= 1270 
vC = 14'b1111101001101000; // vC=-1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b1111101011101000; // vC=-1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110111; // iC= 1335 
vC = 14'b1111101011001000; // vC=-1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111010; // iC= 1274 
vC = 14'b1111101011011111; // vC=-1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001100; // iC= 1356 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001000; // iC= 1288 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110010; // iC= 1330 
vC = 14'b1111101011100010; // vC=-1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100001; // iC= 1377 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000111; // iC= 1351 
vC = 14'b1111101010001101; // vC=-1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101100; // iC= 1324 
vC = 14'b1111101010101100; // vC=-1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101010; // iC= 1450 
vC = 14'b1111101011100100; // vC=-1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100000; // iC= 1440 
vC = 14'b1111101011010010; // vC=-1326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100101; // iC= 1509 
vC = 14'b1111101011100011; // vC=-1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000010; // iC= 1474 
vC = 14'b1111101100010010; // vC=-1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001100; // iC= 1484 
vC = 14'b1111101100100100; // vC=-1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100011; // iC= 1443 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110100; // iC= 1524 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110111; // iC= 1527 
vC = 14'b1111101011100110; // vC=-1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110110; // iC= 1526 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b1111101011101110; // vC=-1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110111; // iC= 1527 
vC = 14'b1111101101010101; // vC=-1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b1111101011110100; // vC=-1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b1111101101010110; // vC=-1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100101; // iC= 1637 
vC = 14'b1111101101011000; // vC=-1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111111; // iC= 1663 
vC = 14'b1111101011110110; // vC=-1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000010; // iC= 1730 
vC = 14'b1111101100001100; // vC=-1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100101; // iC= 1637 
vC = 14'b1111101100010000; // vC=-1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b1111101100000010; // vC=-1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100100; // iC= 1636 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b1111101101111100; // vC=-1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b1111101101010000; // vC=-1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100101; // iC= 1765 
vC = 14'b1111101101011100; // vC=-1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000010; // iC= 1730 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b1111101100010011; // vC=-1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b1111101101111000; // vC=-1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b1111101100101100; // vC=-1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b1111101110100001; // vC=-1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011011; // iC= 1819 
vC = 14'b1111101101101000; // vC=-1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b1111101101011101; // vC=-1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011111; // iC= 1759 
vC = 14'b1111101111010110; // vC=-1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101011; // iC= 1835 
vC = 14'b1111101101011110; // vC=-1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011100; // iC= 1820 
vC = 14'b1111101111001011; // vC=-1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110100; // iC= 1780 
vC = 14'b1111101101110010; // vC=-1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b1111101101011010; // vC=-1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100000; // iC= 1824 
vC = 14'b1111101111001001; // vC=-1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b1111101111101110; // vC=-1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111011; // iC= 1851 
vC = 14'b1111101101101100; // vC=-1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111100; // iC= 1788 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b1111101110101100; // vC=-1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011100; // iC= 1884 
vC = 14'b1111101111001011; // vC=-1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b1111101111101001; // vC=-1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111101111010100; // vC=-1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111101110101011; // vC=-1109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b1111101111100111; // vC=-1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111101111000001; // vC=-1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101101; // iC= 1837 
vC = 14'b1111110001000111; // vC= -953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111110000101011; // vC= -981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101010; // iC= 1898 
vC = 14'b1111101111010101; // vC=-1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b1111101111110110; // vC=-1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b1111110000000100; // vC=-1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111101111110011; // vC=-1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111110000111001; // vC= -967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b1111110001011111; // vC= -929 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110000000001; // vC=-1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000111; // iC= 1991 
vC = 14'b1111110001011001; // vC= -935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111110000010000; // vC=-1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111110010000100; // vC= -892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b1111110010110101; // vC= -843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111110001101010; // vC= -918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111110010100000; // vC= -864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111110010001000; // vC= -888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b1111110001111011; // vC= -901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b1111110011000111; // vC= -825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111110010100011; // vC= -861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111110010000001; // vC= -895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111110100000011; // vC= -765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111110011010111; // vC= -809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111110010111000; // vC= -840 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100011; // iC= 2019 
vC = 14'b1111110101000011; // vC= -701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b1111110100001000; // vC= -760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111110100110111; // vC= -713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111110100000111; // vC= -761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111110100000011; // vC= -765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000001; // iC= 2049 
vC = 14'b1111110101010101; // vC= -683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000001; // iC= 2049 
vC = 14'b1111110100001101; // vC= -755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b1111110011101000; // vC= -792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111110101110101; // vC= -651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b1111110101001001; // vC= -695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111110100001001; // vC= -759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b1111110101011010; // vC= -678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b1111110101010001; // vC= -687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001100; // iC= 2060 
vC = 14'b1111110101001001; // vC= -695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b1111110110010010; // vC= -622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111110101100001; // vC= -671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000101; // iC= 2053 
vC = 14'b1111110110101110; // vC= -594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000001; // iC= 2049 
vC = 14'b1111110110000001; // vC= -639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111110101111111; // vC= -641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110101010011; // vC= -685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b1111110110001001; // vC= -631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001110; // iC= 2062 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b1111110111011111; // vC= -545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001111; // iC= 2063 
vC = 14'b1111110110101100; // vC= -596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000010; // iC= 2050 
vC = 14'b1111110110100111; // vC= -601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b1111110101111010; // vC= -646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111110101100011; // vC= -669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b1111110110100100; // vC= -604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111110111110010; // vC= -526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111110111111100; // vC= -516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b1111110111110010; // vC= -526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111110111100101; // vC= -539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011001; // iC= 2073 
vC = 14'b1111110110100111; // vC= -601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110111111010; // vC= -518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b1111110111111001; // vC= -519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111000111110; // vC= -450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001100; // iC= 2060 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b1111110110110100; // vC= -588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b1111111000000100; // vC= -508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111111000000110; // vC= -506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111111000011100; // vC= -484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111110111011111; // vC= -545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111110111110000; // vC= -528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111111001100000; // vC= -416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111110111111110; // vC= -514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001111; // iC= 2063 
vC = 14'b1111111001111100; // vC= -388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111111000001010; // vC= -502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111111000000000; // vC= -512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010011; // iC= 2067 
vC = 14'b1111111001001000; // vC= -440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b1111111001110101; // vC= -395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111111010011101; // vC= -355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010100; // iC= 2068 
vC = 14'b1111111001000010; // vC= -446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111111000011111; // vC= -481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100011; // iC= 2083 
vC = 14'b1111111000110101; // vC= -459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000011; // iC= 2051 
vC = 14'b1111111001110111; // vC= -393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100011; // iC= 2019 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111111000110010; // vC= -462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111111001001111; // vC= -433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000000; // iC= 2048 
vC = 14'b1111111010010100; // vC= -364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000100; // iC= 1924 
vC = 14'b1111111010001001; // vC= -375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000010; // iC= 2050 
vC = 14'b1111111010001000; // vC= -376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b1111111010000100; // vC= -380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111111001110101; // vC= -395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111111010000011; // vC= -381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111111011110101; // vC= -267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111111010100110; // vC= -346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000011; // iC= 2051 
vC = 14'b1111111011011011; // vC= -293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100101; // iC= 2021 
vC = 14'b1111111100011101; // vC= -227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111111100000101; // vC= -251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111000; // iC= 2040 
vC = 14'b1111111011110111; // vC= -265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111111100101011; // vC= -213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b1111111011101100; // vC= -276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111000; // iC= 2040 
vC = 14'b1111111100010010; // vC= -238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011101; // iC= 2077 
vC = 14'b1111111011010111; // vC= -297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111111011110101; // vC= -267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111111100111010; // vC= -198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b1111111011101110; // vC= -274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111111100001000; // vC= -248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111111100000001; // vC= -255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b1111111100011011; // vC= -229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111111101100010; // vC= -158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010101; // iC= 2069 
vC = 14'b1111111100110101; // vC= -203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011001; // iC= 2073 
vC = 14'b1111111110001011; // vC= -117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011101; // iC= 2077 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111111100101110; // vC= -210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111110100100; // vC=  -92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b1111111100110000; // vC= -208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001001; // iC= 2057 
vC = 14'b1111111110010101; // vC= -107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110100; // iC= 1972 
vC = 14'b1111111101110110; // vC= -138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100001; // iC= 2017 
vC = 14'b1111111101101111; // vC= -145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111111101000101; // vC= -187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111000; // iC= 2040 
vC = 14'b1111111110101011; // vC=  -85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111101100000; // vC= -160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b1111111111100001; // vC=  -31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b1111111101110111; // vC= -137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100010; // iC= 2018 
vC = 14'b1111111110110011; // vC=  -77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b1111111111111001; // vC=   -7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b1111111110100011; // vC=  -93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b0000000000000111; // vC=    7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001011; // iC= 2059 
vC = 14'b0000000000100101; // vC=   37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b1111111111000100; // vC=  -60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b0000000000001110; // vC=   14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b0000000000001001; // vC=    9 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111111111011101; // vC=  -35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111111110110101; // vC=  -75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b0000000000010110; // vC=   22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111111010001; // vC=  -47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b0000000000101010; // vC=   42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b0000000001011100; // vC=   92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b0000000000100100; // vC=   36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b0000000000001111; // vC=   15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b0000000000100000; // vC=   32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101101; // iC= 2029 
vC = 14'b0000000010000101; // vC=  133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b0000000001111010; // vC=  122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100011; // iC= 2019 
vC = 14'b0000000011000101; // vC=  197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b0000000011010010; // vC=  210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b0000000011001111; // vC=  207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b0000000010111011; // vC=  187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b0000000011001000; // vC=  200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011100; // iC= 1884 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b0000000010110111; // vC=  183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b0000000010000011; // vC=  131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b0000000011111100; // vC=  252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010100; // iC= 1876 
vC = 14'b0000000011001010; // vC=  202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b0000000010001011; // vC=  139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b0000000100010101; // vC=  277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b0000000011100101; // vC=  229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110010; // iC= 1906 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000010111001; // vC=  185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b0000000010011000; // vC=  152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b0000000100100100; // vC=  292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b0000000101001101; // vC=  333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b0000000101000011; // vC=  323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101100; // iC= 1964 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b0000000011000110; // vC=  198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b0000000101010111; // vC=  343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b0000000011110011; // vC=  243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b0000000101010010; // vC=  338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b0000000011100011; // vC=  227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b0000000101111101; // vC=  381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b0000000100100100; // vC=  292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b0000000101001110; // vC=  334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b0000000100000100; // vC=  260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b0000000110001010; // vC=  394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b0000000100100001; // vC=  289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001111; // iC= 1871 
vC = 14'b0000000100111111; // vC=  319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b0000000101000101; // vC=  325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b0000000100111001; // vC=  313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000101011011; // vC=  347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011011; // iC= 1819 
vC = 14'b0000000101101101; // vC=  365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b0000000110111000; // vC=  440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b0000000110000010; // vC=  386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b0000000110101001; // vC=  425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b0000000110101011; // vC=  427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111001; // iC= 1849 
vC = 14'b0000000110000010; // vC=  386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b0000000101010011; // vC=  339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b0000000101101010; // vC=  362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001011; // iC= 1867 
vC = 14'b0000000101110000; // vC=  368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b0000000110111100; // vC=  444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b0000000111011010; // vC=  474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b0000000111110110; // vC=  502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000111; // iC= 1863 
vC = 14'b0000000110101111; // vC=  431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111011; // iC= 1851 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b0000000110111100; // vC=  444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b0000000110001111; // vC=  399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101101; // iC= 1837 
vC = 14'b0000000111100001; // vC=  481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b0000000111010100; // vC=  468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b0000000111010010; // vC=  466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101000; // iC= 1832 
vC = 14'b0000001000011010; // vC=  538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100011; // iC= 1827 
vC = 14'b0000001000000101; // vC=  517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010101; // iC= 1749 
vC = 14'b0000000110110000; // vC=  432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001011; // iC= 1867 
vC = 14'b0000001000111010; // vC=  570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000001000001100; // vC=  524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011000; // iC= 1752 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001111; // iC= 1871 
vC = 14'b0000001000101010; // vC=  554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000001001100111; // vC=  615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b0000001000101100; // vC=  556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b0000001000101111; // vC=  559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100101; // iC= 1765 
vC = 14'b0000001000110010; // vC=  562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100010; // iC= 1762 
vC = 14'b0000001001110101; // vC=  629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b0000001001111111; // vC=  639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b0000001000001100; // vC=  524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000011; // iC= 1859 
vC = 14'b0000001010100000; // vC=  672 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b0000001010010110; // vC=  662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b0000001010001100; // vC=  652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b0000001001101011; // vC=  619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110001; // iC= 1777 
vC = 14'b0000001010100111; // vC=  679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b0000001001010010; // vC=  594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101101; // iC= 1709 
vC = 14'b0000001000110100; // vC=  564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100011; // iC= 1763 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b0000001011011010; // vC=  730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000001; // iC= 1729 
vC = 14'b0000001011010111; // vC=  727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b0000001010011010; // vC=  666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111010; // iC= 1658 
vC = 14'b0000001011001101; // vC=  717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b0000001011011100; // vC=  732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010010; // iC= 1682 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110000; // iC= 1776 
vC = 14'b0000001011101101; // vC=  749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101001; // iC= 1705 
vC = 14'b0000001100011110; // vC=  798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101101; // iC= 1645 
vC = 14'b0000001011100101; // vC=  741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000110; // iC= 1734 
vC = 14'b0000001010100100; // vC=  676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b0000001011110000; // vC=  752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b0000001010100101; // vC=  677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110000; // iC= 1776 
vC = 14'b0000001100111100; // vC=  828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b0000001011111100; // vC=  764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001110; // iC= 1678 
vC = 14'b0000001100000110; // vC=  774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110011; // iC= 1651 
vC = 14'b0000001011010111; // vC=  727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000001011101100; // vC=  748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101101; // iC= 1709 
vC = 14'b0000001100100010; // vC=  802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110101; // iC= 1653 
vC = 14'b0000001010111110; // vC=  702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110101; // iC= 1653 
vC = 14'b0000001101001100; // vC=  844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001010; // iC= 1610 
vC = 14'b0000001101100011; // vC=  867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001110; // iC= 1742 
vC = 14'b0000001101100110; // vC=  870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b0000001011110010; // vC=  754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110011; // iC= 1651 
vC = 14'b0000001011111000; // vC=  760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110111; // iC= 1591 
vC = 14'b0000001100111111; // vC=  831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b0000001101101001; // vC=  873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001110000001; // vC=  897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101011; // iC= 1643 
vC = 14'b0000001100111000; // vC=  824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010111; // iC= 1623 
vC = 14'b0000001101001101; // vC=  845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b0000001100001101; // vC=  781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001110001010; // vC=  906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010000; // iC= 1552 
vC = 14'b0000001101011110; // vC=  862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101110; // iC= 1646 
vC = 14'b0000001101101111; // vC=  879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000001110010000; // vC=  912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100111; // iC= 1703 
vC = 14'b0000001101011001; // vC=  857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001011; // iC= 1611 
vC = 14'b0000001110110101; // vC=  949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000110; // iC= 1606 
vC = 14'b0000001101100010; // vC=  866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100010; // iC= 1634 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b0000001110000110; // vC=  902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100110; // iC= 1638 
vC = 14'b0000001111010100; // vC=  980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110000; // iC= 1584 
vC = 14'b0000001100111111; // vC=  831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b0000001111001100; // vC=  972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000001110100000; // vC=  928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001110; // iC= 1550 
vC = 14'b0000001110100100; // vC=  932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111010; // iC= 1658 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010110; // iC= 1558 
vC = 14'b0000001110000001; // vC=  897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b0000001110101111; // vC=  943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b0000001101100001; // vC=  865 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110000; // iC= 1648 
vC = 14'b0000001111101110; // vC= 1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101101; // iC= 1517 
vC = 14'b0000001111111110; // vC= 1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100111; // iC= 1575 
vC = 14'b0000001110100110; // vC=  934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110111; // iC= 1527 
vC = 14'b0000001111110011; // vC= 1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b0000010000000100; // vC= 1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111001; // iC= 1593 
vC = 14'b0000001111010110; // vC=  982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b0000001110001010; // vC=  906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010000; // iC= 1616 
vC = 14'b0000001111111010; // vC= 1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010010; // iC= 1554 
vC = 14'b0000001111100100; // vC=  996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101101; // iC= 1517 
vC = 14'b0000001110101100; // vC=  940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001110; // iC= 1486 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011100; // iC= 1564 
vC = 14'b0000001110101100; // vC=  940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100000; // iC= 1568 
vC = 14'b0000001110101100; // vC=  940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111011; // iC= 1531 
vC = 14'b0000001111110010; // vC= 1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101011; // iC= 1451 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101000; // iC= 1448 
vC = 14'b0000010000100000; // vC= 1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111100; // iC= 1532 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010011; // iC= 1491 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111110; // iC= 1406 
vC = 14'b0000001111100110; // vC=  998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b0000010001011001; // vC= 1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001101; // iC= 1485 
vC = 14'b0000001111010100; // vC=  980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110011; // iC= 1523 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001010; // iC= 1418 
vC = 14'b0000010001000111; // vC= 1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101100; // iC= 1452 
vC = 14'b0000010000010001; // vC= 1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110010; // iC= 1458 
vC = 14'b0000010001101111; // vC= 1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100101; // iC= 1381 
vC = 14'b0000010001111111; // vC= 1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101011; // iC= 1515 
vC = 14'b0000001111110100; // vC= 1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000011; // iC= 1411 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010010; // iC= 1490 
vC = 14'b0000010000100110; // vC= 1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b0000010001111001; // vC= 1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101011; // iC= 1515 
vC = 14'b0000010000100000; // vC= 1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100000; // iC= 1504 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001111; // iC= 1359 
vC = 14'b0000010000110100; // vC= 1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011001; // iC= 1497 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000001; // iC= 1345 
vC = 14'b0000010001110110; // vC= 1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001110; // iC= 1358 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010101; // iC= 1365 
vC = 14'b0000010010101100; // vC= 1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011010; // iC= 1370 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100011; // iC= 1379 
vC = 14'b0000010001000001; // vC= 1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010111; // iC= 1431 
vC = 14'b0000010000111101; // vC= 1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010110; // iC= 1302 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001000; // iC= 1416 
vC = 14'b0000010010100010; // vC= 1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010101; // iC= 1429 
vC = 14'b0000010001111000; // vC= 1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111110; // iC= 1342 
vC = 14'b0000010010001101; // vC= 1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001110; // iC= 1358 
vC = 14'b0000010001110111; // vC= 1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101011; // iC= 1323 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011001; // iC= 1305 
vC = 14'b0000010001110011; // vC= 1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010111; // iC= 1367 
vC = 14'b0000010011100111; // vC= 1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010001; // iC= 1361 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111011; // iC= 1275 
vC = 14'b0000010011110100; // vC= 1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101110; // iC= 1262 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101111; // iC= 1263 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001111; // iC= 1359 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000011; // iC= 1283 
vC = 14'b0000010011111001; // vC= 1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100011; // iC= 1379 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111010; // iC= 1338 
vC = 14'b0000010010011011; // vC= 1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001110; // iC= 1294 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010001; // iC= 1233 
vC = 14'b0000010010101100; // vC= 1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001011; // iC= 1291 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110010; // iC= 1266 
vC = 14'b0000010100010000; // vC= 1296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000110; // iC= 1286 
vC = 14'b0000010010010110; // vC= 1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111000; // iC= 1336 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010111; // iC= 1303 
vC = 14'b0000010100000111; // vC= 1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110000; // iC= 1328 
vC = 14'b0000010010101111; // vC= 1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110111; // iC= 1335 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011000; // iC= 1240 
vC = 14'b0000010100100001; // vC= 1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101011; // iC= 1195 
vC = 14'b0000010011110110; // vC= 1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110110; // iC= 1270 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111011; // iC= 1211 
vC = 14'b0000010011011000; // vC= 1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101010; // iC= 1258 
vC = 14'b0000010011111011; // vC= 1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100110; // iC= 1254 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100111; // iC= 1255 
vC = 14'b0000010011111001; // vC= 1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000011; // iC= 1283 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110011; // iC= 1267 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101011; // iC= 1259 
vC = 14'b0000010101011010; // vC= 1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000010011101001; // vC= 1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000001; // iC= 1281 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110011; // iC= 1203 
vC = 14'b0000010011010110; // vC= 1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000010; // iC= 1218 
vC = 14'b0000010011010101; // vC= 1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110010; // iC= 1266 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010011; // iC= 1235 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000011; // iC= 1155 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110011; // iC= 1203 
vC = 14'b0000010101110010; // vC= 1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011101; // iC= 1245 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011010; // iC= 1242 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111011; // iC= 1083 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100010; // iC= 1122 
vC = 14'b0000010110001000; // vC= 1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111110; // iC= 1086 
vC = 14'b0000010101000100; // vC= 1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000011; // iC= 1155 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111001; // iC= 1081 
vC = 14'b0000010101001100; // vC= 1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100110; // iC= 1062 
vC = 14'b0000010100100101; // vC= 1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001010; // iC= 1098 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101000; // iC= 1128 
vC = 14'b0000010100100010; // vC= 1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001111; // iC= 1039 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010010; // iC= 1042 
vC = 14'b0000010110011001; // vC= 1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010100; // iC= 1108 
vC = 14'b0000010100111101; // vC= 1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110111; // iC= 1079 
vC = 14'b0000010100110011; // vC= 1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001101; // iC= 1037 
vC = 14'b0000010110000001; // vC= 1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010011; // iC= 1107 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011011; // iC= 1115 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111010; // iC= 1018 
vC = 14'b0000010101011111; // vC= 1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110101; // iC= 1077 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111001; // iC= 1017 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110110; // iC= 1078 
vC = 14'b0000010101101111; // vC= 1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101011; // iC= 1131 
vC = 14'b0000010100110100; // vC= 1332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000011; // iC= 1027 
vC = 14'b0000010110010110; // vC= 1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110100; // iC= 1076 
vC = 14'b0000010110110110; // vC= 1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100011; // iC= 1123 
vC = 14'b0000010101010011; // vC= 1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010110; // iC= 1046 
vC = 14'b0000010101101001; // vC= 1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101101; // iC= 1069 
vC = 14'b0000010111010010; // vC= 1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111011; // iC=  955 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001111; // iC= 1039 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111010; // iC= 1082 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101011; // iC= 1067 
vC = 14'b0000010110111000; // vC= 1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000001; // iC=  961 
vC = 14'b0000010111011000; // vC= 1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111000; // iC=  952 
vC = 14'b0000010110101101; // vC= 1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010011; // iC= 1043 
vC = 14'b0000010110011001; // vC= 1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110001; // iC= 1009 
vC = 14'b0000010111000101; // vC= 1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100110; // iC=  998 
vC = 14'b0000010111001101; // vC= 1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001011; // iC=  907 
vC = 14'b0000010101100001; // vC= 1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011111; // iC=  991 
vC = 14'b0000010101101100; // vC= 1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b0000010110000001; // vC= 1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000111; // iC= 1031 
vC = 14'b0000010101100001; // vC= 1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101111; // iC=  943 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110000; // iC=  880 
vC = 14'b0000010111101011; // vC= 1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011101; // iC=  925 
vC = 14'b0000010101110000; // vC= 1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111111; // iC=  959 
vC = 14'b0000010110011110; // vC= 1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000111; // iC=  967 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b0000010111000100; // vC= 1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011011; // iC=  923 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110101; // iC=  949 
vC = 14'b0000010101111001; // vC= 1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111100; // iC=  892 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110100; // iC=  948 
vC = 14'b0000010110000101; // vC= 1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b0000010111110101; // vC= 1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101101; // iC=  941 
vC = 14'b0000010110101010; // vC= 1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111010; // iC=  954 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110000; // iC=  816 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010001; // iC=  849 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000111; // iC=  839 
vC = 14'b0000010111110001; // vC= 1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101001; // iC=  937 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100001; // iC=  801 
vC = 14'b0000010110111010; // vC= 1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100010; // iC=  930 
vC = 14'b0000010111001010; // vC= 1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010101; // iC=  917 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100000; // iC=  928 
vC = 14'b0000010111010111; // vC= 1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010100; // iC=  916 
vC = 14'b0000010111110111; // vC= 1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100000; // iC=  800 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101110; // iC=  750 
vC = 14'b0000011000001101; // vC= 1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100101; // iC=  869 
vC = 14'b0000010110111111; // vC= 1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010010; // iC=  786 
vC = 14'b0000011000101011; // vC= 1579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110101; // iC=  821 
vC = 14'b0000011001000010; // vC= 1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110001; // iC=  817 
vC = 14'b0000010111010011; // vC= 1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011011; // iC=  795 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001101; // iC=  717 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001000; // iC=  712 
vC = 14'b0000011001000110; // vC= 1606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010000; // iC=  848 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010001; // iC=  721 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011101; // iC=  733 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110001; // iC=  817 
vC = 14'b0000010111110011; // vC= 1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000000; // iC=  832 
vC = 14'b0000011000110110; // vC= 1590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110100; // iC=  692 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000001; // iC=  769 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100110; // iC=  806 
vC = 14'b0000011001001100; // vC= 1612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100101; // iC=  677 
vC = 14'b0000010111111110; // vC= 1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100110; // iC=  742 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101000; // iC=  680 
vC = 14'b0000011000101100; // vC= 1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010001; // iC=  785 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001100; // iC=  780 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000111; // iC=  711 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111011; // iC=  763 
vC = 14'b0000011001100100; // vC= 1636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101010; // iC=  682 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111000; // iC=  632 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110010; // iC=  690 
vC = 14'b0000010111011000; // vC= 1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110111; // iC=  759 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111011; // iC=  635 
vC = 14'b0000010111101011; // vC= 1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000111; // iC=  647 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111110; // iC=  638 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111001; // iC=  697 
vC = 14'b0000010111110111; // vC= 1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000111; // iC=  583 
vC = 14'b0000010111101100; // vC= 1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101100; // iC=  684 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001010; // iC=  714 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111011; // iC=  635 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110000; // iC=  688 
vC = 14'b0000010111111011; // vC= 1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000001; // iC=  641 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111010; // iC=  698 
vC = 14'b0000011001101000; // vC= 1640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100101; // iC=  613 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000011; // iC=  579 
vC = 14'b0000011000010011; // vC= 1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000010; // iC=  578 
vC = 14'b0000010111111110; // vC= 1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111011; // iC=  635 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101001; // iC=  553 
vC = 14'b0000011001101010; // vC= 1642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111101; // iC=  509 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011011; // iC=  603 
vC = 14'b0000011000101101; // vC= 1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100111; // iC=  551 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111101; // iC=  509 
vC = 14'b0000011001110111; // vC= 1655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100000; // iC=  544 
vC = 14'b0000010111110011; // vC= 1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010101; // iC=  597 
vC = 14'b0000011000111101; // vC= 1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000111; // iC=  583 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100011; // iC=  611 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100001; // iC=  481 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010000; // iC=  592 
vC = 14'b0000011001110011; // vC= 1651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111100; // iC=  444 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011001; // iC=  537 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011011; // iC=  539 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001110; // iC=  590 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101000; // iC=  488 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100110; // iC=  486 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110010; // iC=  498 
vC = 14'b0000011000111000; // vC= 1592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011100; // iC=  476 
vC = 14'b0000011010011110; // vC= 1694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011000; // iC=  536 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110011; // iC=  435 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101100; // iC=  492 
vC = 14'b0000011001111110; // vC= 1662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000011; // iC=  387 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011011; // iC=  411 
vC = 14'b0000011000101101; // vC= 1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101110; // iC=  494 
vC = 14'b0000011001111010; // vC= 1658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000100; // iC=  388 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011111; // iC=  351 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101011; // iC=  363 
vC = 14'b0000011010001011; // vC= 1675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101111; // iC=  431 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010101; // iC=  341 
vC = 14'b0000011001010100; // vC= 1620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010101; // iC=  277 
vC = 14'b0000011000010011; // vC= 1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001010; // iC=  266 
vC = 14'b0000011001010110; // vC= 1622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001000; // iC=  392 
vC = 14'b0000011001000000; // vC= 1600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111110; // iC=  254 
vC = 14'b0000011000011001; // vC= 1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010000; // iC=  336 
vC = 14'b0000011000101100; // vC= 1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110100; // iC=  308 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110010; // iC=  242 
vC = 14'b0000011010100000; // vC= 1696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010000; // iC=  208 
vC = 14'b0000011001110111; // vC= 1655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011111; // iC=  287 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011110; // iC=  158 
vC = 14'b0000011001011001; // vC= 1625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100011; // iC=  227 
vC = 14'b0000011010101110; // vC= 1710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101111; // iC=  175 
vC = 14'b0000011010001110; // vC= 1678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000111; // iC=  199 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000001; // iC=  129 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010001; // iC=  209 
vC = 14'b0000011010001110; // vC= 1678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000011; // iC=  131 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101010; // iC=  170 
vC = 14'b0000011001101001; // vC= 1641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000110; // iC=  134 
vC = 14'b0000011001100010; // vC= 1634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000011; // iC=  131 
vC = 14'b0000011001100001; // vC= 1633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001100; // iC=   12 
vC = 14'b0000011000110100; // vC= 1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001110; // iC=   78 
vC = 14'b0000011010000000; // vC= 1664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011010; // iC=  -38 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001101; // iC=   13 
vC = 14'b0000011001000010; // vC= 1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110000; // iC=  -16 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000101; // iC=    5 
vC = 14'b0000011010101110; // vC= 1710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110111; // iC=  -73 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010111; // iC=  -41 
vC = 14'b0000011010100101; // vC= 1701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000101; // iC=  -59 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010011; // iC= -173 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101000; // iC=  -88 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110100; // iC= -140 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001100; // iC= -116 
vC = 14'b0000011010001110; // vC= 1678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001101; // iC= -243 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000010; // iC= -190 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100001; // iC= -287 
vC = 14'b0000011010001010; // vC= 1674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100011; // iC= -349 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101010; // iC= -342 
vC = 14'b0000011001111010; // vC= 1658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010011; // iC= -237 
vC = 14'b0000011010000111; // vC= 1671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100011; // iC= -413 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010000; // iC= -304 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100100; // iC= -348 
vC = 14'b0000011001000010; // vC= 1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110111; // iC= -393 
vC = 14'b0000011010010101; // vC= 1685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001010; // iC= -374 
vC = 14'b0000011010000001; // vC= 1665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011011; // iC= -421 
vC = 14'b0000011001001100; // vC= 1612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010010; // iC= -494 
vC = 14'b0000011001101000; // vC= 1640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011100; // iC= -484 
vC = 14'b0000011010001001; // vC= 1673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001111; // iC= -497 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011111; // iC= -609 
vC = 14'b0000011001011000; // vC= 1624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001111; // iC= -561 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011111; // iC= -609 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110000; // iC= -528 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101011; // iC= -661 
vC = 14'b0000010111100111; // vC= 1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110000; // iC= -592 
vC = 14'b0000011001011101; // vC= 1629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110111; // iC= -713 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010000; // iC= -624 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101011; // iC= -789 
vC = 14'b0000010111110001; // vC= 1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001101; // iC= -819 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000011; // iC= -829 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100011; // iC= -733 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101000; // iC= -728 
vC = 14'b0000010111101011; // vC= 1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110010; // iC= -846 
vC = 14'b0000011000110100; // vC= 1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100101; // iC= -923 
vC = 14'b0000011000110110; // vC= 1590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101111; // iC= -849 
vC = 14'b0000010111111000; // vC= 1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000111; // iC= -953 
vC = 14'b0000011000000001; // vC= 1537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110100; // iC= -844 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001001; // iC= -887 
vC = 14'b0000010110111111; // vC= 1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010000; // iC= -944 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101100; // iC= -980 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101101; // iC= -915 
vC = 14'b0000010111100001; // vC= 1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001101; // iC=-1011 
vC = 14'b0000011000101100; // vC= 1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100011; // iC= -989 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110001; // iC= -975 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010001; // iC=-1071 
vC = 14'b0000010110101000; // vC= 1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100111; // iC=-1049 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010111; // iC=-1129 
vC = 14'b0000010110110010; // vC= 1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110000; // iC=-1104 
vC = 14'b0000010111110001; // vC= 1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101001; // iC=-1047 
vC = 14'b0000010101111101; // vC= 1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010000; // iC=-1072 
vC = 14'b0000011000011001; // vC= 1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110010; // iC=-1230 
vC = 14'b0000010111001101; // vC= 1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011010; // iC=-1254 
vC = 14'b0000010111001110; // vC= 1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100001; // iC=-1119 
vC = 14'b0000010101101100; // vC= 1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011011; // iC=-1189 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010101; // iC=-1195 
vC = 14'b0000010111010110; // vC= 1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110101; // iC=-1163 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000101; // iC=-1275 
vC = 14'b0000010101111110; // vC= 1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001101; // iC=-1267 
vC = 14'b0000010110001101; // vC= 1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101100; // iC=-1364 
vC = 14'b0000010110111111; // vC= 1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000000; // iC=-1280 
vC = 14'b0000010101101111; // vC= 1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100000; // iC=-1376 
vC = 14'b0000010111011000; // vC= 1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110100; // iC=-1292 
vC = 14'b0000010101010100; // vC= 1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001101; // iC=-1267 
vC = 14'b0000010101101101; // vC= 1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100000; // iC=-1376 
vC = 14'b0000010101010010; // vC= 1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101000; // iC=-1368 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000001; // iC=-1407 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011101; // iC=-1443 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b0000010110110111; // vC= 1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001111; // iC=-1457 
vC = 14'b0000010100111100; // vC= 1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001010; // iC=-1462 
vC = 14'b0000010100011001; // vC= 1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b0000010100100100; // vC= 1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000010; // iC=-1534 
vC = 14'b0000010100111101; // vC= 1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001000; // iC=-1464 
vC = 14'b0000010101001100; // vC= 1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111011; // iC=-1413 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001110; // iC=-1458 
vC = 14'b0000010011111000; // vC= 1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b0000010011111101; // vC= 1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b0000010100111000; // vC= 1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010100; // iC=-1516 
vC = 14'b0000010101001000; // vC= 1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101111; // iC=-1553 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b0000010101011010; // vC= 1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b0000010011011010; // vC= 1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b0000010100101001; // vC= 1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111110; // iC=-1538 
vC = 14'b0000010101001100; // vC= 1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b0000010100101010; // vC= 1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b0000010010100111; // vC= 1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b0000010100000110; // vC= 1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b0000010010101011; // vC= 1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010001; // iC=-1583 
vC = 14'b0000010001111101; // vC= 1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011010; // iC=-1702 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110000; // iC=-1680 
vC = 14'b0000010001111010; // vC= 1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b0000010010101110; // vC= 1198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000010011001111; // vC= 1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b0000010011011001; // vC= 1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011010; // iC=-1702 
vC = 14'b0000010001110000; // vC= 1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000010010000011; // vC= 1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b0000010001000000; // vC= 1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110011; // iC=-1741 
vC = 14'b0000010010100010; // vC= 1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010000; // iC=-1648 
vC = 14'b0000010001111000; // vC= 1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000010001010011; // vC= 1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110000; // iC=-1680 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b0000010001111011; // vC= 1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b0000010000101011; // vC= 1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000001111110010; // vC= 1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000001111100001; // vC=  993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b0000001111010101; // vC=  981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000010000001000; // vC= 1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000001111111000; // vC= 1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000010001010011; // vC= 1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000001111100011; // vC=  995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b0000001111001001; // vC=  969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101010; // iC=-1750 
vC = 14'b0000001110100110; // vC=  934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b0000001111110101; // vC= 1013 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111010; // iC=-1670 
vC = 14'b0000001111100001; // vC=  993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111010; // iC=-1670 
vC = 14'b0000001110111011; // vC=  955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000001111010110; // vC=  982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000001110000100; // vC=  900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000001110100111; // vC=  935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b0000001111110100; // vC= 1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101001; // iC=-1815 
vC = 14'b0000001111000010; // vC=  962 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000001111110011; // vC= 1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000001101011100; // vC=  860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000001101011111; // vC=  863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000001101110000; // vC=  880 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b0000001110011100; // vC=  924 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011000; // iC=-1704 
vC = 14'b0000001110010101; // vC=  917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b0000001110010010; // vC=  914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000001110001010; // vC=  906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011101; // iC=-1827 
vC = 14'b0000001101101011; // vC=  875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000001101010101; // vC=  853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b0000001100011001; // vC=  793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100100; // iC=-1820 
vC = 14'b0000001110000011; // vC=  899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000001101100010; // vC=  866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000001100000111; // vC=  775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000001100010101; // vC=  789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b0000001101100001; // vC=  865 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000001100001011; // vC=  779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000001100010101; // vC=  789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000001100100011; // vC=  803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b0000001100110000; // vC=  816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110110; // iC=-1866 
vC = 14'b0000001011111011; // vC=  763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000001011011111; // vC=  735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000001011101100; // vC=  748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b0000001010110111; // vC=  695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b0000001100011110; // vC=  798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000001011011001; // vC=  729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110100; // iC=-1868 
vC = 14'b0000001100111111; // vC=  831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000001011000110; // vC=  710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000001100010110; // vC=  790 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b0000001011100100; // vC=  740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b0000001010001110; // vC=  654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000001011011111; // vC=  735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111100; // iC=-1860 
vC = 14'b0000001011111000; // vC=  760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000001010110111; // vC=  695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001011010110; // vC=  726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111010; // iC=-1862 
vC = 14'b0000001010010011; // vC=  659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000001011001110; // vC=  718 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100101; // iC=-1883 
vC = 14'b0000001011101011; // vC=  747 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000001001010001; // vC=  593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011101; // iC=-1827 
vC = 14'b0000001010100100; // vC=  676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000001010001101; // vC=  653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001100; // iC=-1844 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b0000001001010000; // vC=  592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000001010000100; // vC=  644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000001001110110; // vC=  630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001010; // iC=-1846 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000001001100110; // vC=  614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000001000101100; // vC=  556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000001010000110; // vC=  646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b0000001000000001; // vC=  513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001000011101; // vC=  541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000001001101001; // vC=  617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b0000000111110100; // vC=  500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100000; // iC=-1888 
vC = 14'b0000001000100001; // vC=  545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101101; // iC=-1875 
vC = 14'b0000001001100101; // vC=  613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b0000001001011010; // vC=  602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b0000001000111010; // vC=  570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110010; // iC=-1870 
vC = 14'b0000001000000110; // vC=  518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010110; // iC=-1898 
vC = 14'b0000001000001110; // vC=  526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100110; // iC=-1882 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001000100111; // vC=  551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000000110110100; // vC=  436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011110; // iC=-1890 
vC = 14'b0000000110010100; // vC=  404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100100; // iC=-1884 
vC = 14'b0000001000101101; // vC=  557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000000110011000; // vC=  408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111110; // iC=-1858 
vC = 14'b0000000111011111; // vC=  479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000000110001011; // vC=  395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000000111111101; // vC=  509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000000110010100; // vC=  404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000110100110; // vC=  422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110011; // iC=-1869 
vC = 14'b0000000110010110; // vC=  406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001100; // iC=-1844 
vC = 14'b0000000110100001; // vC=  417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000000101010001; // vC=  337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010010; // iC=-1902 
vC = 14'b0000000111010100; // vC=  468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b0000000110000100; // vC=  388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b0000000101010110; // vC=  342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111000; // iC=-1864 
vC = 14'b0000000100011100; // vC=  284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000000110000111; // vC=  391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001010; // iC=-1846 
vC = 14'b0000000110000111; // vC=  391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000000101110100; // vC=  372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000000100010100; // vC=  276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000000100110010; // vC=  306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000000011101010; // vC=  234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000000100000101; // vC=  261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000000100011001; // vC=  281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011101; // iC=-1827 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011001; // iC=-1895 
vC = 14'b0000000100111101; // vC=  317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000000011110001; // vC=  241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101101; // iC=-1875 
vC = 14'b0000000011111000; // vC=  248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000000011110110; // vC=  246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b0000000101001001; // vC=  329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011000; // iC=-1896 
vC = 14'b0000000100000101; // vC=  261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111000; // iC=-1864 
vC = 14'b0000000100010110; // vC=  278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000000011010011; // vC=  211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b0000000011101101; // vC=  237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b0000000100011010; // vC=  282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011010; // iC=-1894 
vC = 14'b0000000011001100; // vC=  204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000000010010110; // vC=  150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111111; // iC=-1857 
vC = 14'b0000000010111001; // vC=  185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000000100001110; // vC=  270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111110; // iC=-1858 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000000011000000; // vC=  192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000000010111001; // vC=  185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000000011001000; // vC=  200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000000001110110; // vC=  118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101110; // iC=-1874 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100000; // iC=-1760 
vC = 14'b0000000010000011; // vC=  131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111110; // iC=-1858 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000000001011000; // vC=   88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001011; // iC=-1845 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100101; // iC=-1883 
vC = 14'b0000000000101111; // vC=   47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000000001111010; // vC=  122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000000000011011; // vC=   27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111110; // iC=-1858 
vC = 14'b0000000000110100; // vC=   52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101100; // iC=-1876 
vC = 14'b0000000000111000; // vC=   56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000000000101101; // vC=   45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b1111111111101100; // vC=  -20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101101; // iC=-1875 
vC = 14'b0000000000110111; // vC=   55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110000; // iC=-1872 
vC = 14'b0000000000010110; // vC=   22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000000001000; // vC=    8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000000001000111; // vC=   71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b1111111111010011; // vC=  -45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b1111111111101001; // vC=  -23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000000000010010; // vC=   18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b1111111111011101; // vC=  -35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000000000010010; // vC=   18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100000; // iC=-1824 
vC = 14'b0000000000100011; // vC=   35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b1111111110101100; // vC=  -84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b1111111111011111; // vC=  -33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b1111111111000110; // vC=  -58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b1111111111101010; // vC=  -22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b1111111101111101; // vC= -131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b1111111110011111; // vC=  -97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b1111111101011101; // vC= -163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b1111111110110110; // vC=  -74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b1111111110111111; // vC=  -65 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b1111111111000010; // vC=  -62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b1111111110111111; // vC=  -65 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b1111111111010110; // vC=  -42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b1111111110111100; // vC=  -68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b1111111111000110; // vC=  -58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b1111111101001001; // vC= -183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b1111111101111000; // vC= -136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b1111111100011000; // vC= -232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100100; // iC=-1692 
vC = 14'b1111111100010001; // vC= -239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b1111111100100010; // vC= -222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b1111111101110001; // vC= -143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000100; // iC=-1724 
vC = 14'b1111111101111000; // vC= -136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b1111111110001100; // vC= -116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b1111111011101110; // vC= -274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b1111111011110110; // vC= -266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b1111111100101100; // vC= -212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b1111111101001110; // vC= -178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b1111111100111001; // vC= -199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011000; // iC=-1704 
vC = 14'b1111111100011011; // vC= -229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b1111111011010001; // vC= -303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011000; // iC=-1704 
vC = 14'b1111111101011000; // vC= -168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111100; // iC=-1668 
vC = 14'b1111111011100000; // vC= -288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b1111111101000110; // vC= -186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b1111111100111010; // vC= -198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b1111111011001000; // vC= -312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b1111111010100110; // vC= -346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b1111111010100011; // vC= -349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b1111111100000100; // vC= -252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b1111111010011111; // vC= -353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b1111111010100011; // vC= -349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b1111111011100110; // vC= -282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b1111111100011100; // vC= -228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b1111111011010110; // vC= -298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b1111111100000100; // vC= -252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000100; // iC=-1724 
vC = 14'b1111111010100101; // vC= -347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b1111111011110100; // vC= -268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b1111111001110100; // vC= -396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b1111111010010111; // vC= -361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b1111111010001101; // vC= -371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b1111111001101000; // vC= -408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b1111111010000001; // vC= -383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b1111111010010001; // vC= -367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b1111111001111101; // vC= -387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b1111111001001010; // vC= -438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b1111111000101011; // vC= -469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011001; // iC=-1639 
vC = 14'b1111111010110001; // vC= -335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b1111111000110110; // vC= -458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100100; // iC=-1628 
vC = 14'b1111111000110100; // vC= -460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b1111111001111101; // vC= -387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b1111111001011011; // vC= -421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b1111111001110101; // vC= -395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001101; // iC=-1651 
vC = 14'b1111111001010100; // vC= -428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111010; // iC=-1670 
vC = 14'b1111110111110100; // vC= -524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111001; // iC=-1607 
vC = 14'b1111111001100110; // vC= -410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100000; // iC=-1632 
vC = 14'b1111111000010100; // vC= -492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b1111110111101110; // vC= -530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110001; // iC=-1679 
vC = 14'b1111110111100101; // vC= -539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011001; // iC=-1639 
vC = 14'b1111110111010110; // vC= -554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000001; // iC=-1599 
vC = 14'b1111110111110101; // vC= -523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b1111111000111001; // vC= -455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b1111111000110101; // vC= -459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010111; // iC=-1641 
vC = 14'b1111110111011110; // vC= -546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001110; // iC=-1586 
vC = 14'b1111110111101111; // vC= -529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b1111110111001111; // vC= -561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111111; // iC=-1665 
vC = 14'b1111111001000001; // vC= -447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b1111110110011111; // vC= -609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011110; // iC=-1634 
vC = 14'b1111110111010001; // vC= -559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000111; // iC=-1657 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b1111110111011011; // vC= -549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111111; // iC=-1537 
vC = 14'b1111111000100101; // vC= -475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b1111110111011110; // vC= -546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b1111110110100100; // vC= -604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b1111110111010011; // vC= -557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010111; // iC=-1577 
vC = 14'b1111110110001000; // vC= -632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b1111110110110111; // vC= -585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b1111110111001001; // vC= -567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b1111110110010101; // vC= -619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b1111110111100010; // vC= -542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b1111110110000111; // vC= -633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100100; // iC=-1500 
vC = 14'b1111110111010100; // vC= -556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b1111110110100001; // vC= -607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010111; // iC=-1577 
vC = 14'b1111110111000101; // vC= -571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b1111110110110100; // vC= -588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b1111110110100000; // vC= -608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b1111110110001111; // vC= -625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b1111110101001000; // vC= -696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b1111110100011100; // vC= -740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b1111110100010000; // vC= -752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b1111110101001100; // vC= -692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001101; // iC=-1459 
vC = 14'b1111110101010100; // vC= -684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b1111110101101100; // vC= -660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b1111110100011100; // vC= -740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b1111110011101010; // vC= -790 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b1111110101100000; // vC= -672 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001000; // iC=-1464 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000011; // iC=-1533 
vC = 14'b1111110101011011; // vC= -677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b1111110100000100; // vC= -764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011111; // iC=-1441 
vC = 14'b1111110100110000; // vC= -720 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b1111110011110100; // vC= -780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101001; // iC=-1431 
vC = 14'b1111110100100110; // vC= -730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111111; // iC=-1409 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110001; // iC=-1551 
vC = 14'b1111110010111100; // vC= -836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b1111110011001001; // vC= -823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010100; // iC=-1388 
vC = 14'b1111110011111010; // vC= -774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b1111110011001000; // vC= -824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011000; // iC=-1512 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110000; // iC=-1488 
vC = 14'b1111110100001000; // vC= -760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111011; // iC=-1413 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b1111110100011101; // vC= -739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010110; // iC=-1386 
vC = 14'b1111110100001111; // vC= -753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b1111110011101101; // vC= -787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011110; // iC=-1378 
vC = 14'b1111110100010100; // vC= -748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001111; // iC=-1393 
vC = 14'b1111110010100101; // vC= -859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001111; // iC=-1393 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100000; // iC=-1376 
vC = 14'b1111110100001000; // vC= -760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110110; // iC=-1418 
vC = 14'b1111110010011100; // vC= -868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b1111110010000000; // vC= -896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000100; // iC=-1404 
vC = 14'b1111110010111010; // vC= -838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110011; // iC=-1421 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000110; // iC=-1466 
vC = 14'b1111110001100011; // vC= -925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100100; // iC=-1308 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011011; // iC=-1445 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101010; // iC=-1430 
vC = 14'b1111110001010100; // vC= -940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010110; // iC=-1386 
vC = 14'b1111110001110100; // vC= -908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011101; // iC=-1379 
vC = 14'b1111110011000110; // vC= -826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100110; // iC=-1434 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110101; // iC=-1355 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000110; // iC=-1402 
vC = 14'b1111110000101111; // vC= -977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000111; // iC=-1273 
vC = 14'b1111110001111011; // vC= -901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100000; // iC=-1312 
vC = 14'b1111110001001101; // vC= -947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110100; // iC=-1420 
vC = 14'b1111110010000011; // vC= -893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111111; // iC=-1345 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b1111110010000111; // vC= -889 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001100; // iC=-1396 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011101; // iC=-1379 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011100; // iC=-1252 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110001; // iC=-1359 
vC = 14'b1111110001000000; // vC= -960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b1111110001010100; // vC= -940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111001; // iC=-1351 
vC = 14'b1111110000111011; // vC= -965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111010; // iC=-1350 
vC = 14'b1111110000001110; // vC=-1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110100; // iC=-1228 
vC = 14'b1111110000110111; // vC= -969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110100; // iC=-1356 
vC = 14'b1111101111111101; // vC=-1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011000; // iC=-1320 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011011; // iC=-1317 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001010; // iC=-1206 
vC = 14'b1111101111001100; // vC=-1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111101; // iC=-1347 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001011; // iC=-1269 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101100; // iC=-1300 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111101; // iC=-1219 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101100; // iC=-1236 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110001; // iC=-1231 
vC = 14'b1111101110100111; // vC=-1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010110; // iC=-1322 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010111; // iC=-1193 
vC = 14'b1111101110101101; // vC=-1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100100; // iC=-1244 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101001; // iC=-1239 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101101; // iC=-1235 
vC = 14'b1111101111000010; // vC=-1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101100; // iC=-1300 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010010; // iC=-1262 
vC = 14'b1111101110100100; // vC=-1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110110; // iC=-1290 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001000; // iC=-1144 
vC = 14'b1111101111000010; // vC=-1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000100; // iC=-1212 
vC = 14'b1111101110010011; // vC=-1133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110111; // iC=-1161 
vC = 14'b1111101111100011; // vC=-1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111101; // iC=-1155 
vC = 14'b1111110000001101; // vC=-1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100001; // iC=-1119 
vC = 14'b1111101110010001; // vC=-1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000010; // iC=-1150 
vC = 14'b1111101110001001; // vC=-1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010111; // iC=-1129 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111110; // iC=-1154 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001110; // iC=-1202 
vC = 14'b1111101111010101; // vC=-1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000001; // iC=-1151 
vC = 14'b1111101110111111; // vC=-1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111100; // iC=-1092 
vC = 14'b1111101110011001; // vC=-1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000010; // iC=-1086 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001001; // iC=-1079 
vC = 14'b1111101101101000; // vC=-1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111100; // iC=-1092 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011000; // iC=-1128 
vC = 14'b1111101101101100; // vC=-1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010001; // iC=-1071 
vC = 14'b1111101111011010; // vC=-1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010000; // iC=-1072 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100100; // iC=-1052 
vC = 14'b1111101101111011; // vC=-1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001011; // iC=-1077 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101010; // iC=-1110 
vC = 14'b1111101101001101; // vC=-1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001011; // iC=-1141 
vC = 14'b1111101110101111; // vC=-1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010100; // iC=-1132 
vC = 14'b1111101101110110; // vC=-1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110101; // iC=-1099 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101111; // iC=-1105 
vC = 14'b1111101101000000; // vC=-1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111110; // iC=-1090 
vC = 14'b1111101110101111; // vC=-1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110101; // iC=-1035 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111010; // iC=-1094 
vC = 14'b1111101100011111; // vC=-1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001000; // iC=-1080 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000111; // iC=-1017 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100001; // iC= -991 
vC = 14'b1111101100011101; // vC=-1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001111; // iC=-1009 
vC = 14'b1111101101010100; // vC=-1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100101; // iC= -987 
vC = 14'b1111101101110111; // vC=-1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111100; // iC=-1092 
vC = 14'b1111101100110001; // vC=-1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010010; // iC=-1070 
vC = 14'b1111101100101000; // vC=-1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110101; // iC= -971 
vC = 14'b1111101011111101; // vC=-1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100000; // iC=-1056 
vC = 14'b1111101101000011; // vC=-1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110000; // iC=-1104 
vC = 14'b1111101110001010; // vC=-1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111111; // iC=-1025 
vC = 14'b1111101011111111; // vC=-1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100101; // iC=-1051 
vC = 14'b1111101101001100; // vC=-1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111111; // iC= -961 
vC = 14'b1111101101000000; // vC=-1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100011; // iC= -989 
vC = 14'b1111101100011000; // vC=-1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010010; // iC=-1070 
vC = 14'b1111101011101111; // vC=-1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011111; // iC= -929 
vC = 14'b1111101011011000; // vC=-1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100001; // iC=-1055 
vC = 14'b1111101101001010; // vC=-1206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111111; // iC= -961 
vC = 14'b1111101101100000; // vC=-1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110011; // iC=-1037 
vC = 14'b1111101100011110; // vC=-1250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011111; // iC= -929 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111000; // iC= -904 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111100; // iC=-1028 
vC = 14'b1111101100101011; // vC=-1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010001; // iC= -943 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001000; // iC= -888 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100000; // iC= -992 
vC = 14'b1111101100110011; // vC=-1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011111; // iC= -929 
vC = 14'b1111101100101000; // vC=-1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101111; // iC= -977 
vC = 14'b1111101011111001; // vC=-1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110010; // iC= -910 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001011; // iC=-1013 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001100; // iC= -884 
vC = 14'b1111101101001001; // vC=-1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100010; // iC= -926 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100100; // iC= -924 
vC = 14'b1111101100010000; // vC=-1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001101; // iC= -947 
vC = 14'b1111101011100110; // vC=-1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011111; // iC= -929 
vC = 14'b1111101010011100; // vC=-1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110111; // iC= -905 
vC = 14'b1111101100010010; // vC=-1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111000; // iC= -904 
vC = 14'b1111101011111100; // vC=-1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110010; // iC= -846 
vC = 14'b1111101011101010; // vC=-1302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100010; // iC= -862 
vC = 14'b1111101011001001; // vC=-1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010100; // iC= -876 
vC = 14'b1111101011101000; // vC=-1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000011; // iC= -957 
vC = 14'b1111101011101100; // vC=-1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111001; // iC= -903 
vC = 14'b1111101100011101; // vC=-1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000100; // iC= -892 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111110; // iC= -834 
vC = 14'b1111101010001001; // vC=-1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111111; // iC= -833 
vC = 14'b1111101011111101; // vC=-1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110010; // iC= -782 
vC = 14'b1111101011100111; // vC=-1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011111; // iC= -865 
vC = 14'b1111101010110000; // vC=-1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100000; // iC= -800 
vC = 14'b1111101011001000; // vC=-1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011011; // iC= -805 
vC = 14'b1111101100000011; // vC=-1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111001; // iC= -903 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001110; // iC= -754 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011101; // iC= -739 
vC = 14'b1111101011101100; // vC=-1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010010; // iC= -878 
vC = 14'b1111101011110111; // vC=-1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110111; // iC= -777 
vC = 14'b1111101001101001; // vC=-1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000001; // iC= -831 
vC = 14'b1111101011101111; // vC=-1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001011; // iC= -821 
vC = 14'b1111101010111111; // vC=-1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000000; // iC= -768 
vC = 14'b1111101001101110; // vC=-1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100001; // iC= -735 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110111; // iC= -713 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110011; // iC= -845 
vC = 14'b1111101001110010; // vC=-1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011000; // iC= -744 
vC = 14'b1111101001001101; // vC=-1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111110; // iC= -834 
vC = 14'b1111101010110100; // vC=-1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001111; // iC= -753 
vC = 14'b1111101010001101; // vC=-1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000100; // iC= -764 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001000; // iC= -696 
vC = 14'b1111101010111011; // vC=-1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100100; // iC= -668 
vC = 14'b1111101011001010; // vC=-1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110011; // iC= -653 
vC = 14'b1111101010000000; // vC=-1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000010; // iC= -766 
vC = 14'b1111101001011111; // vC=-1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100111; // iC= -665 
vC = 14'b1111101001101000; // vC=-1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100010; // iC= -670 
vC = 14'b1111101011001000; // vC=-1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101010; // iC= -790 
vC = 14'b1111101011001111; // vC=-1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001110; // iC= -754 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010001; // iC= -623 
vC = 14'b1111101001101101; // vC=-1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111010; // iC= -774 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011010; // iC= -742 
vC = 14'b1111101010001111; // vC=-1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011101; // iC= -675 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010100; // iC= -684 
vC = 14'b1111101001100101; // vC=-1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110100; // iC= -716 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101010; // iC= -598 
vC = 14'b1111101000011111; // vC=-1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010000; // iC= -624 
vC = 14'b1111101010011100; // vC=-1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010001; // iC= -687 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100110; // iC= -666 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011111; // iC= -673 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111011; // iC= -709 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000010; // iC= -574 
vC = 14'b1111101010110001; // vC=-1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011011; // iC= -549 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101100; // iC= -660 
vC = 14'b1111101000001111; // vC=-1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001111; // iC= -689 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001001; // iC= -567 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010000; // iC= -624 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100001; // iC= -671 
vC = 14'b1111101010010101; // vC=-1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101010; // iC= -598 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000000; // iC= -576 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111111; // iC= -641 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101100; // iC= -596 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100111; // iC= -601 
vC = 14'b1111101000100111; // vC=-1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111000; // iC= -584 
vC = 14'b1111100111111101; // vC=-1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100101; // iC= -539 
vC = 14'b1111101000111010; // vC=-1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001100; // iC= -628 
vC = 14'b1111101001001001; // vC=-1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101110; // iC= -466 
vC = 14'b1111101000011111; // vC=-1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000001; // iC= -575 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111001; // iC= -583 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110011; // iC= -589 
vC = 14'b1111101000011011; // vC=-1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000101; // iC= -571 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010010; // iC= -558 
vC = 14'b1111100111101000; // vC=-1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011100; // iC= -484 
vC = 14'b1111101001000100; // vC=-1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100001; // iC= -543 
vC = 14'b1111101001100100; // vC=-1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011100; // iC= -548 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010111; // iC= -553 
vC = 14'b1111101000110000; // vC=-1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010000; // iC= -432 
vC = 14'b1111101000100000; // vC=-1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110011; // iC= -525 
vC = 14'b1111101000100001; // vC=-1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100011; // iC= -477 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000011; // iC= -445 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001101; // iC= -435 
vC = 14'b1111100111100111; // vC=-1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110100; // iC= -460 
vC = 14'b1111100111011100; // vC=-1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001101; // iC= -371 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101110; // iC= -466 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000001; // iC= -511 
vC = 14'b1111100111111001; // vC=-1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100000; // iC= -480 
vC = 14'b1111100111100100; // vC=-1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010111; // iC= -425 
vC = 14'b1111100111111000; // vC=-1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111100; // iC= -388 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101100; // iC= -340 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100010; // iC= -414 
vC = 14'b1111100111011111; // vC=-1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111110; // iC= -450 
vC = 14'b1111101001100100; // vC=-1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010101; // iC= -363 
vC = 14'b1111100111110111; // vC=-1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011110; // iC= -418 
vC = 14'b1111100111011111; // vC=-1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110000; // iC= -336 
vC = 14'b1111101000001000; // vC=-1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010100; // iC= -364 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010100; // iC= -236 
vC = 14'b1111100111011011; // vC=-1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001001; // iC= -375 
vC = 14'b1111101001011110; // vC=-1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111011; // iC= -325 
vC = 14'b1111100111101110; // vC=-1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110100; // iC= -268 
vC = 14'b1111100111101110; // vC=-1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111110; // iC= -194 
vC = 14'b1111101000100001; // vC=-1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001001; // iC= -183 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111001; // iC= -263 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110000; // iC= -144 
vC = 14'b1111100111101010; // vC=-1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011010; // iC= -166 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001111; // iC= -113 
vC = 14'b1111100111100000; // vC=-1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000111; // iC= -185 
vC = 14'b1111101000101111; // vC=-1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010011; // iC= -109 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000000; // iC=  -64 
vC = 14'b1111101000011110; // vC=-1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100000; // iC= -160 
vC = 14'b1111101000010100; // vC=-1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101101; // iC= -147 
vC = 14'b1111100111110101; // vC=-1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110101; // iC=  -75 
vC = 14'b1111100111111100; // vC=-1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000101; // iC= -123 
vC = 14'b1111100111100001; // vC=-1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111110; // iC=   -2 
vC = 14'b1111100111000101; // vC=-1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001111; // iC=   15 
vC = 14'b1111100111100110; // vC=-1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100110; // iC=   38 
vC = 14'b1111101001000011; // vC=-1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101101; // iC=  -19 
vC = 14'b1111100111011101; // vC=-1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011100; // iC=  -36 
vC = 14'b1111101001001001; // vC=-1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100001; // iC=   97 
vC = 14'b1111101000111010; // vC=-1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000001; // iC=   65 
vC = 14'b1111101000000100; // vC=-1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010111; // iC=  151 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101110; // iC=  110 
vC = 14'b1111100111011101; // vC=-1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110110; // iC=  182 
vC = 14'b1111100110111110; // vC=-1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010110; // iC=   86 
vC = 14'b1111100110111110; // vC=-1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101111; // iC=  239 
vC = 14'b1111100111010101; // vC=-1579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001100; // iC=  140 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000111; // iC=  199 
vC = 14'b1111101000001001; // vC=-1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010110; // iC=  278 
vC = 14'b1111100111000000; // vC=-1600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001011; // iC=  267 
vC = 14'b1111100111011011; // vC=-1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101011; // iC=  235 
vC = 14'b1111100111011010; // vC=-1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000000; // iC=  256 
vC = 14'b1111101000011110; // vC=-1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001010; // iC=  266 
vC = 14'b1111100111111001; // vC=-1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010100; // iC=  340 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101101; // iC=  429 
vC = 14'b1111100111010011; // vC=-1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001011; // iC=  459 
vC = 14'b1111101001100101; // vC=-1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100110; // iC=  422 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010010; // iC=  466 
vC = 14'b1111100111110011; // vC=-1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001110; // iC=  398 
vC = 14'b1111101000001111; // vC=-1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011101; // iC=  541 
vC = 14'b1111101000001100; // vC=-1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000010; // iC=  450 
vC = 14'b1111101000011001; // vC=-1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110110; // iC=  502 
vC = 14'b1111100111100001; // vC=-1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100110; // iC=  486 
vC = 14'b1111100111011001; // vC=-1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110010; // iC=  626 
vC = 14'b1111101001110000; // vC=-1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110010; // iC=  626 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010111; // iC=  599 
vC = 14'b1111101000000100; // vC=-1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111101; // iC=  637 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010110; // iC=  662 
vC = 14'b1111101000001010; // vC=-1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101011; // iC=  683 
vC = 14'b1111101000110111; // vC=-1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000111; // iC=  711 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001001; // iC=  713 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001111; // iC=  783 
vC = 14'b1111101000011001; // vC=-1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101000; // iC=  744 
vC = 14'b1111101001111100; // vC=-1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110100; // iC=  820 
vC = 14'b1111101000011011; // vC=-1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100110; // iC=  806 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001100; // iC=  844 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010000; // iC=  848 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011001; // iC=  985 
vC = 14'b1111101000001110; // vC=-1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100010; // iC=  930 
vC = 14'b1111101001111110; // vC=-1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000011; // iC= 1027 
vC = 14'b1111101001000110; // vC=-1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011101; // iC= 1053 
vC = 14'b1111101000111110; // vC=-1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b1111101000001111; // vC=-1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001101; // iC= 1037 
vC = 14'b1111101010001001; // vC=-1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000110; // iC= 1030 
vC = 14'b1111101000011111; // vC=-1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110111; // iC= 1079 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001110; // iC= 1102 
vC = 14'b1111101000100000; // vC=-1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101111; // iC= 1071 
vC = 14'b1111101001001111; // vC=-1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000010; // iC= 1154 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000101; // iC= 1221 
vC = 14'b1111101010101111; // vC=-1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111011; // iC= 1083 
vC = 14'b1111101010111111; // vC=-1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110100; // iC= 1140 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101100; // iC= 1132 
vC = 14'b1111101001100101; // vC=-1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101110; // iC= 1198 
vC = 14'b1111101010111101; // vC=-1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010000; // iC= 1232 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101001; // iC= 1257 
vC = 14'b1111101001111111; // vC=-1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000000; // iC= 1344 
vC = 14'b1111101001110110; // vC=-1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110101; // iC= 1269 
vC = 14'b1111101011001101; // vC=-1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011100; // iC= 1372 
vC = 14'b1111101011000101; // vC=-1339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100011; // iC= 1315 
vC = 14'b1111101001011111; // vC=-1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110000; // iC= 1392 
vC = 14'b1111101010110111; // vC=-1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100001; // iC= 1313 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110101; // iC= 1333 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010100; // iC= 1428 
vC = 14'b1111101011110111; // vC=-1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011000; // iC= 1368 
vC = 14'b1111101011010110; // vC=-1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001011; // iC= 1355 
vC = 14'b1111101010110100; // vC=-1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011001; // iC= 1497 
vC = 14'b1111101011111001; // vC=-1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110000; // iC= 1520 
vC = 14'b1111101011001000; // vC=-1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000001; // iC= 1473 
vC = 14'b1111101100100000; // vC=-1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111001; // iC= 1465 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000001; // iC= 1537 
vC = 14'b1111101100010111; // vC=-1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101011; // iC= 1451 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110101; // iC= 1461 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001000; // iC= 1608 
vC = 14'b1111101011100110; // vC=-1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000100; // iC= 1604 
vC = 14'b1111101011010111; // vC=-1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010000; // iC= 1552 
vC = 14'b1111101101000010; // vC=-1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011010; // iC= 1562 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000110; // iC= 1670 
vC = 14'b1111101011100011; // vC=-1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110110; // iC= 1590 
vC = 14'b1111101100101110; // vC=-1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b1111101100000100; // vC=-1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010011; // iC= 1683 
vC = 14'b1111101011101100; // vC=-1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100001; // iC= 1697 
vC = 14'b1111101100110100; // vC=-1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101111; // iC= 1647 
vC = 14'b1111101101001001; // vC=-1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000001; // iC= 1729 
vC = 14'b1111101011111100; // vC=-1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b1111101011110001; // vC=-1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b1111101011111001; // vC=-1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101100; // iC= 1772 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101101; // iC= 1645 
vC = 14'b1111101100001111; // vC=-1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b1111101101110001; // vC=-1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111111; // iC= 1791 
vC = 14'b1111101100000110; // vC=-1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b1111101110000111; // vC=-1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b1111101110100001; // vC=-1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010001; // iC= 1745 
vC = 14'b1111101101111011; // vC=-1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b1111101101101010; // vC=-1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100100; // iC= 1764 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100000; // iC= 1824 
vC = 14'b1111101110110010; // vC=-1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010000; // iC= 1808 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111101110111000; // vC=-1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b1111101101010011; // vC=-1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b1111101111000111; // vC=-1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b1111101110010110; // vC=-1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010010; // iC= 1874 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111101111001001; // vC=-1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101000; // iC= 1832 
vC = 14'b1111101110000011; // vC=-1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111110000001100; // vC=-1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b1111101111000100; // vC=-1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111110000011010; // vC= -998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111110000000101; // vC=-1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b1111101110100110; // vC=-1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b1111101111100100; // vC=-1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111110; // iC= 1982 
vC = 14'b1111110001001111; // vC= -945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b1111110000110110; // vC= -970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101000; // iC= 1832 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111110000010100; // vC=-1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111110000001000; // vC=-1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b1111101111010001; // vC=-1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b1111101111110011; // vC=-1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b1111101111101011; // vC=-1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b1111110001110110; // vC= -906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b1111110000110011; // vC= -973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b1111110001000111; // vC= -953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b1111110001001010; // vC= -950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111110001101101; // vC= -915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110001011100; // vC= -932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111110000110011; // vC= -973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001011; // iC= 1867 
vC = 14'b1111110010011101; // vC= -867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b1111110000101110; // vC= -978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111110010000100; // vC= -892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111110001111111; // vC= -897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110010001011; // vC= -885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111110011011110; // vC= -802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110111; // iC= 1975 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011000; // iC= 1880 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b1111110010010111; // vC= -873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b1111110011111000; // vC= -776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b1111110010011110; // vC= -866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111110001101101; // vC= -915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111101; // iC= 2045 
vC = 14'b1111110011110010; // vC= -782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b1111110010101101; // vC= -851 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b1111110010011001; // vC= -871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b1111110010010001; // vC= -879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111110011010010; // vC= -814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b1111110010101000; // vC= -856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111000; // iC= 2040 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000001; // iC= 2049 
vC = 14'b1111110011100010; // vC= -798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111110011011101; // vC= -803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111110100011001; // vC= -743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100101; // iC= 2021 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000000; // iC= 2048 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111110011011100; // vC= -804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b1111110100010110; // vC= -746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111110100101011; // vC= -725 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111110101110011; // vC= -653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b1111110110000110; // vC= -634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001111; // iC= 2063 
vC = 14'b1111110100100001; // vC= -735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111110100110110; // vC= -714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111110110101011; // vC= -597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111110101111001; // vC= -647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111110110010001; // vC= -623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111110101011110; // vC= -674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111110101001000; // vC= -696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111110100110110; // vC= -714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111110101110111; // vC= -649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111110101010011; // vC= -685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001101; // iC= 2061 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111110111110011; // vC= -525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b1111110111000111; // vC= -569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010110; // iC= 2070 
vC = 14'b1111110111000010; // vC= -574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000001; // iC= 2049 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111111000000001; // vC= -511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111110111001011; // vC= -565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100000; // iC= 2080 
vC = 14'b1111110110110101; // vC= -587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100111; // iC= 2087 
vC = 14'b1111111000011111; // vC= -481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111110111010111; // vC= -553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b1111110111000010; // vC= -574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001010; // iC= 1994 
vC = 14'b1111110110100101; // vC= -603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010101; // iC= 2069 
vC = 14'b1111111000101101; // vC= -467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111110111001010; // vC= -566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111111000001100; // vC= -500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000010; // iC= 2050 
vC = 14'b1111111000101101; // vC= -467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110010; // iC= 2034 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000101010; // iC= 2090 
vC = 14'b1111111000100001; // vC= -479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111111000111111; // vC= -449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000101101; // iC= 2093 
vC = 14'b1111111001011011; // vC= -421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111111000000111; // vC= -505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000001; // iC= 2049 
vC = 14'b1111110111100100; // vC= -540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111111000101101; // vC= -467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111111000011010; // vC= -486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011011; // iC= 2075 
vC = 14'b1111111000010000; // vC= -496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111111001110011; // vC= -397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000111; // iC= 1991 
vC = 14'b1111111000101111; // vC= -465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111111001111000; // vC= -392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b1111111000100001; // vC= -479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000110011; // iC= 2099 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010101; // iC= 2069 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111111010000111; // vC= -377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111111010010100; // vC= -364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111111001111010; // vC= -390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111111010110100; // vC= -332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b1111111011100110; // vC= -282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000101100; // iC= 2092 
vC = 14'b1111111001111010; // vC= -390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010010; // iC= 2066 
vC = 14'b1111111001100011; // vC= -413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101101; // iC= 2029 
vC = 14'b1111111011101001; // vC= -279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b1111111011101101; // vC= -275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011011; // iC= 2075 
vC = 14'b1111111100001110; // vC= -242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111001; // iC= 2041 
vC = 14'b1111111100010111; // vC= -233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111111100000011; // vC= -253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111011010011; // vC= -301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011111; // iC= 2079 
vC = 14'b1111111010101100; // vC= -340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000101; // iC= 2053 
vC = 14'b1111111010100110; // vC= -346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000101111; // iC= 2095 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001010; // iC= 2058 
vC = 14'b1111111011111011; // vC= -261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111111100001001; // vC= -247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101100; // iC= 1964 
vC = 14'b1111111010111011; // vC= -325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111111100101011; // vC= -213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111111011111011; // vC= -261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000101000; // iC= 2088 
vC = 14'b1111111011010101; // vC= -299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111111011010011; // vC= -301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000101; // iC= 2053 
vC = 14'b1111111101110010; // vC= -142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010001; // iC= 2065 
vC = 14'b1111111011111010; // vC= -262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010000; // iC= 2064 
vC = 14'b1111111011110001; // vC= -271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b1111111011101110; // vC= -274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111100010110; // vC= -234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000100; // iC= 2052 
vC = 14'b1111111101011111; // vC= -161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111111110001100; // vC= -116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111111101100010; // vC= -158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111111100100010; // vC= -222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111111110100100; // vC=  -92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111111101100111; // vC= -153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111110; // iC= 1982 
vC = 14'b1111111100110101; // vC= -203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b1111111101001111; // vC= -177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111111100111001; // vC= -199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011000; // iC= 2072 
vC = 14'b1111111111010001; // vC=  -47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101111; // iC= 2031 
vC = 14'b1111111110111011; // vC=  -69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111111110010110; // vC= -106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111110001100; // vC= -116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111111101110001; // vC= -143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b1111111111111100; // vC=   -4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111111111110001; // vC=  -15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111111110100110; // vC=  -90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b1111111110101010; // vC=  -86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b0000000000101001; // vC=   41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b0000000000100100; // vC=   36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010110; // iC= 2070 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111111111011001; // vC=  -39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111111111111001; // vC=   -7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b0000000000011000; // vC=   24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111101; // iC= 2045 
vC = 14'b1111111111111011; // vC=   -5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b0000000000001001; // vC=    9 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b0000000000110101; // vC=   53 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111111; // iC= 2047 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011011; // iC= 2011 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b0000000000111011; // vC=   59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100101; // iC= 2021 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001100; // iC= 2060 
vC = 14'b0000000000010111; // vC=   23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001011; // iC= 2059 
vC = 14'b0000000010001111; // vC=  143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b0000000001111001; // vC=  121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b0000000001110111; // vC=  119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b0000000001000111; // vC=   71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b0000000001111111; // vC=  127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b0000000011001011; // vC=  203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b0000000010000100; // vC=  132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b0000000010010011; // vC=  147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b0000000011001100; // vC=  204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b0000000010111001; // vC=  185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b0000000001111011; // vC=  123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b0000000010110011; // vC=  179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b0000000010110101; // vC=  181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b0000000011110011; // vC=  243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b0000000100101000; // vC=  296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b0000000100000110; // vC=  262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b0000000011001011; // vC=  203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b0000000011100111; // vC=  231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000000011111001; // vC=  249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b0000000010111110; // vC=  190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010010; // iC= 1874 
vC = 14'b0000000100001101; // vC=  269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b0000000100001101; // vC=  269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b0000000011111111; // vC=  255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b0000000100111101; // vC=  317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b0000000100011101; // vC=  285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000000101110100; // vC=  372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001010; // iC= 1994 
vC = 14'b0000000011111101; // vC=  253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b0000000100111111; // vC=  319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111011; // iC= 1851 
vC = 14'b0000000101011001; // vC=  345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b0000000110011000; // vC=  408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b0000000100100000; // vC=  288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b0000000101110110; // vC=  374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110001; // iC= 1841 
vC = 14'b0000000101110011; // vC=  371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b0000000101001010; // vC=  330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000000101100100; // vC=  356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b0000000101000001; // vC=  321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011100; // iC= 1948 
vC = 14'b0000000101001011; // vC=  331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b0000000110100011; // vC=  419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b0000000111010000; // vC=  464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001011; // iC= 1867 
vC = 14'b0000000101100010; // vC=  354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b0000000111010001; // vC=  465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b0000000110101001; // vC=  425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b0000000101101101; // vC=  365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b0000000111101000; // vC=  488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b0000000111111100; // vC=  508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b0000000111101011; // vC=  491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b0000001000000001; // vC=  513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b0000000110111001; // vC=  441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000111; // iC= 1799 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000000111001001; // vC=  457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b0000001000111110; // vC=  574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000101; // iC= 1797 
vC = 14'b0000000111101100; // vC=  492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b0000000111110010; // vC=  498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b0000000111011010; // vC=  474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b0000000111000111; // vC=  455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b0000001000111100; // vC=  572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b0000001001001001; // vC=  585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b0000001000111110; // vC=  574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b0000001001011110; // vC=  606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b0000001001010011; // vC=  595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111110; // iC= 1790 
vC = 14'b0000001001101101; // vC=  621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b0000000111111111; // vC=  511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101001; // iC= 1833 
vC = 14'b0000001000001010; // vC=  522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b0000001001111011; // vC=  635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b0000001000100111; // vC=  551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b0000001010000101; // vC=  645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110101; // iC= 1781 
vC = 14'b0000001001011010; // vC=  602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b0000001010000101; // vC=  645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b0000001010101101; // vC=  685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b0000001010011111; // vC=  671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011111; // iC= 1759 
vC = 14'b0000001001101100; // vC=  620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b0000001011001001; // vC=  713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b0000001001111000; // vC=  632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000001000111001; // vC=  569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b0000001001010010; // vC=  594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b0000001011001001; // vC=  713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b0000001010100101; // vC=  677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101011; // iC= 1707 
vC = 14'b0000001001100101; // vC=  613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101110; // iC= 1838 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000011; // iC= 1795 
vC = 14'b0000001010011001; // vC=  665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b0000001011110010; // vC=  754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b0000001011111011; // vC=  763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100010; // iC= 1826 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000001100001011; // vC=  779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000001010101111; // vC=  687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b0000001010000001; // vC=  641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b0000001011000100; // vC=  708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b0000001010111010; // vC=  698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b0000001100011110; // vC=  798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100011; // iC= 1763 
vC = 14'b0000001100000101; // vC=  773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b0000001100101010; // vC=  810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b0000001011001111; // vC=  719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b0000001011101001; // vC=  745 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000001011000000; // vC=  704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000001; // iC= 1665 
vC = 14'b0000001100000011; // vC=  771 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100101; // iC= 1765 
vC = 14'b0000001101001100; // vC=  844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b0000001100101110; // vC=  814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100111; // iC= 1703 
vC = 14'b0000001100101111; // vC=  815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b0000001011111001; // vC=  761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010001; // iC= 1745 
vC = 14'b0000001011100101; // vC=  741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010011; // iC= 1683 
vC = 14'b0000001100111010; // vC=  826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b0000001100001010; // vC=  778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111110; // iC= 1662 
vC = 14'b0000001100000011; // vC=  771 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b0000001101100010; // vC=  866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b0000001100001110; // vC=  782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101010; // iC= 1642 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000000; // iC= 1664 
vC = 14'b0000001100011100; // vC=  796 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b0000001110010000; // vC=  912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b0000001101001001; // vC=  841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b0000001110011101; // vC=  925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100011; // iC= 1571 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b0000001101000111; // vC=  839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100110; // iC= 1702 
vC = 14'b0000001101111001; // vC=  889 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b0000001110000000; // vC=  896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011001; // iC= 1625 
vC = 14'b0000001110001001; // vC=  905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b0000001110100101; // vC=  933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110101; // iC= 1653 
vC = 14'b0000001101010111; // vC=  855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101001; // iC= 1641 
vC = 14'b0000001110011111; // vC=  927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001011; // iC= 1675 
vC = 14'b0000001101111000; // vC=  888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101011; // iC= 1579 
vC = 14'b0000001111100110; // vC=  998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001100; // iC= 1612 
vC = 14'b0000001110001111; // vC=  911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b0000001110010111; // vC=  919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110110; // iC= 1590 
vC = 14'b0000001110111000; // vC=  952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000100; // iC= 1604 
vC = 14'b0000001110000101; // vC=  901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101000; // iC= 1640 
vC = 14'b0000001110010100; // vC=  916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111010; // iC= 1658 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101010; // iC= 1514 
vC = 14'b0000001111111100; // vC= 1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000001; // iC= 1601 
vC = 14'b0000001101111011; // vC=  891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110001; // iC= 1649 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b0000001110101101; // vC=  941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b0000001110000010; // vC=  898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b0000001110011001; // vC=  921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011101; // iC= 1629 
vC = 14'b0000010000001010; // vC= 1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010100; // iC= 1492 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100100; // iC= 1572 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000001111101011; // vC= 1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010111; // iC= 1495 
vC = 14'b0000001110100011; // vC=  931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000101; // iC= 1605 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001010; // iC= 1482 
vC = 14'b0000010000111101; // vC= 1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010001; // iC= 1553 
vC = 14'b0000001111010011; // vC=  979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010100; // iC= 1492 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001011; // iC= 1483 
vC = 14'b0000010000011010; // vC= 1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010101; // iC= 1493 
vC = 14'b0000001111100001; // vC=  993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011111; // iC= 1567 
vC = 14'b0000010000000001; // vC= 1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101110; // iC= 1582 
vC = 14'b0000001111010110; // vC=  982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100011; // iC= 1571 
vC = 14'b0000010000001110; // vC= 1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101101; // iC= 1453 
vC = 14'b0000010001010110; // vC= 1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100011; // iC= 1443 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100101; // iC= 1573 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010111; // iC= 1431 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110010; // iC= 1522 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010001; // iC= 1489 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101100; // iC= 1516 
vC = 14'b0000010001001000; // vC= 1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101001; // iC= 1513 
vC = 14'b0000010000110110; // vC= 1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110001; // iC= 1393 
vC = 14'b0000010010011001; // vC= 1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110011; // iC= 1459 
vC = 14'b0000010010001100; // vC= 1164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001001; // iC= 1481 
vC = 14'b0000010001101000; // vC= 1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111001; // iC= 1465 
vC = 14'b0000010000111101; // vC= 1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010111; // iC= 1431 
vC = 14'b0000010010011011; // vC= 1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111010; // iC= 1466 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101100; // iC= 1516 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001010; // iC= 1354 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100001; // iC= 1441 
vC = 14'b0000010001011110; // vC= 1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011111; // iC= 1375 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101001; // iC= 1385 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001111; // iC= 1423 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000010; // iC= 1474 
vC = 14'b0000010001101000; // vC= 1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000000; // iC= 1344 
vC = 14'b0000010001001000; // vC= 1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000100; // iC= 1412 
vC = 14'b0000010010000010; // vC= 1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100101; // iC= 1445 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111111; // iC= 1471 
vC = 14'b0000010011100100; // vC= 1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111001; // iC= 1337 
vC = 14'b0000010001110110; // vC= 1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000110; // iC= 1350 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100011; // iC= 1379 
vC = 14'b0000010001111101; // vC= 1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111010; // iC= 1402 
vC = 14'b0000010001101110; // vC= 1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001010; // iC= 1290 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110100; // iC= 1396 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100010; // iC= 1378 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110000; // iC= 1328 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100100; // iC= 1380 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000001; // iC= 1345 
vC = 14'b0000010011100110; // vC= 1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100011; // iC= 1315 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001000; // iC= 1416 
vC = 14'b0000010011101000; // vC= 1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011100; // iC= 1372 
vC = 14'b0000010011011100; // vC= 1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111011; // iC= 1339 
vC = 14'b0000010010000101; // vC= 1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101101; // iC= 1389 
vC = 14'b0000010011100110; // vC= 1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100100; // iC= 1252 
vC = 14'b0000010011100101; // vC= 1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000010; // iC= 1282 
vC = 14'b0000010011101111; // vC= 1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010000; // iC= 1296 
vC = 14'b0000010011110100; // vC= 1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011100; // iC= 1244 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010001; // iC= 1361 
vC = 14'b0000010100011000; // vC= 1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100000; // iC= 1248 
vC = 14'b0000010011101110; // vC= 1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110011; // iC= 1331 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111011; // iC= 1211 
vC = 14'b0000010011101001; // vC= 1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000101; // iC= 1285 
vC = 14'b0000010011001110; // vC= 1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111100; // iC= 1276 
vC = 14'b0000010011111100; // vC= 1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100100; // iC= 1252 
vC = 14'b0000010100000110; // vC= 1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111111; // iC= 1215 
vC = 14'b0000010101010011; // vC= 1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101101; // iC= 1197 
vC = 14'b0000010101010111; // vC= 1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010101; // iC= 1237 
vC = 14'b0000010100110011; // vC= 1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100100; // iC= 1252 
vC = 14'b0000010011011001; // vC= 1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111010; // iC= 1274 
vC = 14'b0000010011110111; // vC= 1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100100; // iC= 1188 
vC = 14'b0000010011100001; // vC= 1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110110; // iC= 1206 
vC = 14'b0000010101011100; // vC= 1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101110; // iC= 1198 
vC = 14'b0000010011100111; // vC= 1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100011; // iC= 1251 
vC = 14'b0000010101101111; // vC= 1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100101; // iC= 1253 
vC = 14'b0000010100110001; // vC= 1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011001; // iC= 1241 
vC = 14'b0000010101011111; // vC= 1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000010100101011; // vC= 1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110000; // iC= 1136 
vC = 14'b0000010100111001; // vC= 1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010110; // iC= 1174 
vC = 14'b0000010100010100; // vC= 1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010101; // iC= 1237 
vC = 14'b0000010110001010; // vC= 1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101111; // iC= 1199 
vC = 14'b0000010100111010; // vC= 1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011101; // iC= 1117 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010110; // iC= 1174 
vC = 14'b0000010110001100; // vC= 1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100101; // iC= 1125 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010101; // iC= 1173 
vC = 14'b0000010101110111; // vC= 1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100010; // iC= 1122 
vC = 14'b0000010110010000; // vC= 1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111100; // iC= 1084 
vC = 14'b0000010110100101; // vC= 1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110100; // iC= 1140 
vC = 14'b0000010101111110; // vC= 1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001011; // iC= 1163 
vC = 14'b0000010100111010; // vC= 1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000111; // iC= 1159 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110100; // iC= 1140 
vC = 14'b0000010100101100; // vC= 1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110010; // iC= 1138 
vC = 14'b0000010110011011; // vC= 1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010111; // iC= 1111 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010011; // iC= 1043 
vC = 14'b0000010110010100; // vC= 1428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011010; // iC= 1114 
vC = 14'b0000010110011011; // vC= 1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011010; // iC= 1114 
vC = 14'b0000010101100010; // vC= 1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010001; // iC= 1105 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100001; // iC= 1121 
vC = 14'b0000010111000000; // vC= 1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010101; // iC= 1173 
vC = 14'b0000010101000110; // vC= 1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000110; // iC= 1030 
vC = 14'b0000010111001111; // vC= 1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001100; // iC= 1036 
vC = 14'b0000010101101001; // vC= 1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010000; // iC= 1104 
vC = 14'b0000010111001111; // vC= 1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010000; // iC= 1040 
vC = 14'b0000010101111010; // vC= 1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001010; // iC= 1034 
vC = 14'b0000010101100110; // vC= 1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100000; // iC= 1120 
vC = 14'b0000010110110000; // vC= 1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001010; // iC= 1034 
vC = 14'b0000010101111001; // vC= 1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010011; // iC= 1107 
vC = 14'b0000010111010110; // vC= 1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101101; // iC= 1005 
vC = 14'b0000010110100010; // vC= 1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001100; // iC= 1100 
vC = 14'b0000010101001100; // vC= 1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111000; // iC= 1016 
vC = 14'b0000010110110010; // vC= 1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010011; // iC= 1107 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100010; // iC=  994 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110101; // iC= 1077 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100101; // iC=  933 
vC = 14'b0000010110111001; // vC= 1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011010; // iC=  986 
vC = 14'b0000010110010011; // vC= 1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011101; // iC= 1053 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101001; // iC= 1001 
vC = 14'b0000010111101011; // vC= 1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010101; // iC=  917 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000110; // iC=  966 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000000; // iC=  960 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111000; // iC=  952 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101001; // iC= 1001 
vC = 14'b0000010111111101; // vC= 1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110111; // iC=  951 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000101; // iC= 1029 
vC = 14'b0000010111100111; // vC= 1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000111; // iC= 1031 
vC = 14'b0000010110001100; // vC= 1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111111; // iC=  895 
vC = 14'b0000010111011011; // vC= 1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110001; // iC=  881 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100101; // iC=  933 
vC = 14'b0000010110001111; // vC= 1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100100; // iC=  932 
vC = 14'b0000010110100000; // vC= 1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100110; // iC=  934 
vC = 14'b0000011000011001; // vC= 1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111100; // iC=  956 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001101; // iC=  973 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010110; // iC=  854 
vC = 14'b0000010111001110; // vC= 1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001011; // iC=  971 
vC = 14'b0000011000101100; // vC= 1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101000; // iC=  936 
vC = 14'b0000011000110101; // vC= 1589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110001; // iC=  945 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010110; // iC=  854 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100000; // iC=  800 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001111; // iC=  847 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110100; // iC=  948 
vC = 14'b0000010111001110; // vC= 1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011111; // iC=  927 
vC = 14'b0000011000111110; // vC= 1598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001010; // iC=  842 
vC = 14'b0000010111010000; // vC= 1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010000; // iC=  784 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111101; // iC=  893 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011000; // iC=  920 
vC = 14'b0000011000101010; // vC= 1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100100; // iC=  868 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010100; // iC=  852 
vC = 14'b0000010111001001; // vC= 1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011000; // iC=  856 
vC = 14'b0000010111010111; // vC= 1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110100; // iC=  820 
vC = 14'b0000010111000000; // vC= 1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101101; // iC=  877 
vC = 14'b0000011000111101; // vC= 1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101011; // iC=  875 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000100; // iC=  772 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010001; // iC=  849 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000101; // iC=  837 
vC = 14'b0000010111010101; // vC= 1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001111; // iC=  783 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111100; // iC=  700 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100000; // iC=  800 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111001; // iC=  825 
vC = 14'b0000010111100001; // vC= 1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101000; // iC=  808 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100111; // iC=  679 
vC = 14'b0000010111011000; // vC= 1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011110; // iC=  670 
vC = 14'b0000010111100010; // vC= 1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011000; // iC=  664 
vC = 14'b0000011001100011; // vC= 1635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000001; // iC=  705 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010010; // iC=  722 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111000; // iC=  696 
vC = 14'b0000011001111001; // vC= 1657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110110; // iC=  758 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111000; // iC=  632 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100000; // iC=  672 
vC = 14'b0000010111100010; // vC= 1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001101; // iC=  781 
vC = 14'b0000011000101101; // vC= 1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111100; // iC=  764 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101100; // iC=  748 
vC = 14'b0000011001110010; // vC= 1650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001110; // iC=  718 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100100; // iC=  612 
vC = 14'b0000011001110011; // vC= 1651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011010; // iC=  666 
vC = 14'b0000011001111011; // vC= 1659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010011; // iC=  659 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000101; // iC=  581 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100001; // iC=  609 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010010; // iC=  722 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000111; // iC=  711 
vC = 14'b0000011001110001; // vC= 1649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100011; // iC=  675 
vC = 14'b0000011001010001; // vC= 1617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001000; // iC=  648 
vC = 14'b0000011010000101; // vC= 1669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101001; // iC=  553 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110000; // iC=  688 
vC = 14'b0000011001110111; // vC= 1655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011110; // iC=  670 
vC = 14'b0000010111111011; // vC= 1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101111; // iC=  687 
vC = 14'b0000011001010100; // vC= 1620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010100; // iC=  660 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101001; // iC=  617 
vC = 14'b0000011010011101; // vC= 1693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100011; // iC=  611 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000101; // iC=  517 
vC = 14'b0000011010100011; // vC= 1699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011000; // iC=  536 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010101; // iC=  597 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001001; // iC=  521 
vC = 14'b0000011000111000; // vC= 1592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111010; // iC=  634 
vC = 14'b0000011010100111; // vC= 1703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101110; // iC=  558 
vC = 14'b0000011010001010; // vC= 1674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101000; // iC=  552 
vC = 14'b0000011001000011; // vC= 1603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001101; // iC=  525 
vC = 14'b0000011000110010; // vC= 1586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000000; // iC=  576 
vC = 14'b0000011010110000; // vC= 1712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001110; // iC=  462 
vC = 14'b0000011001101010; // vC= 1642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000100; // iC=  452 
vC = 14'b0000011001010100; // vC= 1620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111000; // iC=  504 
vC = 14'b0000011010011101; // vC= 1693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101000; // iC=  552 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001000; // iC=  584 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111011; // iC=  443 
vC = 14'b0000011001101001; // vC= 1641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110110; // iC=  438 
vC = 14'b0000011010011111; // vC= 1695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000001; // iC=  449 
vC = 14'b0000011010000100; // vC= 1668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100011; // iC=  547 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100111; // iC=  423 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101100; // iC=  492 
vC = 14'b0000011010000011; // vC= 1667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111001; // iC=  441 
vC = 14'b0000011001011101; // vC= 1629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010011; // iC=  467 
vC = 14'b0000011001110111; // vC= 1655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111000; // iC=  504 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011101; // iC=  349 
vC = 14'b0000011010011011; // vC= 1691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110111; // iC=  375 
vC = 14'b0000011010100010; // vC= 1698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010011; // iC=  339 
vC = 14'b0000011010111010; // vC= 1722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010001; // iC=  337 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000111; // iC=  391 
vC = 14'b0000011010001000; // vC= 1672 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111101; // iC=  381 
vC = 14'b0000011010001010; // vC= 1674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000010; // iC=  386 
vC = 14'b0000011001011001; // vC= 1625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100111; // iC=  295 
vC = 14'b0000011010110101; // vC= 1717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000100; // iC=  260 
vC = 14'b0000011001100101; // vC= 1637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100110; // iC=  294 
vC = 14'b0000011010011111; // vC= 1695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110010; // iC=  370 
vC = 14'b0000011001110110; // vC= 1654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000111; // iC=  327 
vC = 14'b0000011010010000; // vC= 1680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001100; // iC=  332 
vC = 14'b0000011001011101; // vC= 1629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111100; // iC=  188 
vC = 14'b0000011000111000; // vC= 1592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100101; // iC=  293 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100101; // iC=  229 
vC = 14'b0000011010011010; // vC= 1690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011101; // iC=  221 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110001; // iC=  241 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000101; // iC=  133 
vC = 14'b0000011010100000; // vC= 1696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101010; // iC=  106 
vC = 14'b0000011001000110; // vC= 1606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011101; // iC=  157 
vC = 14'b0000011010110001; // vC= 1713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011100; // iC=  156 
vC = 14'b0000011010010110; // vC= 1686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000111; // iC=  199 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111011; // iC=  123 
vC = 14'b0000011001010100; // vC= 1620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011110; // iC=   30 
vC = 14'b0000011001110011; // vC= 1651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011110; // iC=   30 
vC = 14'b0000011011000110; // vC= 1734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101010; // iC=  -22 
vC = 14'b0000011000111101; // vC= 1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011110; // iC=  -34 
vC = 14'b0000011011000011; // vC= 1731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100100; // iC=   36 
vC = 14'b0000011001011110; // vC= 1630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111001; // iC=  -71 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000011; // iC=  -61 
vC = 14'b0000011010011101; // vC= 1693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011101; // iC=  -35 
vC = 14'b0000011010001111; // vC= 1679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000101; // iC=  -59 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100010; // iC=  -94 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011110; // iC= -162 
vC = 14'b0000011010110010; // vC= 1714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110000; // iC=  -80 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000100; // iC= -124 
vC = 14'b0000011001111110; // vC= 1662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101110; // iC= -210 
vC = 14'b0000011001010111; // vC= 1623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011111; // iC= -161 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001111; // iC= -177 
vC = 14'b0000011010010000; // vC= 1680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111000; // iC= -264 
vC = 14'b0000011010010001; // vC= 1681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100100; // iC= -220 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011110; // iC= -290 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111111; // iC= -321 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100100; // iC= -348 
vC = 14'b0000011000101000; // vC= 1576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011010; // iC= -358 
vC = 14'b0000011000101100; // vC= 1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011101; // iC= -419 
vC = 14'b0000011001000000; // vC= 1600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000000; // iC= -320 
vC = 14'b0000011010001100; // vC= 1676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001010; // iC= -374 
vC = 14'b0000011000101111; // vC= 1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010100; // iC= -428 
vC = 14'b0000011001101100; // vC= 1644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011111; // iC= -481 
vC = 14'b0000011000110010; // vC= 1586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000011; // iC= -445 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000001; // iC= -511 
vC = 14'b0000011010100001; // vC= 1697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101101; // iC= -595 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011001; // iC= -487 
vC = 14'b0000011001011001; // vC= 1625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111000; // iC= -520 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001111; // iC= -561 
vC = 14'b0000011010000111; // vC= 1671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101101; // iC= -595 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110001; // iC= -591 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011011; // iC= -741 
vC = 14'b0000011001100010; // vC= 1634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001110; // iC= -626 
vC = 14'b0000011010000011; // vC= 1667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010100; // iC= -684 
vC = 14'b0000011001110110; // vC= 1654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010010; // iC= -686 
vC = 14'b0000011001110011; // vC= 1651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110001; // iC= -783 
vC = 14'b0000011001000010; // vC= 1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111011; // iC= -837 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000101; // iC= -827 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111011; // iC= -773 
vC = 14'b0000011001100010; // vC= 1634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101001; // iC= -791 
vC = 14'b0000010111011101; // vC= 1501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001000; // iC= -824 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010101; // iC= -875 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110110; // iC= -842 
vC = 14'b0000010111001000; // vC= 1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110000; // iC= -912 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110011; // iC= -909 
vC = 14'b0000010111011110; // vC= 1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111001; // iC=-1031 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011001; // iC= -999 
vC = 14'b0000010111110111; // vC= 1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010011; // iC= -941 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111110; // iC= -962 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000001; // iC=-1023 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110110; // iC=-1098 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100010; // iC=-1118 
vC = 14'b0000010111110100; // vC= 1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010101; // iC=-1067 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011101; // iC=-1059 
vC = 14'b0000010111110100; // vC= 1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001101; // iC=-1139 
vC = 14'b0000010110010111; // vC= 1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011111; // iC=-1185 
vC = 14'b0000011000101010; // vC= 1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101110; // iC=-1106 
vC = 14'b0000010111100110; // vC= 1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101100; // iC=-1108 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100101; // iC=-1179 
vC = 14'b0000010110101000; // vC= 1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110001; // iC=-1231 
vC = 14'b0000010111111111; // vC= 1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001001; // iC=-1271 
vC = 14'b0000010111000100; // vC= 1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100100; // iC=-1180 
vC = 14'b0000010110110110; // vC= 1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011110; // iC=-1186 
vC = 14'b0000010110001111; // vC= 1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000001; // iC=-1215 
vC = 14'b0000010111001010; // vC= 1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000011; // iC=-1213 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011100; // iC=-1252 
vC = 14'b0000010111000011; // vC= 1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100110; // iC=-1242 
vC = 14'b0000010111000011; // vC= 1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010011; // iC=-1325 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b0000010101010010; // vC= 1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001100; // iC=-1396 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011101; // iC=-1443 
vC = 14'b0000010110000100; // vC= 1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000111; // iC=-1401 
vC = 14'b0000010101101010; // vC= 1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101111; // iC=-1361 
vC = 14'b0000010101111001; // vC= 1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011011; // iC=-1381 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111011; // iC=-1413 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001110; // iC=-1458 
vC = 14'b0000010100011111; // vC= 1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b0000010110011010; // vC= 1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b0000010100100010; // vC= 1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b0000010100100100; // vC= 1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b0000010101111001; // vC= 1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b0000010101001011; // vC= 1355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b0000010101011100; // vC= 1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b0000010100110011; // vC= 1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b0000010011010111; // vC= 1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b0000010100111110; // vC= 1342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b0000010100011111; // vC= 1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b0000010011100000; // vC= 1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110111; // iC=-1673 
vC = 14'b0000010100111111; // vC= 1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b0000010010110011; // vC= 1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b0000010100001101; // vC= 1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b0000010010110011; // vC= 1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b0000010010110001; // vC= 1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010011; // iC=-1581 
vC = 14'b0000010011001111; // vC= 1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000010010010101; // vC= 1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b0000010010000001; // vC= 1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b0000010011000100; // vC= 1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000010010011011; // vC= 1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001101; // iC=-1651 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000010010110011; // vC= 1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b0000010011000001; // vC= 1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011000; // iC=-1704 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b0000010010110111; // vC= 1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000010011001101; // vC= 1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000010001000011; // vC= 1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000010010001111; // vC= 1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000010000100101; // vC= 1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b0000010000011001; // vC= 1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000010000111100; // vC= 1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b0000010001101011; // vC= 1131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000010001011010; // vC= 1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b0000010000111000; // vC= 1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b0000001110111010; // vC=  954 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b0000001111010100; // vC=  980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001111111000; // vC= 1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000001110101000; // vC=  936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000001111101101; // vC= 1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110001; // iC=-1679 
vC = 14'b0000001111100011; // vC=  995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000001111111000; // vC= 1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b0000001110010101; // vC=  917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000001111111100; // vC= 1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000001110011000; // vC=  920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111011; // iC=-1797 
vC = 14'b0000001111010001; // vC=  977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b0000001110011101; // vC=  925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000001101100101; // vC=  869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000001101100010; // vC=  866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001011; // iC=-1845 
vC = 14'b0000001111011111; // vC=  991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011010; // iC=-1830 
vC = 14'b0000001101111101; // vC=  893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000001101100000; // vC=  864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000001101010010; // vC=  850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000001101101010; // vC=  874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011101; // iC=-1699 
vC = 14'b0000001110110111; // vC=  951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000001110101110; // vC=  942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000001110000100; // vC=  900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000001110100110; // vC=  934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001100011000; // vC=  792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b0000001101110111; // vC=  887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000001101110111; // vC=  887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000001100110000; // vC=  816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000010; // iC=-1854 
vC = 14'b0000001110000110; // vC=  902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001100000110; // vC=  774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000001011011010; // vC=  730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000001011011100; // vC=  732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000001100110101; // vC=  821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000001010111111; // vC=  703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000001100011000; // vC=  792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000001011000010; // vC=  706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000001100001010; // vC=  778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000001010010101; // vC=  661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000001010111100; // vC=  700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000001010111001; // vC=  697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101101; // iC=-1875 
vC = 14'b0000001010100100; // vC=  676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011100; // iC=-1892 
vC = 14'b0000001011010101; // vC=  725 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000001011001101; // vC=  717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100101; // iC=-1883 
vC = 14'b0000001001110000; // vC=  624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000001001111110; // vC=  638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b0000001011100111; // vC=  743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001110; // iC=-1842 
vC = 14'b0000001011010110; // vC=  726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000001010000110; // vC=  646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100000; // iC=-1888 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000001001110110; // vC=  630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b0000001001100010; // vC=  610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000001010001101; // vC=  653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000001000111001; // vC=  569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000001010111010; // vC=  698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000001001101001; // vC=  617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b0000001001111001; // vC=  633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001111; // iC=-1841 
vC = 14'b0000001001010001; // vC=  593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011101; // iC=-1827 
vC = 14'b0000001001011110; // vC=  606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011011; // iC=-1893 
vC = 14'b0000001010001010; // vC=  650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001110; // iC=-1842 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b0000000111101101; // vC=  493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010001; // iC=-1903 
vC = 14'b0000000111011011; // vC=  475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b0000001000111001; // vC=  569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000000111100001; // vC=  481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000000111011101; // vC=  477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010001011; // iC=-1909 
vC = 14'b0000000111101011; // vC=  491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011111; // iC=-1889 
vC = 14'b0000000111001001; // vC=  457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000000111111010; // vC=  506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000111011101; // vC=  477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000001000101100; // vC=  556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000000111100010; // vC=  482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011111; // iC=-1889 
vC = 14'b0000000110001111; // vC=  399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000000111000101; // vC=  453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001000100100; // vC=  548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110011; // iC=-1869 
vC = 14'b0000001000011101; // vC=  541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111011; // iC=-1861 
vC = 14'b0000000110110100; // vC=  436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101011; // iC=-1877 
vC = 14'b0000000111101100; // vC=  492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010100; // iC=-1900 
vC = 14'b0000000110011011; // vC=  411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111011; // iC=-1861 
vC = 14'b0000000110010000; // vC=  400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000000111000100; // vC=  452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000101011101; // vC=  349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000000110101110; // vC=  430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b0000000110011110; // vC=  414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000000101100100; // vC=  356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000000110110100; // vC=  436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000000110101001; // vC=  425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010001111; // iC=-1905 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110011; // iC=-1869 
vC = 14'b0000000101111101; // vC=  381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000000101100100; // vC=  356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b0000000100101101; // vC=  301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010001101; // iC=-1907 
vC = 14'b0000000101101011; // vC=  363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b0000000110010011; // vC=  403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010001000; // iC=-1912 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100111; // iC=-1881 
vC = 14'b0000000100001001; // vC=  265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000000100111011; // vC=  315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b0000000100010010; // vC=  274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101000; // iC=-1880 
vC = 14'b0000000100111100; // vC=  316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b0000000101011100; // vC=  348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011010; // iC=-1894 
vC = 14'b0000000011001111; // vC=  207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000000; // iC=-1792 
vC = 14'b0000000011000110; // vC=  198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100000; // iC=-1760 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000000100110010; // vC=  306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000000011101000; // vC=  232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010111; // iC=-1897 
vC = 14'b0000000101000001; // vC=  321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010100; // iC=-1836 
vC = 14'b0000000100110111; // vC=  311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011110; // iC=-1890 
vC = 14'b0000000011000111; // vC=  199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100000; // iC=-1888 
vC = 14'b0000000011111111; // vC=  255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000000011100110; // vC=  230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000011; // iC=-1853 
vC = 14'b0000000011111010; // vC=  250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b0000000010010010; // vC=  146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010110; // iC=-1898 
vC = 14'b0000000011001011; // vC=  203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100110; // iC=-1882 
vC = 14'b0000000010101000; // vC=  168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000011010010; // vC=  210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000000001011101; // vC=   93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b0000000001010000; // vC=   80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101101; // iC=-1875 
vC = 14'b0000000011000011; // vC=  195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000000001000111; // vC=   71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000000001011010; // vC=   90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000000000110100; // vC=   52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000000000101010; // vC=   42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000000010000011; // vC=  131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000000001010100; // vC=   84 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110010; // iC=-1870 
vC = 14'b0000000000011010; // vC=   26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110010; // iC=-1806 
vC = 14'b1111111111101100; // vC=  -20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000000001101011; // vC=  107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100000; // iC=-1824 
vC = 14'b0000000000011101; // vC=   29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b1111111111000011; // vC=  -61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b1111111111000110; // vC=  -58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b1111111111001000; // vC=  -56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000011; // iC=-1853 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110000; // iC=-1872 
vC = 14'b0000000000011010; // vC=   26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b1111111111110000; // vC=  -16 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b1111111110101011; // vC=  -85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000000000101101; // vC=   45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b1111111110101110; // vC=  -82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b0000000000000110; // vC=    6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b1111111111000111; // vC=  -57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b1111111111010101; // vC=  -43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b1111111111000101; // vC=  -59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b1111111111100111; // vC=  -25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b1111111111101000; // vC=  -24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010100; // iC=-1836 
vC = 14'b1111111111101110; // vC=  -18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b1111111110110001; // vC=  -79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010011; // iC=-1837 
vC = 14'b1111111111000010; // vC=  -62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b1111111110010111; // vC= -105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b1111111101101011; // vC= -149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b1111111101010001; // vC= -175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b1111111110110001; // vC=  -79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b1111111101110100; // vC= -140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b1111111110100101; // vC=  -91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b1111111110001101; // vC= -115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b1111111100111001; // vC= -199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b1111111110001110; // vC= -114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b1111111100100000; // vC= -224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100100; // iC=-1820 
vC = 14'b1111111011111010; // vC= -262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b1111111100011101; // vC= -227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111101; // iC=-1667 
vC = 14'b1111111100010100; // vC= -236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b1111111101001111; // vC= -177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100100; // iC=-1820 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100101; // iC=-1691 
vC = 14'b1111111100101001; // vC= -215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b1111111011010010; // vC= -302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b1111111100001001; // vC= -247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001000; // iC=-1656 
vC = 14'b1111111100111011; // vC= -197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101101; // iC=-1683 
vC = 14'b1111111011100110; // vC= -282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b1111111011110111; // vC= -265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111101; // iC=-1667 
vC = 14'b1111111100100101; // vC= -219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b1111111100101001; // vC= -215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010100; // iC=-1644 
vC = 14'b1111111100101010; // vC= -214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101010; // iC=-1750 
vC = 14'b1111111100001010; // vC= -246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001000; // iC=-1656 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b1111111011011001; // vC= -295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b1111111011011100; // vC= -292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b1111111011001101; // vC= -307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b1111111011110001; // vC= -271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b1111111001111101; // vC= -387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010100; // iC=-1644 
vC = 14'b1111111001110000; // vC= -400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b1111111010101101; // vC= -339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b1111111010100011; // vC= -349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b1111111010111100; // vC= -324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101010; // iC=-1686 
vC = 14'b1111111001110100; // vC= -396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b1111111001101100; // vC= -404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b1111111011010001; // vC= -303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b1111111001111011; // vC= -389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011111; // iC=-1633 
vC = 14'b1111111010111001; // vC= -327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b1111111000111100; // vC= -452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b1111111010100011; // vC= -349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b1111111000101001; // vC= -471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b1111111000111010; // vC= -454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100011; // iC=-1629 
vC = 14'b1111111000010000; // vC= -496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b1111111001110111; // vC= -393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b1111111001010011; // vC= -429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b1111111000101111; // vC= -465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b1111110111101100; // vC= -532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b1111111001010011; // vC= -429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001101; // iC=-1651 
vC = 14'b1111111000010000; // vC= -496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b1111111000010000; // vC= -496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b1111111000101000; // vC= -472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b1111111001001001; // vC= -439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b1111110111010011; // vC= -557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111111; // iC=-1665 
vC = 14'b1111110111110100; // vC= -524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b1111111000111111; // vC= -449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011101; // iC=-1571 
vC = 14'b1111110111001110; // vC= -562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100101; // iC=-1691 
vC = 14'b1111110110110001; // vC= -591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b1111111000001011; // vC= -501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b1111111000101110; // vC= -466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010011; // iC=-1581 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b1111111000011001; // vC= -487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b1111111000010100; // vC= -492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b1111111000000101; // vC= -507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b1111111000011010; // vC= -486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b1111110110111000; // vC= -584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b1111110111001111; // vC= -561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b1111110110110011; // vC= -589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100011; // iC=-1565 
vC = 14'b1111110110110010; // vC= -590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110001; // iC=-1615 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011111; // iC=-1505 
vC = 14'b1111110111000111; // vC= -569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b1111110101111101; // vC= -643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010010; // iC=-1646 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b1111110111010001; // vC= -559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b1111110110000111; // vC= -633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110101; // iC=-1611 
vC = 14'b1111110101010011; // vC= -685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b1111110101000011; // vC= -701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b1111110110000110; // vC= -634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b1111110101011010; // vC= -678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000101; // iC=-1595 
vC = 14'b1111110100101110; // vC= -722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b1111110100101000; // vC= -728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101011; // iC=-1493 
vC = 14'b1111110110000000; // vC= -640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100100; // iC=-1500 
vC = 14'b1111110100111010; // vC= -710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b1111110100101101; // vC= -723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b1111110110000110; // vC= -634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b1111110011111010; // vC= -774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000110; // iC=-1466 
vC = 14'b1111110101000001; // vC= -703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b1111110100110111; // vC= -713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b1111110101111101; // vC= -643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110110; // iC=-1482 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100011; // iC=-1565 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100111; // iC=-1497 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111111; // iC=-1473 
vC = 14'b1111110011001101; // vC= -819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b1111110100010000; // vC= -752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011100; // iC=-1444 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b1111110100000000; // vC= -768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000100; // iC=-1468 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110110; // iC=-1418 
vC = 14'b1111110011110111; // vC= -777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b1111110100010110; // vC= -746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110111; // iC=-1481 
vC = 14'b1111110010101111; // vC= -849 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b1111110100001110; // vC= -754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b1111110100110001; // vC= -719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101011; // iC=-1429 
vC = 14'b1111110011011100; // vC= -804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111000; // iC=-1416 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101101; // iC=-1491 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b1111110010100011; // vC= -861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010111; // iC=-1385 
vC = 14'b1111110011110101; // vC= -779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b1111110011010001; // vC= -815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b1111110010000110; // vC= -890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b1111110011011111; // vC= -801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000110; // iC=-1466 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101000; // iC=-1432 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110101; // iC=-1419 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111000; // iC=-1352 
vC = 14'b1111110001101010; // vC= -918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001111; // iC=-1393 
vC = 14'b1111110010010010; // vC= -878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111101; // iC=-1475 
vC = 14'b1111110011100010; // vC= -798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000101; // iC=-1339 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b1111110001111011; // vC= -901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001010; // iC=-1398 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001011; // iC=-1397 
vC = 14'b1111110000111100; // vC= -964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b1111110011000010; // vC= -830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010110; // iC=-1322 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001110; // iC=-1394 
vC = 14'b1111110000111111; // vC= -961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011110; // iC=-1442 
vC = 14'b1111110000101011; // vC= -981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100100; // iC=-1372 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100100; // iC=-1436 
vC = 14'b1111110001000101; // vC= -955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110010; // iC=-1294 
vC = 14'b1111110000111100; // vC= -964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011101; // iC=-1379 
vC = 14'b1111110000100111; // vC= -985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101111; // iC=-1361 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010111; // iC=-1321 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000000; // iC=-1344 
vC = 14'b1111110001101111; // vC= -913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111100; // iC=-1284 
vC = 14'b1111110001001111; // vC= -945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111101; // iC=-1347 
vC = 14'b1111101111111010; // vC=-1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100100; // iC=-1244 
vC = 14'b1111110000111111; // vC= -961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001010; // iC=-1334 
vC = 14'b1111110000011000; // vC=-1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000111; // iC=-1337 
vC = 14'b1111101111110011; // vC=-1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000000; // iC=-1344 
vC = 14'b1111101111101111; // vC=-1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100110; // iC=-1306 
vC = 14'b1111110000001001; // vC=-1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010100; // iC=-1324 
vC = 14'b1111110001000010; // vC= -958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000010; // iC=-1342 
vC = 14'b1111110000101101; // vC= -979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111100; // iC=-1348 
vC = 14'b1111101111111111; // vC=-1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110100; // iC=-1292 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110110; // iC=-1226 
vC = 14'b1111110001001110; // vC= -946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110100; // iC=-1228 
vC = 14'b1111101111001101; // vC=-1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100000; // iC=-1312 
vC = 14'b1111110000011010; // vC= -998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110011; // iC=-1229 
vC = 14'b1111110000010101; // vC=-1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111110001000010; // vC= -958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001111; // iC=-1265 
vC = 14'b1111110000110100; // vC= -972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000111; // iC=-1337 
vC = 14'b1111101111011001; // vC=-1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010000; // iC=-1264 
vC = 14'b1111101110111111; // vC=-1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011111; // iC=-1313 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101000; // iC=-1176 
vC = 14'b1111101110100110; // vC=-1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000101; // iC=-1211 
vC = 14'b1111101111001100; // vC=-1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100001; // iC=-1247 
vC = 14'b1111101110101001; // vC=-1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011111; // iC=-1185 
vC = 14'b1111101110010100; // vC=-1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b1111101110110000; // vC=-1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001100; // iC=-1268 
vC = 14'b1111101111111010; // vC=-1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000111; // iC=-1145 
vC = 14'b1111101111110110; // vC=-1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000100; // iC=-1276 
vC = 14'b1111101111111101; // vC=-1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010000; // iC=-1200 
vC = 14'b1111101110011111; // vC=-1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101010; // iC=-1238 
vC = 14'b1111101111101100; // vC=-1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011111; // iC=-1121 
vC = 14'b1111101111000011; // vC=-1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101011; // iC=-1173 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001111; // iC=-1265 
vC = 14'b1111101110101000; // vC=-1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111100; // iC=-1156 
vC = 14'b1111101110101000; // vC=-1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101011; // iC=-1237 
vC = 14'b1111101110100101; // vC=-1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011110; // iC=-1186 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011010; // iC=-1126 
vC = 14'b1111101111000111; // vC=-1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101100; // iC=-1172 
vC = 14'b1111101111100000; // vC=-1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000110; // iC=-1210 
vC = 14'b1111101101111110; // vC=-1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001010; // iC=-1206 
vC = 14'b1111101110010010; // vC=-1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000110; // iC=-1082 
vC = 14'b1111101110101110; // vC=-1106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011000; // iC=-1192 
vC = 14'b1111101110101101; // vC=-1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111100; // iC=-1220 
vC = 14'b1111101101010000; // vC=-1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000000; // iC=-1152 
vC = 14'b1111101101010011; // vC=-1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000101; // iC=-1211 
vC = 14'b1111101110110001; // vC=-1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011001; // iC=-1191 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001011; // iC=-1077 
vC = 14'b1111101101100100; // vC=-1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000001; // iC=-1087 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001110; // iC=-1074 
vC = 14'b1111101110110100; // vC=-1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000011; // iC=-1149 
vC = 14'b1111101100100000; // vC=-1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010111; // iC=-1065 
vC = 14'b1111101110001001; // vC=-1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000000; // iC=-1152 
vC = 14'b1111101100101001; // vC=-1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101000; // iC=-1112 
vC = 14'b1111101110010110; // vC=-1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010000; // iC=-1136 
vC = 14'b1111101110001111; // vC=-1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100101; // iC=-1051 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011101; // iC=-1059 
vC = 14'b1111101110000110; // vC=-1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011011; // iC= -997 
vC = 14'b1111101101110111; // vC=-1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001011; // iC=-1013 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001001; // iC=-1015 
vC = 14'b1111101110000111; // vC=-1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101110; // iC= -978 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101001; // iC= -983 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110011; // iC= -973 
vC = 14'b1111101100100100; // vC=-1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111101101100010; // vC=-1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101010; // iC=-1110 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000110; // iC=-1082 
vC = 14'b1111101100010000; // vC=-1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001000; // iC= -952 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011111; // iC=-1057 
vC = 14'b1111101011100010; // vC=-1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010001; // iC= -943 
vC = 14'b1111101100100110; // vC=-1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101111; // iC=-1041 
vC = 14'b1111101100000111; // vC=-1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000001; // iC= -959 
vC = 14'b1111101100110111; // vC=-1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000010; // iC= -958 
vC = 14'b1111101011101010; // vC=-1302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110110; // iC=-1034 
vC = 14'b1111101100101001; // vC=-1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100101; // iC=-1051 
vC = 14'b1111101101000010; // vC=-1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010000; // iC= -944 
vC = 14'b1111101011001001; // vC=-1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001111; // iC=-1009 
vC = 14'b1111101011110111; // vC=-1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101111; // iC= -977 
vC = 14'b1111101100000111; // vC=-1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011010; // iC= -934 
vC = 14'b1111101101011010; // vC=-1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001000; // iC= -952 
vC = 14'b1111101101010011; // vC=-1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000111; // iC= -889 
vC = 14'b1111101100111101; // vC=-1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111100; // iC=-1028 
vC = 14'b1111101011111111; // vC=-1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000101; // iC= -955 
vC = 14'b1111101101000001; // vC=-1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b1111101101001000; // vC=-1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000000; // iC= -960 
vC = 14'b1111101011101111; // vC=-1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101001; // iC= -983 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111110; // iC= -962 
vC = 14'b1111101011110101; // vC=-1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011111; // iC= -865 
vC = 14'b1111101100101000; // vC=-1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110011; // iC= -909 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011111; // iC= -865 
vC = 14'b1111101100100011; // vC=-1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011011; // iC= -869 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101101; // iC= -979 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010110; // iC= -938 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000011; // iC= -893 
vC = 14'b1111101010001111; // vC=-1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110010; // iC= -910 
vC = 14'b1111101010010101; // vC=-1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001000; // iC= -952 
vC = 14'b1111101011111110; // vC=-1282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101001; // iC= -919 
vC = 14'b1111101011110111; // vC=-1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101100; // iC= -852 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010010; // iC= -878 
vC = 14'b1111101010111011; // vC=-1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111011; // iC= -901 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110101; // iC= -843 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110111; // iC= -777 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110100; // iC= -780 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111101; // iC= -771 
vC = 14'b1111101011100100; // vC=-1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000111; // iC= -889 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101011; // iC= -789 
vC = 14'b1111101010000011; // vC=-1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111111; // iC= -897 
vC = 14'b1111101001111101; // vC=-1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111101; // iC= -835 
vC = 14'b1111101001110001; // vC=-1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001101; // iC= -883 
vC = 14'b1111101010111010; // vC=-1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111100; // iC= -836 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111110; // iC= -834 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010010; // iC= -814 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001100; // iC= -756 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100111; // iC= -729 
vC = 14'b1111101001100110; // vC=-1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100010; // iC= -734 
vC = 14'b1111101011010110; // vC=-1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100111; // iC= -729 
vC = 14'b1111101010000010; // vC=-1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001000; // iC= -696 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100101; // iC= -795 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001000; // iC= -760 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100000; // iC= -800 
vC = 14'b1111101010100100; // vC=-1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100111; // iC= -729 
vC = 14'b1111101000110110; // vC=-1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111101; // iC= -707 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011010; // iC= -806 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001110; // iC= -690 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101001; // iC= -791 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100100; // iC= -732 
vC = 14'b1111101000110111; // vC=-1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111000; // iC= -648 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010111; // iC= -745 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010010; // iC= -686 
vC = 14'b1111101010110101; // vC=-1355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110001; // iC= -655 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010111; // iC= -617 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101101; // iC= -659 
vC = 14'b1111101000110001; // vC=-1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100000; // iC= -672 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100001; // iC= -671 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100001; // iC= -735 
vC = 14'b1111101001110101; // vC=-1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110110; // iC= -714 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001000; // iC= -568 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001010; // iC= -694 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100000; // iC= -672 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101100; // iC= -660 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010010; // iC= -686 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010000; // iC= -560 
vC = 14'b1111101000000011; // vC=-1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111011; // iC= -645 
vC = 14'b1111101000010010; // vC=-1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010001; // iC= -559 
vC = 14'b1111101010011010; // vC=-1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100111; // iC= -601 
vC = 14'b1111101001101001; // vC=-1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010101; // iC= -619 
vC = 14'b1111101001111110; // vC=-1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000001; // iC= -639 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010101; // iC= -619 
vC = 14'b1111101010010001; // vC=-1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000101; // iC= -571 
vC = 14'b1111101010001011; // vC=-1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000111; // iC= -505 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111111; // iC= -513 
vC = 14'b1111101001110011; // vC=-1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000111; // iC= -569 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100011; // iC= -541 
vC = 14'b1111101001011110; // vC=-1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010110; // iC= -490 
vC = 14'b1111100111110000; // vC=-1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100110; // iC= -538 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001001; // iC= -567 
vC = 14'b1111100111111100; // vC=-1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101000; // iC= -472 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101111; // iC= -465 
vC = 14'b1111100111110100; // vC=-1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000101; // iC= -571 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110110; // iC= -586 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001111; // iC= -433 
vC = 14'b1111100111100011; // vC=-1565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100011; // iC= -477 
vC = 14'b1111100111100010; // vC=-1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101011; // iC= -469 
vC = 14'b1111101001101110; // vC=-1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011101; // iC= -483 
vC = 14'b1111101001100111; // vC=-1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000010; // iC= -510 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100101; // iC= -411 
vC = 14'b1111100111011101; // vC=-1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000011; // iC= -509 
vC = 14'b1111101000110110; // vC=-1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100010; // iC= -478 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000100; // iC= -508 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010101; // iC= -427 
vC = 14'b1111101001001111; // vC=-1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000111; // iC= -505 
vC = 14'b1111101000001001; // vC=-1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101001; // iC= -471 
vC = 14'b1111101000111011; // vC=-1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111010; // iC= -454 
vC = 14'b1111101000001101; // vC=-1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010110; // iC= -426 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010110001; // iC= -335 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010100; // iC= -428 
vC = 14'b1111100111110100; // vC=-1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111001; // iC= -391 
vC = 14'b1111100111010110; // vC=-1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011000; // iC= -424 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000100; // iC= -316 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000101; // iC= -251 
vC = 14'b1111100111101001; // vC=-1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000110; // iC= -378 
vC = 14'b1111101000010001; // vC=-1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010010; // iC= -238 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100001; // iC= -351 
vC = 14'b1111100111000011; // vC=-1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101000; // iC= -216 
vC = 14'b1111101000010111; // vC=-1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000100; // iC= -188 
vC = 14'b1111100111001001; // vC=-1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000001; // iC= -255 
vC = 14'b1111100111010111; // vC=-1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011010; // iC= -230 
vC = 14'b1111100111100001; // vC=-1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110000; // iC= -208 
vC = 14'b1111100111110101; // vC=-1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101001; // iC= -215 
vC = 14'b1111101000110111; // vC=-1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100001; // iC= -159 
vC = 14'b1111100111110000; // vC=-1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010101; // iC= -107 
vC = 14'b1111100111011010; // vC=-1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111100; // iC= -132 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111000; // iC=  -72 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011001; // iC= -103 
vC = 14'b1111101000011001; // vC=-1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100101; // iC= -155 
vC = 14'b1111100111001100; // vC=-1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000010; // iC= -126 
vC = 14'b1111100111111011; // vC=-1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100111; // iC=  -89 
vC = 14'b1111101001000110; // vC=-1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111010; // iC= -134 
vC = 14'b1111100111101011; // vC=-1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101101; // iC=  -19 
vC = 14'b1111101001000000; // vC=-1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011101; // iC=   29 
vC = 14'b1111100111000001; // vC=-1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000001; // iC=    1 
vC = 14'b1111101000010010; // vC=-1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010010; // iC=   18 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001011; // iC=   75 
vC = 14'b1111101000000001; // vC=-1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110101; // iC=  -11 
vC = 14'b1111101000010101; // vC=-1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001101; // iC=   77 
vC = 14'b1111100111010111; // vC=-1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001110; // iC=  142 
vC = 14'b1111101000000100; // vC=-1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110011; // iC=   51 
vC = 14'b1111100111100110; // vC=-1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000111; // iC=  199 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110110; // iC=  118 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001110; // iC=  206 
vC = 14'b1111101001001110; // vC=-1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111101; // iC=  189 
vC = 14'b1111100111011111; // vC=-1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000110; // iC=  326 
vC = 14'b1111101000111010; // vC=-1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000101; // iC=  197 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010010; // iC=  210 
vC = 14'b1111101000111110; // vC=-1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101011; // iC=  299 
vC = 14'b1111101000000010; // vC=-1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000001; // iC=  385 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100011; // iC=  355 
vC = 14'b1111100111100100; // vC=-1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101100; // iC=  428 
vC = 14'b1111101001001000; // vC=-1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011101; // iC=  349 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011001; // iC=  473 
vC = 14'b1111101000001111; // vC=-1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110110; // iC=  438 
vC = 14'b1111101000011101; // vC=-1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001000; // iC=  456 
vC = 14'b1111101001001111; // vC=-1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100100; // iC=  548 
vC = 14'b1111101000011100; // vC=-1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111000; // iC=  504 
vC = 14'b1111100111101110; // vC=-1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111001; // iC=  505 
vC = 14'b1111100111010110; // vC=-1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001000; // iC=  520 
vC = 14'b1111101001001111; // vC=-1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110101; // iC=  629 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110011; // iC=  691 
vC = 14'b1111101001001001; // vC=-1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101101; // iC=  621 
vC = 14'b1111100111110010; // vC=-1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010111; // iC=  727 
vC = 14'b1111101000000000; // vC=-1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001101; // iC=  717 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010101; // iC=  661 
vC = 14'b1111100111111110; // vC=-1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010111; // iC=  791 
vC = 14'b1111101000101100; // vC=-1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101001; // iC=  745 
vC = 14'b1111100111101101; // vC=-1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111011; // iC=  763 
vC = 14'b1111101001110000; // vC=-1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110110; // iC=  758 
vC = 14'b1111100111111101; // vC=-1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011100; // iC=  860 
vC = 14'b1111101000000010; // vC=-1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000101; // iC=  773 
vC = 14'b1111101001100101; // vC=-1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110011; // iC=  947 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010001; // iC=  977 
vC = 14'b1111101000011111; // vC=-1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010001; // iC=  913 
vC = 14'b1111101000000100; // vC=-1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110111; // iC=  887 
vC = 14'b1111101000110001; // vC=-1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001001; // iC=  905 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000100; // iC= 1028 
vC = 14'b1111101001101101; // vC=-1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110010; // iC= 1074 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100001; // iC= 1057 
vC = 14'b1111101001011001; // vC=-1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001100; // iC=  972 
vC = 14'b1111101010010110; // vC=-1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110001; // iC= 1137 
vC = 14'b1111101010101100; // vC=-1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010100; // iC= 1044 
vC = 14'b1111101001100100; // vC=-1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000111; // iC= 1095 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110010; // iC= 1074 
vC = 14'b1111101010000010; // vC=-1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100100; // iC= 1124 
vC = 14'b1111101010101010; // vC=-1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110101; // iC= 1205 
vC = 14'b1111101000101100; // vC=-1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001111; // iC= 1231 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110111; // iC= 1271 
vC = 14'b1111101000110000; // vC=-1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000101; // iC= 1285 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101001; // iC= 1193 
vC = 14'b1111101010010010; // vC=-1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101011; // iC= 1323 
vC = 14'b1111101010010111; // vC=-1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011111; // iC= 1247 
vC = 14'b1111101001011000; // vC=-1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100001; // iC= 1313 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001011; // iC= 1291 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001001; // iC= 1289 
vC = 14'b1111101001111101; // vC=-1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001011; // iC= 1291 
vC = 14'b1111101001100100; // vC=-1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000101; // iC= 1349 
vC = 14'b1111101010111100; // vC=-1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100010; // iC= 1442 
vC = 14'b1111101010010110; // vC=-1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b1111101011101110; // vC=-1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000100; // iC= 1412 
vC = 14'b1111101010010000; // vC=-1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000100; // iC= 1476 
vC = 14'b1111101010010010; // vC=-1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111001; // iC= 1465 
vC = 14'b1111101011101010; // vC=-1302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010011; // iC= 1427 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111110; // iC= 1534 
vC = 14'b1111101011011000; // vC=-1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010111; // iC= 1431 
vC = 14'b1111101011000001; // vC=-1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000101; // iC= 1477 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111000; // iC= 1592 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110000; // iC= 1584 
vC = 14'b1111101010100111; // vC=-1369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b1111101011001111; // vC=-1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111100; // iC= 1596 
vC = 14'b1111101100011000; // vC=-1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110011; // iC= 1587 
vC = 14'b1111101100100101; // vC=-1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110100; // iC= 1652 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011111; // iC= 1567 
vC = 14'b1111101101001001; // vC=-1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011010; // iC= 1562 
vC = 14'b1111101011101001; // vC=-1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101001; // iC= 1705 
vC = 14'b1111101011010111; // vC=-1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b1111101011010010; // vC=-1326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010001; // iC= 1745 
vC = 14'b1111101100011000; // vC=-1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000010; // iC= 1730 
vC = 14'b1111101011011011; // vC=-1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100000; // iC= 1632 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100001; // iC= 1633 
vC = 14'b1111101101111110; // vC=-1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b1111101110000110; // vC=-1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b1111101011101111; // vC=-1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111101101110110; // vC=-1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000101; // iC= 1797 
vC = 14'b1111101101100011; // vC=-1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111110; // iC= 1790 
vC = 14'b1111101101110010; // vC=-1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101110; // iC= 1710 
vC = 14'b1111101100111010; // vC=-1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b1111101110101100; // vC=-1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b1111101110011110; // vC=-1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b1111101100101001; // vC=-1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100000; // iC= 1824 
vC = 14'b1111101101100101; // vC=-1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111101101001001; // vC=-1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111101101111000; // vC=-1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b1111101110100000; // vC=-1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110110; // iC= 1846 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110110; // iC= 1846 
vC = 14'b1111101111111001; // vC=-1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b1111101110100010; // vC=-1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b1111101111111111; // vC=-1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111101111010111; // vC=-1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111110000001111; // vC=-1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b1111101111110101; // vC=-1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b1111110000000111; // vC=-1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b1111101111010001; // vC=-1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b1111101110100010; // vC=-1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b1111110000001110; // vC=-1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010010; // iC= 1874 
vC = 14'b1111101111001101; // vC=-1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b1111101111110010; // vC=-1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111110000100101; // vC= -987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b1111101111011101; // vC=-1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b1111101111111101; // vC=-1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110010; // iC= 1906 
vC = 14'b1111110001100000; // vC= -928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b1111110001000011; // vC= -957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111101111111000; // vC=-1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b1111110000110101; // vC= -971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b1111110000111111; // vC= -961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b1111110001100000; // vC= -928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111110010010001; // vC= -879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011101; // iC= 2013 
vC = 14'b1111110001110010; // vC= -910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110100; // iC= 1972 
vC = 14'b1111110010000111; // vC= -889 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100001; // iC= 2017 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b1111110000111111; // vC= -961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111110000100100; // vC= -988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111110010000101; // vC= -891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b1111110011000010; // vC= -830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111110; // iC= 1982 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111110001000110; // vC= -954 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111110011011001; // vC= -807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111110001111100; // vC= -900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111110011100111; // vC= -793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000011; // iC= 2051 
vC = 14'b1111110011001001; // vC= -823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b1111110001111111; // vC= -897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111110010001111; // vC= -881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111110100000100; // vC= -764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111110010011101; // vC= -867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111110100001111; // vC= -753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b1111110011000010; // vC= -830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111110011001111; // vC= -817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111110100000101; // vC= -763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b1111110100011101; // vC= -739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111110011110100; // vC= -780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110011001001; // vC= -823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b1111110100101100; // vC= -724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111110100111101; // vC= -707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111110100000100; // vC= -764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010001; // iC= 2065 
vC = 14'b1111110101010001; // vC= -687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111110100111110; // vC= -706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b1111110101000001; // vC= -703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111101; // iC= 2045 
vC = 14'b1111110101010100; // vC= -684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000000; // iC= 2048 
vC = 14'b1111110100011110; // vC= -738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b1111110101000001; // vC= -703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001110; // iC= 2062 
vC = 14'b1111110110010011; // vC= -621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100001; // iC= 2017 
vC = 14'b1111110110110101; // vC= -587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111110110010010; // vC= -622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011010; // iC= 2074 
vC = 14'b1111110101111010; // vC= -646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101111; // iC= 2031 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b1111110101110011; // vC= -653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111110111110100; // vC= -524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111110111011001; // vC= -551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b1111110111111101; // vC= -515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010110; // iC= 2070 
vC = 14'b1111110111001110; // vC= -562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111110111001010; // vC= -566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101011; // iC= 2027 
vC = 14'b1111111000001010; // vC= -502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b1111110111101111; // vC= -529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111110110110000; // vC= -592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111110110011011; // vC= -613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111110111001011; // vC= -565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111110111110010; // vC= -526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100110; // iC= 2086 
vC = 14'b1111111000000000; // vC= -512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111111000001111; // vC= -497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100011; // iC= 2083 
vC = 14'b1111111001001111; // vC= -433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000101101; // iC= 2093 
vC = 14'b1111110111111010; // vC= -518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111110111011000; // vC= -552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000110010; // iC= 2098 
vC = 14'b1111111000110110; // vC= -458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000110100; // iC= 2100 
vC = 14'b1111111000111110; // vC= -450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111111000010101; // vC= -491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001010; // iC= 1994 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000000; // iC= 1984 
vC = 14'b1111111000110001; // vC= -463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111111010001011; // vC= -373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b1111111001111010; // vC= -390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111111001111100; // vC= -388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b1111111010011100; // vC= -356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000100; // iC= 2052 
vC = 14'b1111111001010101; // vC= -427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b1111111000111010; // vC= -454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111111001010111; // vC= -425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111111000111001; // vC= -455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111111010010011; // vC= -365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101101; // iC= 2029 
vC = 14'b1111111010011100; // vC= -356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111111010111101; // vC= -323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111111010100111; // vC= -345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111111010011111; // vC= -353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011110; // iC= 2078 
vC = 14'b1111111001111001; // vC= -391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100110; // iC= 2086 
vC = 14'b1111111010001000; // vC= -376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111111011000110; // vC= -314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000110000; // iC= 2096 
vC = 14'b1111111011010111; // vC= -297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b1111111010001110; // vC= -370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111111001110011; // vC= -397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000101010; // iC= 2090 
vC = 14'b1111111100001111; // vC= -241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111111010111000; // vC= -328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100110; // iC= 2086 
vC = 14'b1111111010001001; // vC= -375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111010100100; // vC= -348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010100; // iC= 2068 
vC = 14'b1111111010110000; // vC= -336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000101; // iC= 2053 
vC = 14'b1111111010110011; // vC= -333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111111100001011; // vC= -245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011100; // iC= 1948 
vC = 14'b1111111010111000; // vC= -328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111111011110011; // vC= -269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111111100110100; // vC= -204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000110010; // iC= 2098 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b1111111100011010; // vC= -230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111111011111011; // vC= -261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010001; // iC= 2065 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b1111111011110100; // vC= -268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111100001011; // vC= -245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100011; // iC= 2083 
vC = 14'b1111111011111101; // vC= -259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010100; // iC= 2068 
vC = 14'b1111111101100000; // vC= -160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b1111111101001011; // vC= -181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000011; // iC= 2051 
vC = 14'b1111111101100100; // vC= -156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111111101001000; // vC= -184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111111101110100; // vC= -140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111111101111011; // vC= -133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100111; // iC= 2087 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111111110001110; // vC= -114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010011; // iC= 2067 
vC = 14'b1111111110111101; // vC=  -67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111111101000110; // vC= -186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111111101011111; // vC= -161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010110; // iC= 2070 
vC = 14'b1111111101010010; // vC= -174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b1111111101011101; // vC= -163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001010; // iC= 2058 
vC = 14'b1111111110011100; // vC= -100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010100; // iC= 2004 
vC = 14'b1111111111111000; // vC=   -8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110010; // iC= 2034 
vC = 14'b1111111110100001; // vC=  -95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b1111111110110011; // vC=  -77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b1111111110111011; // vC=  -69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b0000000000010111; // vC=   23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111111110110011; // vC=  -77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001010; // iC= 2058 
vC = 14'b0000000000010100; // vC=   20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110010; // iC= 2034 
vC = 14'b1111111111110111; // vC=   -9 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b0000000000101010; // vC=   42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b0000000000101000; // vC=   40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110010; // iC= 2034 
vC = 14'b1111111111110101; // vC=  -11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b1111111111011011; // vC=  -37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b0000000000111000; // vC=   56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b1111111111111010; // vC=   -6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b1111111111011101; // vC=  -35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001010; // iC= 1994 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111111111100110; // vC=  -26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000011; // iC= 2051 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001011; // iC= 2059 
vC = 14'b0000000000000101; // vC=    5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011011; // iC= 2011 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000111; // iC= 1991 
vC = 14'b0000000000111101; // vC=   61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010100; // iC= 2004 
vC = 14'b0000000000011101; // vC=   29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b0000000000001110; // vC=   14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000111; // iC= 2055 
vC = 14'b0000000000110111; // vC=   55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b0000000000110101; // vC=   53 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b0000000010001100; // vC=  140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101111; // iC= 2031 
vC = 14'b0000000010011000; // vC=  152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000001; // iC= 2049 
vC = 14'b0000000000111011; // vC=   59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b0000000001101011; // vC=  107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b0000000011000111; // vC=  199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b0000000001111001; // vC=  121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b0000000001010111; // vC=   87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b0000000010101110; // vC=  174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b0000000011101000; // vC=  232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b0000000001111000; // vC=  120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001010; // iC= 1994 
vC = 14'b0000000010011000; // vC=  152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b0000000010000011; // vC=  131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100010; // iC= 2018 
vC = 14'b0000000010001101; // vC=  141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b0000000010001101; // vC=  141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b0000000010010111; // vC=  151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b0000000010000101; // vC=  133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101100; // iC= 1964 
vC = 14'b0000000010010111; // vC=  151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b0000000010010111; // vC=  151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b0000000100000000; // vC=  256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b0000000100010010; // vC=  274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b0000000011000101; // vC=  197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011000; // iC= 1880 
vC = 14'b0000000011100001; // vC=  225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b0000000011110011; // vC=  243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b0000000010111111; // vC=  191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010010; // iC= 1874 
vC = 14'b0000000101001111; // vC=  335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b0000000100011110; // vC=  286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b0000000100110110; // vC=  310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b0000000011100111; // vC=  231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b0000000100101101; // vC=  301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b0000000100100001; // vC=  289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b0000000101000001; // vC=  321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b0000000101010011; // vC=  339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b0000000110001010; // vC=  394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010100; // iC= 1876 
vC = 14'b0000000100100000; // vC=  288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b0000000110011010; // vC=  410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b0000000100010111; // vC=  279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b0000000101000110; // vC=  326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b0000000101101101; // vC=  365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b0000000101100000; // vC=  352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010001; // iC= 1873 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b0000000111001100; // vC=  460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b0000000110100111; // vC=  423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b0000000101000010; // vC=  322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b0000000110101001; // vC=  425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b0000000110101101; // vC=  429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b0000000111101010; // vC=  490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b0000000110011010; // vC=  410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b0000000101100010; // vC=  354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000000111010100; // vC=  468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000101; // iC= 1797 
vC = 14'b0000000111100010; // vC=  482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b0000001000000110; // vC=  518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b0000001000010111; // vC=  535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b0000000111111000; // vC=  504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b0000000111100101; // vC=  485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b0000000111111101; // vC=  509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b0000001000100000; // vC=  544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000000110101111; // vC=  431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b0000000110110111; // vC=  439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000010; // iC= 1858 
vC = 14'b0000000110111001; // vC=  441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b0000000111000111; // vC=  455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000001000010101; // vC=  533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b0000001001011100; // vC=  604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b0000001001101001; // vC=  617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b0000001000111101; // vC=  573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011000; // iC= 1880 
vC = 14'b0000000111101101; // vC=  493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b0000001000111011; // vC=  571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111101; // iC= 1853 
vC = 14'b0000001000101010; // vC=  554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101011; // iC= 1835 
vC = 14'b0000000111101010; // vC=  490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110001; // iC= 1777 
vC = 14'b0000001001101110; // vC=  622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b0000001000001001; // vC=  521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b0000001001000011; // vC=  579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b0000000111111101; // vC=  509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011000; // iC= 1752 
vC = 14'b0000001000101001; // vC=  553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b0000001010000100; // vC=  644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000001000111000; // vC=  568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b0000001000101110; // vC=  558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111100; // iC= 1724 
vC = 14'b0000001001100111; // vC=  615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b0000001001101000; // vC=  616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b0000001010010000; // vC=  656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000110; // iC= 1798 
vC = 14'b0000001001110011; // vC=  627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b0000001010010110; // vC=  662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b0000001001001010; // vC=  586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001001; // iC= 1737 
vC = 14'b0000001010100100; // vC=  676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111011; // iC= 1851 
vC = 14'b0000001011011010; // vC=  730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000110; // iC= 1798 
vC = 14'b0000001011100011; // vC=  739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000110; // iC= 1734 
vC = 14'b0000001011001010; // vC=  714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b0000001001111101; // vC=  637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b0000001010111111; // vC=  703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b0000001100001000; // vC=  776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b0000001001110110; // vC=  630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b0000001011010000; // vC=  720 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100011; // iC= 1699 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111000; // iC= 1720 
vC = 14'b0000001010001001; // vC=  649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b0000001010010000; // vC=  656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b0000001100000111; // vC=  775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b0000001011011011; // vC=  731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000000; // iC= 1664 
vC = 14'b0000001011101100; // vC=  748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000001011011100; // vC=  732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101001; // iC= 1705 
vC = 14'b0000001011011111; // vC=  735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000001101011110; // vC=  862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010100; // iC= 1620 
vC = 14'b0000001011100101; // vC=  741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101011; // iC= 1707 
vC = 14'b0000001100111010; // vC=  826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100010; // iC= 1634 
vC = 14'b0000001101100100; // vC=  868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000001100011011; // vC=  795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011110; // iC= 1630 
vC = 14'b0000001011110111; // vC=  759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b0000001101100101; // vC=  869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100010; // iC= 1634 
vC = 14'b0000001101110001; // vC=  881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110011; // iC= 1651 
vC = 14'b0000001110000011; // vC=  899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000000; // iC= 1600 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101110; // iC= 1582 
vC = 14'b0000001100010001; // vC=  785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000110; // iC= 1606 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001011; // iC= 1611 
vC = 14'b0000001101111000; // vC=  888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101011; // iC= 1579 
vC = 14'b0000001110000111; // vC=  903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101001; // iC= 1577 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010001; // iC= 1617 
vC = 14'b0000001101010100; // vC=  852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101100; // iC= 1580 
vC = 14'b0000001101111000; // vC=  888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101111; // iC= 1647 
vC = 14'b0000001101111111; // vC=  895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100110; // iC= 1574 
vC = 14'b0000001101010010; // vC=  850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b0000001110110101; // vC=  949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000101; // iC= 1605 
vC = 14'b0000001110000100; // vC=  900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000010; // iC= 1538 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001111011101; // vC=  989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110101; // iC= 1653 
vC = 14'b0000001111101100; // vC= 1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001101110101; // vC=  885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b0000001101100001; // vC=  865 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011100; // iC= 1628 
vC = 14'b0000001101100100; // vC=  868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010001; // iC= 1553 
vC = 14'b0000001111111001; // vC= 1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111011; // iC= 1595 
vC = 14'b0000001101111111; // vC=  895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010100; // iC= 1620 
vC = 14'b0000001101111001; // vC=  889 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b0000001101110011; // vC=  883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011100; // iC= 1564 
vC = 14'b0000001110001110; // vC=  910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000001111010101; // vC=  981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110100; // iC= 1524 
vC = 14'b0000001110100110; // vC=  934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101000; // iC= 1512 
vC = 14'b0000001110111000; // vC=  952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100101; // iC= 1509 
vC = 14'b0000001110101101; // vC=  941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100101; // iC= 1509 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010111; // iC= 1559 
vC = 14'b0000010000100000; // vC= 1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001111101011; // vC= 1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010100; // iC= 1556 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111000; // iC= 1528 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001010; // iC= 1482 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101011; // iC= 1579 
vC = 14'b0000001111001100; // vC=  972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100101; // iC= 1509 
vC = 14'b0000001111101001; // vC= 1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101001; // iC= 1577 
vC = 14'b0000010000001001; // vC= 1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101001; // iC= 1449 
vC = 14'b0000010001011100; // vC= 1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101000; // iC= 1448 
vC = 14'b0000010000100110; // vC= 1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100111; // iC= 1575 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100101; // iC= 1509 
vC = 14'b0000010001000111; // vC= 1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b0000010000110000; // vC= 1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010100; // iC= 1428 
vC = 14'b0000010001101101; // vC= 1133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011001; // iC= 1433 
vC = 14'b0000010000110100; // vC= 1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001100; // iC= 1484 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101101; // iC= 1453 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010111; // iC= 1495 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100101; // iC= 1509 
vC = 14'b0000010000101011; // vC= 1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101010; // iC= 1514 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111110; // iC= 1406 
vC = 14'b0000010001111011; // vC= 1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001111; // iC= 1487 
vC = 14'b0000010000000101; // vC= 1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000010; // iC= 1410 
vC = 14'b0000010001000000; // vC= 1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101010; // iC= 1386 
vC = 14'b0000010010101001; // vC= 1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111111; // iC= 1471 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100100; // iC= 1444 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011100; // iC= 1500 
vC = 14'b0000010001100001; // vC= 1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001101; // iC= 1357 
vC = 14'b0000010000101111; // vC= 1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001100; // iC= 1420 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000101; // iC= 1477 
vC = 14'b0000010010011010; // vC= 1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100000; // iC= 1440 
vC = 14'b0000010001110000; // vC= 1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101111; // iC= 1455 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000100; // iC= 1348 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011000; // iC= 1432 
vC = 14'b0000010001001110; // vC= 1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010010; // iC= 1426 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011101; // iC= 1373 
vC = 14'b0000010011001011; // vC= 1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100001; // iC= 1313 
vC = 14'b0000010010100010; // vC= 1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000001; // iC= 1345 
vC = 14'b0000010011001100; // vC= 1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110010; // iC= 1394 
vC = 14'b0000010011010110; // vC= 1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010101; // iC= 1429 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101001; // iC= 1385 
vC = 14'b0000010011101111; // vC= 1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100010; // iC= 1378 
vC = 14'b0000010001101100; // vC= 1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111101; // iC= 1405 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110101; // iC= 1333 
vC = 14'b0000010010010100; // vC= 1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011000; // iC= 1368 
vC = 14'b0000010100001000; // vC= 1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001111; // iC= 1295 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111100; // iC= 1276 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101100; // iC= 1324 
vC = 14'b0000010011100010; // vC= 1250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011111; // iC= 1247 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100100; // iC= 1316 
vC = 14'b0000010011101110; // vC= 1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001111; // iC= 1231 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111101; // iC= 1277 
vC = 14'b0000010010001111; // vC= 1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001010; // iC= 1290 
vC = 14'b0000010010100000; // vC= 1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110001; // iC= 1265 
vC = 14'b0000010011100001; // vC= 1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100011; // iC= 1315 
vC = 14'b0000010100101100; // vC= 1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100111; // iC= 1255 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101010; // iC= 1322 
vC = 14'b0000010010101100; // vC= 1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111001; // iC= 1209 
vC = 14'b0000010010111111; // vC= 1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000010; // iC= 1218 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001111; // iC= 1231 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101110; // iC= 1262 
vC = 14'b0000010010110001; // vC= 1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000001; // iC= 1281 
vC = 14'b0000010011100011; // vC= 1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010011; // iC= 1235 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001100; // iC= 1228 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001110; // iC= 1294 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100010; // iC= 1186 
vC = 14'b0000010011001111; // vC= 1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110110; // iC= 1206 
vC = 14'b0000010100100101; // vC= 1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000101; // iC= 1285 
vC = 14'b0000010100001101; // vC= 1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100111; // iC= 1255 
vC = 14'b0000010101100011; // vC= 1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110100; // iC= 1268 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101011; // iC= 1131 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000010; // iC= 1282 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110001; // iC= 1201 
vC = 14'b0000010100011100; // vC= 1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110101; // iC= 1141 
vC = 14'b0000010101100011; // vC= 1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001011; // iC= 1227 
vC = 14'b0000010101100100; // vC= 1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111001; // iC= 1145 
vC = 14'b0000010011111011; // vC= 1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010110; // iC= 1174 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111110; // iC= 1214 
vC = 14'b0000010011110101; // vC= 1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100110; // iC= 1190 
vC = 14'b0000010100101011; // vC= 1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000010100000001; // vC= 1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001101; // iC= 1101 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011101; // iC= 1117 
vC = 14'b0000010101111010; // vC= 1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110011; // iC= 1075 
vC = 14'b0000010101001001; // vC= 1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001110; // iC= 1166 
vC = 14'b0000010101010110; // vC= 1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101101; // iC= 1069 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110111; // iC= 1207 
vC = 14'b0000010100100111; // vC= 1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000001; // iC= 1089 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101100; // iC= 1068 
vC = 14'b0000010101001001; // vC= 1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001001; // iC= 1161 
vC = 14'b0000010101011100; // vC= 1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011100; // iC= 1116 
vC = 14'b0000010101110001; // vC= 1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010011; // iC= 1043 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001001; // iC= 1033 
vC = 14'b0000010111000001; // vC= 1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010111; // iC= 1111 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100000; // iC= 1056 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010110; // iC= 1046 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100100; // iC= 1124 
vC = 14'b0000010101101011; // vC= 1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100111; // iC= 1063 
vC = 14'b0000010110010000; // vC= 1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100101; // iC=  997 
vC = 14'b0000010110001101; // vC= 1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101101; // iC= 1005 
vC = 14'b0000010101001000; // vC= 1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111010; // iC= 1082 
vC = 14'b0000010101110101; // vC= 1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100001; // iC= 1057 
vC = 14'b0000010101101100; // vC= 1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001110; // iC= 1102 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010110; // iC= 1046 
vC = 14'b0000010101011000; // vC= 1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000000; // iC= 1088 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101010; // iC= 1002 
vC = 14'b0000010110100010; // vC= 1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111101; // iC= 1021 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111001; // iC= 1081 
vC = 14'b0000010111001010; // vC= 1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011010; // iC= 1050 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111111; // iC= 1087 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000001; // iC= 1025 
vC = 14'b0000010111010101; // vC= 1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100101; // iC=  997 
vC = 14'b0000010101101100; // vC= 1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110111; // iC=  951 
vC = 14'b0000010111100101; // vC= 1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011110; // iC=  926 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100011; // iC= 1059 
vC = 14'b0000010111100100; // vC= 1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011111; // iC=  927 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101100; // iC=  940 
vC = 14'b0000010110000100; // vC= 1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110101; // iC=  949 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010101; // iC=  981 
vC = 14'b0000010111111011; // vC= 1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110001; // iC= 1009 
vC = 14'b0000010111111000; // vC= 1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111110; // iC= 1022 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100111; // iC=  999 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101001; // iC= 1001 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000100; // iC=  964 
vC = 14'b0000010111010111; // vC= 1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011010; // iC=  922 
vC = 14'b0000010111100101; // vC= 1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001100; // iC=  972 
vC = 14'b0000010110100101; // vC= 1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010010; // iC=  914 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011000; // iC=  856 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010101; // iC=  917 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110000; // iC=  880 
vC = 14'b0000010111111001; // vC= 1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110110; // iC=  822 
vC = 14'b0000010110010110; // vC= 1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000001; // iC=  897 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100101; // iC=  805 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011010; // iC=  794 
vC = 14'b0000011000101111; // vC= 1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111111; // iC=  895 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101001; // iC=  873 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110101; // iC=  821 
vC = 14'b0000010111001111; // vC= 1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100010; // iC=  802 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001111; // iC=  847 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011010; // iC=  858 
vC = 14'b0000010110101010; // vC= 1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101011; // iC=  811 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100010; // iC=  866 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100001; // iC=  865 
vC = 14'b0000010110110100; // vC= 1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111010; // iC=  762 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011100; // iC=  860 
vC = 14'b0000010111101010; // vC= 1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010010; // iC=  850 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010001; // iC=  849 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110111; // iC=  823 
vC = 14'b0000011000011001; // vC= 1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010000; // iC=  784 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100100; // iC=  740 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000100; // iC=  836 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110101; // iC=  821 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000111; // iC=  775 
vC = 14'b0000010111110001; // vC= 1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100010; // iC=  738 
vC = 14'b0000010111111000; // vC= 1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001111; // iC=  783 
vC = 14'b0000010111010101; // vC= 1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001001; // iC=  777 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111001; // iC=  761 
vC = 14'b0000011001100110; // vC= 1638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110010; // iC=  690 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011111; // iC=  671 
vC = 14'b0000011001101001; // vC= 1641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101000; // iC=  744 
vC = 14'b0000011000111000; // vC= 1592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100000; // iC=  736 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001001; // iC=  713 
vC = 14'b0000011000110110; // vC= 1590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100010; // iC=  738 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100101; // iC=  741 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011100; // iC=  732 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001001; // iC=  649 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111111; // iC=  639 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001001; // iC=  649 
vC = 14'b0000011001101100; // vC= 1644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100001; // iC=  673 
vC = 14'b0000011001110000; // vC= 1648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010001; // iC=  721 
vC = 14'b0000011000110100; // vC= 1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111101; // iC=  637 
vC = 14'b0000011001110100; // vC= 1652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111100; // iC=  700 
vC = 14'b0000011001100100; // vC= 1636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111001; // iC=  697 
vC = 14'b0000011000101111; // vC= 1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000111; // iC=  647 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100100; // iC=  676 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000000; // iC=  640 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010100; // iC=  660 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101110; // iC=  622 
vC = 14'b0000011001100100; // vC= 1636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100000; // iC=  672 
vC = 14'b0000011001100100; // vC= 1636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010100; // iC=  532 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101011; // iC=  555 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111010; // iC=  570 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011011; // iC=  539 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101100; // iC=  556 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000010; // iC=  514 
vC = 14'b0000011001011010; // vC= 1626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110111; // iC=  567 
vC = 14'b0000011000101101; // vC= 1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111011; // iC=  635 
vC = 14'b0000011000101100; // vC= 1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101011; // iC=  491 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111111; // iC=  575 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010101; // iC=  597 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001111; // iC=  463 
vC = 14'b0000011010011000; // vC= 1688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001000; // iC=  456 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010000; // iC=  592 
vC = 14'b0000011001011010; // vC= 1626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111000; // iC=  504 
vC = 14'b0000011001111101; // vC= 1661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000101; // iC=  453 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001011; // iC=  459 
vC = 14'b0000011001101110; // vC= 1646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010110; // iC=  470 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001011; // iC=  459 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001111; // iC=  527 
vC = 14'b0000011001100011; // vC= 1635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010001; // iC=  465 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110111; // iC=  439 
vC = 14'b0000011010101100; // vC= 1708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110001; // iC=  433 
vC = 14'b0000011000110110; // vC= 1590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101101; // iC=  493 
vC = 14'b0000011001010010; // vC= 1618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101000; // iC=  488 
vC = 14'b0000011000010111; // vC= 1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100111; // iC=  359 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010111; // iC=  471 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101011; // iC=  363 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011111; // iC=  351 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100010; // iC=  418 
vC = 14'b0000011000110101; // vC= 1589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010111; // iC=  343 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010110; // iC=  278 
vC = 14'b0000011010000010; // vC= 1666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110111; // iC=  375 
vC = 14'b0000011010011110; // vC= 1694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001001; // iC=  329 
vC = 14'b0000011000110101; // vC= 1589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001111; // iC=  335 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010100; // iC=  340 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100101; // iC=  229 
vC = 14'b0000011001011100; // vC= 1628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000001; // iC=  321 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001000; // iC=  200 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011011; // iC=  283 
vC = 14'b0000011001011011; // vC= 1627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111010; // iC=  186 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100000; // iC=  160 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010000; // iC=  144 
vC = 14'b0000011010100100; // vC= 1700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011111; // iC=   95 
vC = 14'b0000011010111011; // vC= 1723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011000; // iC=   88 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010001; // iC=  209 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101111; // iC=  175 
vC = 14'b0000011010111100; // vC= 1724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011011; // iC=  155 
vC = 14'b0000011010001101; // vC= 1677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011011; // iC=   91 
vC = 14'b0000011010011101; // vC= 1693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101001; // iC=  105 
vC = 14'b0000011010001110; // vC= 1678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000111; // iC=    7 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010100; // iC=   20 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101001; // iC=   41 
vC = 14'b0000011001011100; // vC= 1628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011111; // iC=   31 
vC = 14'b0000011010001010; // vC= 1674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000011; // iC=  -61 
vC = 14'b0000011001100111; // vC= 1639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001100; // iC=  -52 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010111; // iC=  -41 
vC = 14'b0000011001000101; // vC= 1605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101100; // iC=  -84 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100111; // iC=  -89 
vC = 14'b0000011010001001; // vC= 1673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111000; // iC= -200 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001110; // iC= -178 
vC = 14'b0000011001011100; // vC= 1628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001010; // iC= -182 
vC = 14'b0000011001111101; // vC= 1661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001110; // iC= -242 
vC = 14'b0000011010010110; // vC= 1686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100001; // iC= -159 
vC = 14'b0000011010010000; // vC= 1680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010010; // iC= -174 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000111; // iC= -185 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110100; // iC= -268 
vC = 14'b0000011010000100; // vC= 1668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001001; // iC= -247 
vC = 14'b0000011010010101; // vC= 1685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111001; // iC= -263 
vC = 14'b0000011010010000; // vC= 1680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001001; // iC= -311 
vC = 14'b0000011001010110; // vC= 1622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111011; // iC= -325 
vC = 14'b0000011001100101; // vC= 1637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000011; // iC= -445 
vC = 14'b0000011001111001; // vC= 1657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111010; // iC= -390 
vC = 14'b0000011010001110; // vC= 1678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111111; // iC= -385 
vC = 14'b0000011010010011; // vC= 1683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111100; // iC= -452 
vC = 14'b0000011001110001; // vC= 1649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110011; // iC= -525 
vC = 14'b0000011001110010; // vC= 1650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000110; // iC= -506 
vC = 14'b0000011010000111; // vC= 1671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011101; // iC= -483 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001000; // iC= -568 
vC = 14'b0000011010001101; // vC= 1677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111011; // iC= -581 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001111; // iC= -561 
vC = 14'b0000011001111001; // vC= 1657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010100; // iC= -620 
vC = 14'b0000011001110100; // vC= 1652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110001; // iC= -719 
vC = 14'b0000011001000101; // vC= 1605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101100; // iC= -596 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110100; // iC= -716 
vC = 14'b0000011000101101; // vC= 1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011010; // iC= -678 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111111; // iC= -705 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111110; // iC= -706 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000111; // iC= -825 
vC = 14'b0000011000110100; // vC= 1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100101; // iC= -795 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100000; // iC= -864 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111101; // iC= -835 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101000; // iC= -856 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001010; // iC= -886 
vC = 14'b0000011000110100; // vC= 1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001010; // iC= -822 
vC = 14'b0000010111001001; // vC= 1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100011; // iC= -861 
vC = 14'b0000010111011011; // vC= 1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010111; // iC= -873 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011110; // iC= -930 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010101; // iC= -939 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101011; // iC= -917 
vC = 14'b0000011001000101; // vC= 1605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101100; // iC= -980 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011000; // iC=-1000 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111110; // iC=-1090 
vC = 14'b0000010110100000; // vC= 1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111001; // iC=-1031 
vC = 14'b0000010111000000; // vC= 1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101010; // iC=-1110 
vC = 14'b0000010111001011; // vC= 1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100010; // iC=-1118 
vC = 14'b0000010111010010; // vC= 1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101010; // iC=-1046 
vC = 14'b0000010111000001; // vC= 1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111010; // iC=-1158 
vC = 14'b0000010111011001; // vC= 1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001110; // iC=-1138 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101110; // iC=-1170 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110001; // iC=-1231 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001100; // iC=-1268 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111100; // iC=-1220 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111100; // iC=-1284 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b0000010111000010; // vC= 1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010111; // iC=-1193 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001000; // iC=-1208 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000000; // iC=-1344 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100000; // iC=-1312 
vC = 14'b0000010111100001; // vC= 1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100000; // iC=-1376 
vC = 14'b0000010110010111; // vC= 1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001101; // iC=-1331 
vC = 14'b0000010111010111; // vC= 1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101001; // iC=-1431 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101000; // iC=-1368 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101000; // iC=-1304 
vC = 14'b0000010101001000; // vC= 1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111001; // iC=-1351 
vC = 14'b0000010110011001; // vC= 1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111011; // iC=-1413 
vC = 14'b0000010110001111; // vC= 1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110011; // iC=-1357 
vC = 14'b0000010100110110; // vC= 1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b0000010110101101; // vC= 1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b0000010101010110; // vC= 1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001011; // iC=-1397 
vC = 14'b0000010101001101; // vC= 1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111100; // iC=-1476 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100110; // iC=-1562 
vC = 14'b0000010101000000; // vC= 1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101101; // iC=-1555 
vC = 14'b0000010100101100; // vC= 1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b0000010100011100; // vC= 1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b0000010011110010; // vC= 1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b0000010011110000; // vC= 1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001010; // iC=-1526 
vC = 14'b0000010100001110; // vC= 1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b0000010101100111; // vC= 1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010100; // iC=-1580 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b0000010100111001; // vC= 1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b0000010100001110; // vC= 1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000111; // iC=-1657 
vC = 14'b0000010100001101; // vC= 1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100011; // iC=-1629 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000010011111001; // vC= 1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b0000010100001110; // vC= 1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011110; // iC=-1634 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b0000010011110100; // vC= 1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101011; // iC=-1557 
vC = 14'b0000010010101110; // vC= 1198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000010011001101; // vC= 1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100100; // iC=-1692 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000111; // iC=-1657 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101101; // iC=-1619 
vC = 14'b0000010011100001; // vC= 1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110110; // iC=-1610 
vC = 14'b0000010010010100; // vC= 1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b0000010011111000; // vC= 1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b0000010010011110; // vC= 1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111001; // iC=-1607 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101101; // iC=-1619 
vC = 14'b0000010010100000; // vC= 1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100000; // iC=-1760 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011111; // iC=-1633 
vC = 14'b0000010001101101; // vC= 1133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b0000010010101011; // vC= 1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000010000100100; // vC= 1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b0000010010000101; // vC= 1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000010001010100; // vC= 1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100000; // iC=-1632 
vC = 14'b0000010000101110; // vC= 1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011001; // iC=-1639 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000010001000110; // vC= 1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101010; // iC=-1686 
vC = 14'b0000010000110000; // vC= 1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000010001111100; // vC= 1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000001111110010; // vC= 1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b0000010001100000; // vC= 1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000010000100110; // vC= 1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b0000001111101100; // vC= 1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b0000001111000010; // vC=  962 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b0000010000011010; // vC= 1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000001110111000; // vC=  952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000001111101100; // vC= 1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b0000001110111000; // vC=  952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000001111111011; // vC= 1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000001110001110; // vC=  910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000001110001100; // vC=  908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000001111110110; // vC= 1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000001111011111; // vC=  991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100000; // iC=-1760 
vC = 14'b0000001110001111; // vC=  911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000001111111110; // vC= 1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000001111010011; // vC=  979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000001111000101; // vC=  965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b0000001101111011; // vC=  891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b0000001110001010; // vC=  906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000001101101100; // vC=  876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000001110110100; // vC=  948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000001110000001; // vC=  897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b0000001100110001; // vC=  817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000001100100000; // vC=  800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000001110000110; // vC=  902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000001101011100; // vC=  860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000001101111000; // vC=  888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000001110011011; // vC=  923 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000001100100111; // vC=  807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000001101011111; // vC=  863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000001101001011; // vC=  843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000001011011111; // vC=  735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101111; // iC=-1873 
vC = 14'b0000001100110000; // vC=  816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b0000001100001110; // vC=  782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000001011001100; // vC=  716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001011101100; // vC=  748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110110; // iC=-1866 
vC = 14'b0000001101000001; // vC=  833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b0000001011110110; // vC=  758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000001011110010; // vC=  754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101001; // iC=-1879 
vC = 14'b0000001011001100; // vC=  716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000001011000001; // vC=  705 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000001011001101; // vC=  717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000001010011010; // vC=  666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000001010011000; // vC=  664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111111; // iC=-1857 
vC = 14'b0000001100000111; // vC=  775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000001010001010; // vC=  650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000011; // iC=-1853 
vC = 14'b0000001100001011; // vC=  779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111110; // iC=-1858 
vC = 14'b0000001011001011; // vC=  715 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000001011100111; // vC=  743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000001011010001; // vC=  721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000001001100111; // vC=  615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100010; // iC=-1886 
vC = 14'b0000001001011001; // vC=  601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000001011010011; // vC=  723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000001010100010; // vC=  674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110110; // iC=-1866 
vC = 14'b0000001001101110; // vC=  622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000001000101110; // vC=  558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101001; // iC=-1879 
vC = 14'b0000001010101010; // vC=  682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111111; // iC=-1857 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000001000011010; // vC=  538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b0000001001110000; // vC=  624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000001000001110; // vC=  526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000001000100111; // vC=  551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101110; // iC=-1874 
vC = 14'b0000001001010010; // vC=  594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100110; // iC=-1882 
vC = 14'b0000000111101000; // vC=  488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000000111101011; // vC=  491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001000001001; // vC=  521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110011; // iC=-1869 
vC = 14'b0000001000000010; // vC=  514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000001001000011; // vC=  579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b0000000111100110; // vC=  486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b0000000111101111; // vC=  495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101000; // iC=-1880 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000001000100000; // vC=  544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100010; // iC=-1886 
vC = 14'b0000000111010101; // vC=  469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000011; // iC=-1853 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010101; // iC=-1899 
vC = 14'b0000000110110100; // vC=  436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000000111001000; // vC=  456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011000; // iC=-1896 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101001; // iC=-1879 
vC = 14'b0000000110110100; // vC=  436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000000111111111; // vC=  511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000000111010101; // vC=  469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101011; // iC=-1877 
vC = 14'b0000000110111011; // vC=  443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000000111000000; // vC=  448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000000110110111; // vC=  439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111101; // iC=-1859 
vC = 14'b0000000101010100; // vC=  340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100001; // iC=-1887 
vC = 14'b0000000101111101; // vC=  381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000000110011011; // vC=  411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000000101111011; // vC=  379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000000110110000; // vC=  432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000000110111011; // vC=  443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b0000000100101011; // vC=  299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000000110101001; // vC=  425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010001011; // iC=-1909 
vC = 14'b0000000100011101; // vC=  285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000000100010110; // vC=  278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000000101111101; // vC=  381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111010; // iC=-1862 
vC = 14'b0000000011110101; // vC=  245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100100; // iC=-1820 
vC = 14'b0000000101101010; // vC=  362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000011; // iC=-1853 
vC = 14'b0000000101001110; // vC=  334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011000; // iC=-1896 
vC = 14'b0000000011111100; // vC=  252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000000100100100; // vC=  292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000000100110010; // vC=  306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100000; // iC=-1760 
vC = 14'b0000000101011011; // vC=  347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000000100011000; // vC=  280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011101; // iC=-1827 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000101000110; // vC=  326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000000101000000; // vC=  320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000000011111101; // vC=  253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000000011111010; // vC=  250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000000011011001; // vC=  217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011101; // iC=-1891 
vC = 14'b0000000010111011; // vC=  187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000100010011; // vC=  275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b0000000011010011; // vC=  211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100110; // iC=-1882 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011101; // iC=-1827 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101010; // iC=-1878 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011110; // iC=-1890 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000000010001111; // vC=  143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000000011101001; // vC=  233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000000001011111; // vC=   95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000000001010011; // vC=   83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000000001110101; // vC=  117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000000000100110; // vC=   38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000000; // iC=-1792 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000000010011000; // vC=  152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000000001000101; // vC=   69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000000000100101; // vC=   37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000000001011011; // vC=   91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b0000000000101000; // vC=   40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b0000000001111011; // vC=  123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010011; // iC=-1837 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b0000000000011010; // vC=   26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b1111111111010111; // vC=  -41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b1111111111010110; // vC=  -42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b1111111111100110; // vC=  -26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b1111111111001101; // vC=  -51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b1111111111011001; // vC=  -39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b1111111111010011; // vC=  -45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b1111111111101011; // vC=  -21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010000; // iC=-1840 
vC = 14'b1111111110101101; // vC=  -83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000000000001011; // vC=   11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000000000010111; // vC=   23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000000000101011; // vC=   43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000000000010111; // vC=   23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011110; // iC=-1698 
vC = 14'b1111111110010000; // vC= -112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b1111111110111100; // vC=  -68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b1111111111001101; // vC=  -51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b1111111101100110; // vC= -154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b1111111111100001; // vC=  -31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b1111111110101001; // vC=  -87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b1111111101011100; // vC= -164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b1111111101110111; // vC= -137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b1111111110110101; // vC=  -75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b1111111110001111; // vC= -113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b1111111110010110; // vC= -106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011101; // iC=-1827 
vC = 14'b1111111101110100; // vC= -140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b1111111101100000; // vC= -160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b1111111100111001; // vC= -199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110010; // iC=-1806 
vC = 14'b1111111101101011; // vC= -149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110001; // iC=-1679 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b1111111101100100; // vC= -156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b1111111110011100; // vC= -100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b1111111100001011; // vC= -245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b1111111101001001; // vC= -183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b1111111100010001; // vC= -239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b1111111101000001; // vC= -191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101010; // iC=-1686 
vC = 14'b1111111100110110; // vC= -202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b1111111101100110; // vC= -154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b1111111101000000; // vC= -192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b1111111100011011; // vC= -229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111100; // iC=-1668 
vC = 14'b1111111100100100; // vC= -220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b1111111101001001; // vC= -183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b1111111101010010; // vC= -174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b1111111100101011; // vC= -213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b1111111011110011; // vC= -269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b1111111011001010; // vC= -310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b1111111100010011; // vC= -237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100011; // iC=-1693 
vC = 14'b1111111011110010; // vC= -270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b1111111100011111; // vC= -225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b1111111010101010; // vC= -342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b1111111010001000; // vC= -376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b1111111010110111; // vC= -329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b1111111011000110; // vC= -314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101000; // iC=-1688 
vC = 14'b1111111011100001; // vC= -287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b1111111010010011; // vC= -365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b1111111010001001; // vC= -375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b1111111011101010; // vC= -278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b1111111011011100; // vC= -292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b1111111001011011; // vC= -421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111111; // iC=-1665 
vC = 14'b1111111001000111; // vC= -441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011000; // iC=-1704 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b1111111001100110; // vC= -410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b1111111011000001; // vC= -319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b1111111011000010; // vC= -318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110000; // iC=-1680 
vC = 14'b1111111010101001; // vC= -343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101000; // iC=-1688 
vC = 14'b1111111010000100; // vC= -380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b1111111010011011; // vC= -357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b1111111010100011; // vC= -349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b1111111001101001; // vC= -407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b1111111001111100; // vC= -388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b1111111001000101; // vC= -443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b1111111001000101; // vC= -443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b1111111001101101; // vC= -403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b1111111000110001; // vC= -463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011101; // iC=-1571 
vC = 14'b1111111000001011; // vC= -501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110000; // iC=-1680 
vC = 14'b1111111000001101; // vC= -499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b1111110111111111; // vC= -513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100110; // iC=-1562 
vC = 14'b1111110111010110; // vC= -554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110100; // iC=-1612 
vC = 14'b1111111000001000; // vC= -504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001100; // iC=-1588 
vC = 14'b1111111000001111; // vC= -497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b1111111000111100; // vC= -452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b1111111001000100; // vC= -444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b1111110110111011; // vC= -581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b1111110110111001; // vC= -583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100100; // iC=-1692 
vC = 14'b1111110111011001; // vC= -551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b1111111000101110; // vC= -466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b1111110110110100; // vC= -588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b1111110110110011; // vC= -589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b1111110110001110; // vC= -626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b1111110111110010; // vC= -526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b1111110101110000; // vC= -656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b1111110110100110; // vC= -602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010000; // iC=-1648 
vC = 14'b1111110111110111; // vC= -521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b1111110110010101; // vC= -619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b1111110111001001; // vC= -567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101101; // iC=-1555 
vC = 14'b1111110101100101; // vC= -667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011101; // iC=-1571 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111110; // iC=-1538 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b1111110101010001; // vC= -687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b1111110101111100; // vC= -644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b1111110101101010; // vC= -662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001000; // iC=-1464 
vC = 14'b1111110100101110; // vC= -722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000010; // iC=-1470 
vC = 14'b1111110100100110; // vC= -730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011111; // iC=-1505 
vC = 14'b1111110101110110; // vC= -650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b1111110110100101; // vC= -603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b1111110110100111; // vC= -601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b1111110101010000; // vC= -688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b1111110100001111; // vC= -753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011000; // iC=-1512 
vC = 14'b1111110100011110; // vC= -738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b1111110100011111; // vC= -737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110001; // iC=-1551 
vC = 14'b1111110100111100; // vC= -708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111010; // iC=-1478 
vC = 14'b1111110011110010; // vC= -782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111111; // iC=-1473 
vC = 14'b1111110011101011; // vC= -789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001110; // iC=-1458 
vC = 14'b1111110101100011; // vC= -669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011011; // iC=-1445 
vC = 14'b1111110011011101; // vC= -803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b1111110100010001; // vC= -751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001110; // iC=-1458 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101100; // iC=-1428 
vC = 14'b1111110011111011; // vC= -773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111011; // iC=-1413 
vC = 14'b1111110100010100; // vC= -748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111010; // iC=-1478 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b1111110100100000; // vC= -736 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111100; // iC=-1412 
vC = 14'b1111110011101011; // vC= -789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b1111110011100100; // vC= -796 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101011; // iC=-1493 
vC = 14'b1111110100110111; // vC= -713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111001; // iC=-1479 
vC = 14'b1111110100111000; // vC= -712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b1111110010101011; // vC= -853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000001; // iC=-1407 
vC = 14'b1111110011110011; // vC= -781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111101; // iC=-1411 
vC = 14'b1111110010001110; // vC= -882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010100; // iC=-1388 
vC = 14'b1111110011010110; // vC= -810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100100; // iC=-1436 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001101; // iC=-1459 
vC = 14'b1111110011101000; // vC= -792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100101; // iC=-1371 
vC = 14'b1111110010010110; // vC= -874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100011; // iC=-1373 
vC = 14'b1111110100001101; // vC= -755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111000; // iC=-1416 
vC = 14'b1111110100000110; // vC= -762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011011; // iC=-1381 
vC = 14'b1111110011110111; // vC= -777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111001; // iC=-1479 
vC = 14'b1111110001100001; // vC= -927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111011; // iC=-1413 
vC = 14'b1111110001001110; // vC= -946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000011; // iC=-1405 
vC = 14'b1111110010001111; // vC= -881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111000; // iC=-1352 
vC = 14'b1111110010101001; // vC= -855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b1111110001110100; // vC= -908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001100; // iC=-1332 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100011; // iC=-1309 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110101; // iC=-1419 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101011; // iC=-1301 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100110; // iC=-1434 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000001; // iC=-1407 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100110; // iC=-1306 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000000; // iC=-1280 
vC = 14'b1111110001100001; // vC= -927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000100; // iC=-1276 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011101; // iC=-1315 
vC = 14'b1111110000101000; // vC= -984 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101001; // iC=-1303 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010001; // iC=-1263 
vC = 14'b1111110000110100; // vC= -972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101100; // iC=-1364 
vC = 14'b1111110010000000; // vC= -896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011010; // iC=-1254 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101011; // iC=-1237 
vC = 14'b1111110000010101; // vC=-1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110011; // iC=-1357 
vC = 14'b1111110000101110; // vC= -978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001110; // iC=-1330 
vC = 14'b1111110000001001; // vC=-1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101100; // iC=-1300 
vC = 14'b1111110001000010; // vC= -958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101000; // iC=-1368 
vC = 14'b1111101111011000; // vC=-1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000010; // iC=-1278 
vC = 14'b1111110000010000; // vC=-1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111001; // iC=-1351 
vC = 14'b1111101111100001; // vC=-1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010100; // iC=-1260 
vC = 14'b1111110000111110; // vC= -962 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101001; // iC=-1239 
vC = 14'b1111101111101111; // vC=-1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100111; // iC=-1305 
vC = 14'b1111110000010011; // vC=-1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100110; // iC=-1242 
vC = 14'b1111101111000101; // vC=-1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110011; // iC=-1293 
vC = 14'b1111110000101110; // vC= -978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001100; // iC=-1332 
vC = 14'b1111110000001101; // vC=-1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111101; // iC=-1283 
vC = 14'b1111101110110101; // vC=-1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001001; // iC=-1271 
vC = 14'b1111110000101110; // vC= -978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110011; // iC=-1293 
vC = 14'b1111110000001000; // vC=-1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010000; // iC=-1200 
vC = 14'b1111101110101010; // vC=-1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011000; // iC=-1192 
vC = 14'b1111101110101001; // vC=-1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100011; // iC=-1245 
vC = 14'b1111101110100100; // vC=-1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001100; // iC=-1204 
vC = 14'b1111101111001101; // vC=-1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001000; // iC=-1208 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001011; // iC=-1141 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111110; // iC=-1218 
vC = 14'b1111110000100010; // vC= -990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101001; // iC=-1175 
vC = 14'b1111101111000000; // vC=-1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010111; // iC=-1129 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101000; // iC=-1176 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101001; // iC=-1175 
vC = 14'b1111101111101110; // vC=-1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100010; // iC=-1246 
vC = 14'b1111101111111011; // vC=-1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011101; // iC=-1251 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101110; // iC=-1234 
vC = 14'b1111101111001000; // vC=-1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010000; // iC=-1136 
vC = 14'b1111101110100000; // vC=-1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011000; // iC=-1192 
vC = 14'b1111101101100110; // vC=-1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000100; // iC=-1212 
vC = 14'b1111101111100000; // vC=-1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100111; // iC=-1177 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100010; // iC=-1118 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111001; // iC=-1095 
vC = 14'b1111101111101101; // vC=-1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010101; // iC=-1131 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001001; // iC=-1143 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010000; // iC=-1136 
vC = 14'b1111101101110110; // vC=-1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101010; // iC=-1110 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100100; // iC=-1116 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100101; // iC=-1179 
vC = 14'b1111101101000010; // vC=-1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010000; // iC=-1136 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011011; // iC=-1189 
vC = 14'b1111101110011110; // vC=-1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000111; // iC=-1145 
vC = 14'b1111101110001111; // vC=-1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100111; // iC=-1177 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010011; // iC=-1069 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001111; // iC=-1073 
vC = 14'b1111101110011011; // vC=-1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011110; // iC=-1122 
vC = 14'b1111101101000010; // vC=-1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010100; // iC=-1132 
vC = 14'b1111101110001101; // vC=-1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100011; // iC=-1117 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001001; // iC=-1079 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001000; // iC=-1144 
vC = 14'b1111101101100000; // vC=-1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010101; // iC=-1003 
vC = 14'b1111101110010111; // vC=-1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011010; // iC=-1062 
vC = 14'b1111101101000000; // vC=-1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011110; // iC=-1122 
vC = 14'b1111101100010001; // vC=-1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111111; // iC=-1025 
vC = 14'b1111101100110001; // vC=-1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111000; // iC=-1032 
vC = 14'b1111101101111011; // vC=-1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110100; // iC=-1036 
vC = 14'b1111101110001100; // vC=-1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000100; // iC= -956 
vC = 14'b1111101101100110; // vC=-1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101111; // iC= -977 
vC = 14'b1111101011110100; // vC=-1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010100; // iC=-1068 
vC = 14'b1111101100111100; // vC=-1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011000; // iC=-1064 
vC = 14'b1111101101001000; // vC=-1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011010; // iC=-1062 
vC = 14'b1111101011100010; // vC=-1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010100; // iC=-1068 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111011; // iC=-1029 
vC = 14'b1111101100001000; // vC=-1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011001; // iC= -935 
vC = 14'b1111101100111100; // vC=-1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111010; // iC=-1030 
vC = 14'b1111101100000111; // vC=-1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101000; // iC= -984 
vC = 14'b1111101011001110; // vC=-1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011110; // iC=-1058 
vC = 14'b1111101011101001; // vC=-1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011001; // iC= -935 
vC = 14'b1111101100011111; // vC=-1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001100; // iC=-1012 
vC = 14'b1111101011000010; // vC=-1342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101000; // iC= -984 
vC = 14'b1111101100101001; // vC=-1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100101; // iC= -923 
vC = 14'b1111101100101011; // vC=-1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010111; // iC= -873 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000110; // iC=-1018 
vC = 14'b1111101100001010; // vC=-1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011000; // iC=-1000 
vC = 14'b1111101011111101; // vC=-1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101011; // iC= -917 
vC = 14'b1111101010111011; // vC=-1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111101; // iC= -899 
vC = 14'b1111101100111000; // vC=-1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001111; // iC= -945 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100000; // iC= -992 
vC = 14'b1111101100110000; // vC=-1232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111100; // iC= -836 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011010; // iC= -870 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000011; // iC= -957 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110100; // iC= -972 
vC = 14'b1111101011111010; // vC=-1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011101; // iC= -867 
vC = 14'b1111101100101110; // vC=-1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100000; // iC= -864 
vC = 14'b1111101010010111; // vC=-1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000110; // iC= -826 
vC = 14'b1111101100010100; // vC=-1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010000; // iC= -816 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111110; // iC= -834 
vC = 14'b1111101010111110; // vC=-1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100111; // iC= -857 
vC = 14'b1111101010110111; // vC=-1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011101; // iC= -803 
vC = 14'b1111101100000001; // vC=-1279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100010; // iC= -798 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110110; // iC= -778 
vC = 14'b1111101010010000; // vC=-1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000000; // iC= -896 
vC = 14'b1111101011101111; // vC=-1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111010; // iC= -774 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010101; // iC= -811 
vC = 14'b1111101011111010; // vC=-1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100010; // iC= -798 
vC = 14'b1111101001101111; // vC=-1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001101; // iC= -883 
vC = 14'b1111101010111111; // vC=-1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000011; // iC= -893 
vC = 14'b1111101011110010; // vC=-1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100001; // iC= -735 
vC = 14'b1111101001110100; // vC=-1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101000; // iC= -728 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000010; // iC= -766 
vC = 14'b1111101010111011; // vC=-1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000011; // iC= -829 
vC = 14'b1111101001111011; // vC=-1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100100; // iC= -796 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111011; // iC= -837 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001001; // iC= -759 
vC = 14'b1111101010010000; // vC=-1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000100; // iC= -828 
vC = 14'b1111101011100011; // vC=-1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110001; // iC= -847 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000100; // iC= -700 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001001; // iC= -695 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010100; // iC= -748 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001001; // iC= -695 
vC = 14'b1111101001111101; // vC=-1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011100; // iC= -804 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000010; // iC= -766 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010110; // iC= -810 
vC = 14'b1111101010001001; // vC=-1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011000; // iC= -744 
vC = 14'b1111101010111010; // vC=-1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110100; // iC= -652 
vC = 14'b1111101010100100; // vC=-1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101111; // iC= -657 
vC = 14'b1111101010001010; // vC=-1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101100; // iC= -660 
vC = 14'b1111101001101100; // vC=-1428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100010; // iC= -734 
vC = 14'b1111101001001000; // vC=-1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000101; // iC= -635 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011110; // iC= -738 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010010; // iC= -686 
vC = 14'b1111101010110010; // vC=-1358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001101; // iC= -755 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101110; // iC= -658 
vC = 14'b1111101010110001; // vC=-1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111111; // iC= -641 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110000; // iC= -592 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100000; // iC= -672 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101101; // iC= -659 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000000; // iC= -704 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010001; // iC= -623 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001111; // iC= -561 
vC = 14'b1111101000100101; // vC=-1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101111; // iC= -657 
vC = 14'b1111101000111001; // vC=-1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010100; // iC= -556 
vC = 14'b1111101000010110; // vC=-1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100001; // iC= -671 
vC = 14'b1111101010101100; // vC=-1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110100; // iC= -588 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111111; // iC= -577 
vC = 14'b1111101001100111; // vC=-1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110110; // iC= -586 
vC = 14'b1111101010010001; // vC=-1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110001; // iC= -527 
vC = 14'b1111101000001111; // vC=-1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b1111101010011101; // vC=-1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011110; // iC= -546 
vC = 14'b1111101000011110; // vC=-1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000011; // iC= -637 
vC = 14'b1111101000111111; // vC=-1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010111; // iC= -553 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111010; // iC= -518 
vC = 14'b1111101001011111; // vC=-1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111110; // iC= -578 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111100; // iC= -516 
vC = 14'b1111101010001010; // vC=-1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101111; // iC= -593 
vC = 14'b1111101000010011; // vC=-1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111011; // iC= -517 
vC = 14'b1111101001111100; // vC=-1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011001; // iC= -551 
vC = 14'b1111101001000000; // vC=-1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001000; // iC= -504 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001011; // iC= -501 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000100; // iC= -444 
vC = 14'b1111101010001011; // vC=-1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100100; // iC= -540 
vC = 14'b1111101000010011; // vC=-1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001111; // iC= -561 
vC = 14'b1111101001111100; // vC=-1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111010; // iC= -518 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110110; // iC= -458 
vC = 14'b1111100111111111; // vC=-1537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101000; // iC= -536 
vC = 14'b1111100111100110; // vC=-1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111111; // iC= -513 
vC = 14'b1111101001001000; // vC=-1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010011; // iC= -429 
vC = 14'b1111100111111111; // vC=-1537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010000; // iC= -432 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101110; // iC= -466 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011110; // iC= -418 
vC = 14'b1111101000001111; // vC=-1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010111; // iC= -361 
vC = 14'b1111100111110011; // vC=-1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111110; // iC= -450 
vC = 14'b1111100111011110; // vC=-1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101010; // iC= -470 
vC = 14'b1111101000011011; // vC=-1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111101; // iC= -451 
vC = 14'b1111100111111010; // vC=-1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010010; // iC= -366 
vC = 14'b1111101001001101; // vC=-1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001110; // iC= -306 
vC = 14'b1111100111010100; // vC=-1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110100; // iC= -396 
vC = 14'b1111100111101001; // vC=-1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010011; // iC= -365 
vC = 14'b1111101000100010; // vC=-1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111100; // iC= -324 
vC = 14'b1111101001000011; // vC=-1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000001; // iC= -319 
vC = 14'b1111101001011110; // vC=-1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110000; // iC= -272 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010011; // iC= -237 
vC = 14'b1111100111011001; // vC=-1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111111; // iC= -257 
vC = 14'b1111101001101001; // vC=-1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111010; // iC= -262 
vC = 14'b1111100111100011; // vC=-1565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111010; // iC= -262 
vC = 14'b1111100111010101; // vC=-1579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101011; // iC= -149 
vC = 14'b1111101001100101; // vC=-1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011010; // iC= -166 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010110; // iC= -170 
vC = 14'b1111101000111010; // vC=-1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011011; // iC= -229 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001011; // iC= -181 
vC = 14'b1111101000001100; // vC=-1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010100; // iC= -172 
vC = 14'b1111100111100101; // vC=-1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011101; // iC=  -99 
vC = 14'b1111100111100001; // vC=-1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000101; // iC= -187 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111110; // iC= -130 
vC = 14'b1111101000111111; // vC=-1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110101; // iC= -139 
vC = 14'b1111101001011110; // vC=-1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111010; // iC=   -6 
vC = 14'b1111101000111001; // vC=-1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101100; // iC=  -20 
vC = 14'b1111101001000000; // vC=-1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101010; // iC=   42 
vC = 14'b1111100111111110; // vC=-1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001110; // iC=   14 
vC = 14'b1111101000011101; // vC=-1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010000; // iC=  -48 
vC = 14'b1111101000100111; // vC=-1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011110; // iC=  -34 
vC = 14'b1111101001100100; // vC=-1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100101; // iC=  -27 
vC = 14'b1111100111001111; // vC=-1585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111011; // iC=   59 
vC = 14'b1111101000111001; // vC=-1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001100; // iC=  140 
vC = 14'b1111101000011110; // vC=-1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011101; // iC=  157 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011000; // iC=   88 
vC = 14'b1111100111110000; // vC=-1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111100; // iC=  188 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101000; // iC=  232 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101111; // iC=  175 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001110; // iC=  270 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011110; // iC=  222 
vC = 14'b1111101000000000; // vC=-1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000100; // iC=  324 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010010; // iC=  274 
vC = 14'b1111100111110010; // vC=-1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011111; // iC=  287 
vC = 14'b1111100111010010; // vC=-1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011101; // iC=  349 
vC = 14'b1111101001011111; // vC=-1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011011; // iC=  347 
vC = 14'b1111101000110011; // vC=-1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101001; // iC=  297 
vC = 14'b1111100111010011; // vC=-1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100101; // iC=  421 
vC = 14'b1111100111110101; // vC=-1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010100; // iC=  468 
vC = 14'b1111100111100000; // vC=-1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011001; // iC=  473 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111001; // iC=  505 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101000; // iC=  424 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100111; // iC=  487 
vC = 14'b1111101001001110; // vC=-1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010110; // iC=  534 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111110; // iC=  574 
vC = 14'b1111100111101111; // vC=-1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110100; // iC=  564 
vC = 14'b1111101000000110; // vC=-1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100110; // iC=  614 
vC = 14'b1111101000010010; // vC=-1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011010; // iC=  602 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100101; // iC=  677 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110100; // iC=  692 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101011; // iC=  747 
vC = 14'b1111100111110110; // vC=-1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101101; // iC=  685 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010011; // iC=  723 
vC = 14'b1111101000110110; // vC=-1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100111; // iC=  743 
vC = 14'b1111101000000110; // vC=-1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011101; // iC=  861 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010110; // iC=  790 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010001; // iC=  913 
vC = 14'b1111101001000100; // vC=-1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011101; // iC=  861 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010100; // iC=  852 
vC = 14'b1111101010100101; // vC=-1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000110; // iC=  902 
vC = 14'b1111101010010101; // vC=-1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101101; // iC=  941 
vC = 14'b1111101000010000; // vC=-1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111000; // iC= 1016 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110010; // iC= 1010 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100100; // iC=  932 
vC = 14'b1111101001011110; // vC=-1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100010; // iC= 1058 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001010; // iC= 1098 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010111; // iC= 1111 
vC = 14'b1111101010000011; // vC=-1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010001; // iC= 1105 
vC = 14'b1111101010011010; // vC=-1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110001; // iC= 1137 
vC = 14'b1111101010010100; // vC=-1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000001; // iC= 1089 
vC = 14'b1111101011001010; // vC=-1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001010; // iC= 1162 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011001; // iC= 1177 
vC = 14'b1111101011010000; // vC=-1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000101; // iC= 1157 
vC = 14'b1111101001110100; // vC=-1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010101; // iC= 1173 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010011; // iC= 1235 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000011; // iC= 1155 
vC = 14'b1111101010110111; // vC=-1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011100; // iC= 1244 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100101; // iC= 1189 
vC = 14'b1111101011101111; // vC=-1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101111; // iC= 1327 
vC = 14'b1111101011110011; // vC=-1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110011; // iC= 1331 
vC = 14'b1111101011110101; // vC=-1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011010; // iC= 1370 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001000; // iC= 1288 
vC = 14'b1111101001100001; // vC=-1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011001; // iC= 1305 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001011; // iC= 1419 
vC = 14'b1111101001111111; // vC=-1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000110; // iC= 1414 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001111; // iC= 1487 
vC = 14'b1111101100001110; // vC=-1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110000; // iC= 1392 
vC = 14'b1111101010111010; // vC=-1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101010; // iC= 1514 
vC = 14'b1111101001111101; // vC=-1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011001; // iC= 1433 
vC = 14'b1111101100011001; // vC=-1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110001; // iC= 1393 
vC = 14'b1111101010010010; // vC=-1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000001; // iC= 1537 
vC = 14'b1111101011100100; // vC=-1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110111; // iC= 1463 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110110; // iC= 1462 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100011; // iC= 1507 
vC = 14'b1111101101000000; // vC=-1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011111; // iC= 1567 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010010; // iC= 1618 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101001; // iC= 1641 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000110; // iC= 1542 
vC = 14'b1111101011010111; // vC=-1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101111; // iC= 1647 
vC = 14'b1111101011100011; // vC=-1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101101; // iC= 1645 
vC = 14'b1111101100000111; // vC=-1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101110; // iC= 1710 
vC = 14'b1111101011010101; // vC=-1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000001; // iC= 1729 
vC = 14'b1111101100111000; // vC=-1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b1111101100101011; // vC=-1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011001; // iC= 1625 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111101101111100; // vC=-1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b1111101101010011; // vC=-1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b1111101101011111; // vC=-1185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b1111101101111001; // vC=-1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110010; // iC= 1778 
vC = 14'b1111101100101010; // vC=-1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001100; // iC= 1740 
vC = 14'b1111101101100101; // vC=-1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001110; // iC= 1742 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b1111101110011111; // vC=-1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b1111101101100101; // vC=-1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001111; // iC= 1871 
vC = 14'b1111101101100110; // vC=-1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101110; // iC= 1774 
vC = 14'b1111101110000111; // vC=-1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b1111101110111100; // vC=-1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111100; // iC= 1788 
vC = 14'b1111101111011111; // vC=-1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000101; // iC= 1861 
vC = 14'b1111101111000011; // vC=-1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b1111101101101100; // vC=-1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b1111101111110100; // vC=-1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b1111101110100111; // vC=-1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b1111101101101100; // vC=-1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110101; // iC= 1845 
vC = 14'b1111101111100100; // vC=-1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000010; // iC= 1858 
vC = 14'b1111101110011010; // vC=-1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b1111101110110000; // vC=-1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101001; // iC= 1833 
vC = 14'b1111101111000011; // vC=-1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b1111101111000101; // vC=-1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b1111110000000100; // vC=-1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b1111101110100001; // vC=-1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110000110100; // vC= -972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b1111101110111001; // vC=-1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b1111110000111111; // vC= -961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111110001100011; // vC= -925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111110000010011; // vC=-1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111110; // iC= 1982 
vC = 14'b1111110001101010; // vC= -918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111110001000000; // vC= -960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b1111101111111101; // vC=-1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111110000100001; // vC= -991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111110000001100; // vC=-1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110010; // iC= 1906 
vC = 14'b1111110000100010; // vC= -990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b1111110000100000; // vC= -992 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111110000100000; // vC= -992 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111110001110011; // vC= -909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001000; // iC= 1864 
vC = 14'b1111110010001000; // vC= -888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b1111110001101100; // vC= -916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111110001111001; // vC= -903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b1111110011101001; // vC= -791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100010; // iC= 2018 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111110001101100; // vC= -916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111110011110011; // vC= -781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111000; // iC= 2040 
vC = 14'b1111110011000110; // vC= -826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b1111110100010111; // vC= -745 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000000; // iC= 1984 
vC = 14'b1111110011000101; // vC= -827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111110100000110; // vC= -762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110100101110; // vC= -722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111110100100000; // vC= -736 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b1111110011001100; // vC= -820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000111; // iC= 2055 
vC = 14'b1111110100001100; // vC= -756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111110101011000; // vC= -680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b1111110011101110; // vC= -786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110011110111; // vC= -777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b1111110100101110; // vC= -722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b1111110101111000; // vC= -648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111110100000001; // vC= -767 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b1111110100000111; // vC= -761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111110101110001; // vC= -655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010100; // iC= 2068 
vC = 14'b1111110100101000; // vC= -728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111110100010111; // vC= -745 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111110101111001; // vC= -647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111110101011110; // vC= -674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011101; // iC= 2013 
vC = 14'b1111110110000000; // vC= -640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b1111110101011010; // vC= -678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001000; // iC= 2056 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110100; // iC= 1972 
vC = 14'b1111110101000010; // vC= -702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111110101110000; // vC= -656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011001; // iC= 2073 
vC = 14'b1111110101001011; // vC= -693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111110101111011; // vC= -645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100000; // iC= 2080 
vC = 14'b1111110101011110; // vC= -674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010111; // iC= 2071 
vC = 14'b1111110111101110; // vC= -530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b1111110111100000; // vC= -544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111000; // iC= 2040 
vC = 14'b1111110110110011; // vC= -589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b1111110110000011; // vC= -637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111110110010000; // vC= -624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b1111110110100011; // vC= -605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b1111110111011110; // vC= -546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100101; // iC= 2085 
vC = 14'b1111110111001101; // vC= -563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111110111001001; // vC= -567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111110111100001; // vC= -543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000010; // iC= 2050 
vC = 14'b1111111000100101; // vC= -475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111111000111001; // vC= -455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111110111100000; // vC= -544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011101; // iC= 2013 
vC = 14'b1111111000111000; // vC= -456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100101; // iC= 2021 
vC = 14'b1111110111101000; // vC= -536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010100; // iC= 2004 
vC = 14'b1111111001011001; // vC= -423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011010; // iC= 2074 
vC = 14'b1111111001000111; // vC= -441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111111000010100; // vC= -492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001111; // iC= 2063 
vC = 14'b1111111000101001; // vC= -471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111111000100100; // vC= -476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111111000111011; // vC= -453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000100; // iC= 2052 
vC = 14'b1111111000110010; // vC= -462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111111000000111; // vC= -505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111111; // iC= 2047 
vC = 14'b1111111000011110; // vC= -482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100110; // iC= 2086 
vC = 14'b1111111000111011; // vC= -453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100010; // iC= 2082 
vC = 14'b1111111001000010; // vC= -446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011011; // iC= 2075 
vC = 14'b1111111000111011; // vC= -453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111111001010010; // vC= -430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101011; // iC= 2027 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b1111111000111011; // vC= -453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001100; // iC= 2060 
vC = 14'b1111111011001011; // vC= -309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100111; // iC= 2087 
vC = 14'b1111111001010100; // vC= -428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111111010100011; // vC= -349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011100; // iC= 1948 
vC = 14'b1111111011010001; // vC= -303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111111011000110; // vC= -314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010100; // iC= 2068 
vC = 14'b1111111010110010; // vC= -334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111111011101111; // vC= -273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111111010011000; // vC= -360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b1111111011011100; // vC= -292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b1111111011011101; // vC= -291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100110; // iC= 2086 
vC = 14'b1111111011100011; // vC= -285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001110; // iC= 2062 
vC = 14'b1111111011101111; // vC= -273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111111010110011; // vC= -333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111111010011100; // vC= -356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111111100011111; // vC= -225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b1111111011100000; // vC= -288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111111100111100; // vC= -196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111011111011; // vC= -261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000101; // iC= 2053 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110010; // iC= 2034 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010000; // iC= 2064 
vC = 14'b1111111100100100; // vC= -220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111101001000; // vC= -184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111111101110010; // vC= -142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100101; // iC= 2021 
vC = 14'b1111111101001011; // vC= -181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111101011101; // vC= -163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111001; // iC= 2041 
vC = 14'b1111111011110010; // vC= -270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111111101011111; // vC= -161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b1111111101011010; // vC= -166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b1111111101011011; // vC= -165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000010; // iC= 2050 
vC = 14'b1111111110100111; // vC=  -89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b1111111101010001; // vC= -175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011100; // iC= 2076 
vC = 14'b1111111101001110; // vC= -178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010101; // iC= 2069 
vC = 14'b1111111100111001; // vC= -199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100010; // iC= 2018 
vC = 14'b1111111101000110; // vC= -186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000011; // iC= 2051 
vC = 14'b1111111111011010; // vC=  -38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111111110100100; // vC=  -92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111111111001110; // vC=  -50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b1111111111101110; // vC=  -18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b1111111110100001; // vC=  -95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b1111111110010100; // vC= -108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b1111111110111100; // vC=  -68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111001; // iC= 2041 
vC = 14'b0000000000001011; // vC=   11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b1111111111000110; // vC=  -58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b0000000000001110; // vC=   14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111111110011100; // vC= -100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000100; // iC= 2052 
vC = 14'b1111111110101001; // vC=  -87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111111111010101; // vC=  -43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b0000000000101001; // vC=   41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b1111111110111110; // vC=  -66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b1111111111100000; // vC=  -32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111100; // iC= 2044 
vC = 14'b1111111111101110; // vC=  -18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111111111101110; // vC=  -18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111111111011; // vC=   -5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b0000000001111000; // vC=  120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b0000000000101010; // vC=   42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000100; // iC= 1924 
vC = 14'b1111111111110000; // vC=  -16 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b0000000001010010; // vC=   82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b0000000001001001; // vC=   73 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b0000000010100101; // vC=  165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001010; // iC= 1994 
vC = 14'b0000000001001110; // vC=   78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b0000000001110101; // vC=  117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b0000000010101100; // vC=  172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b0000000011000110; // vC=  198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b0000000011010110; // vC=  214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b0000000010110001; // vC=  177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b0000000010000101; // vC=  133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b0000000010000110; // vC=  134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b0000000011101100; // vC=  236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b0000000011000000; // vC=  192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b0000000011011100; // vC=  220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001111; // iC= 1871 
vC = 14'b0000000100000110; // vC=  262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b0000000010100010; // vC=  162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b0000000011110011; // vC=  243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b0000000100011010; // vC=  282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b0000000011111011; // vC=  251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b0000000100000011; // vC=  259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b0000000100010010; // vC=  274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000000011111011; // vC=  251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b0000000101000100; // vC=  324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b0000000101001101; // vC=  333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000111; // iC= 1991 
vC = 14'b0000000101001110; // vC=  334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000000100101001; // vC=  297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b0000000011101001; // vC=  233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b0000000100100101; // vC=  293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b0000000100100011; // vC=  291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b0000000110011001; // vC=  409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b0000000100000011; // vC=  259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b0000000101010110; // vC=  342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b0000000110101101; // vC=  429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b0000000100100100; // vC=  292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b0000000110011000; // vC=  408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b0000000110011001; // vC=  409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b0000000111000001; // vC=  449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b0000000111000111; // vC=  455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b0000000110010000; // vC=  400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b0000000101001010; // vC=  330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b0000000101100011; // vC=  355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b0000000111000111; // vC=  455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000000110111110; // vC=  446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b0000000110100101; // vC=  421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b0000000110111101; // vC=  445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010000; // iC= 1808 
vC = 14'b0000000111111100; // vC=  508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b0000001000000010; // vC=  514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000110; // iC= 1798 
vC = 14'b0000000110111011; // vC=  443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010001; // iC= 1873 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b0000001000000011; // vC=  515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b0000000110101111; // vC=  431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b0000000111010101; // vC=  469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100011; // iC= 1827 
vC = 14'b0000001000011010; // vC=  538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b0000000111101100; // vC=  492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000010; // iC= 1794 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111011; // iC= 1851 
vC = 14'b0000001000100111; // vC=  551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000010; // iC= 1794 
vC = 14'b0000001000101111; // vC=  559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000010; // iC= 1858 
vC = 14'b0000001000000100; // vC=  516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111001; // iC= 1849 
vC = 14'b0000000111110010; // vC=  498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b0000001000001100; // vC=  524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000001000010010; // vC=  530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b0000001001010110; // vC=  598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110110; // iC= 1846 
vC = 14'b0000001001010011; // vC=  595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000001000001110; // vC=  526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b0000001001110101; // vC=  629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b0000001001001101; // vC=  589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111000; // iC= 1720 
vC = 14'b0000001000010010; // vC=  530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b0000001001011110; // vC=  606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b0000001000010010; // vC=  530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100010; // iC= 1826 
vC = 14'b0000001010100111; // vC=  679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101101; // iC= 1709 
vC = 14'b0000001010110010; // vC=  690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b0000001001010011; // vC=  595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b0000001001100100; // vC=  612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b0000001001011110; // vC=  606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b0000001001111000; // vC=  632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001100; // iC= 1804 
vC = 14'b0000001011001111; // vC=  719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b0000001001011101; // vC=  605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000011; // iC= 1795 
vC = 14'b0000001010101010; // vC=  682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b0000001001011010; // vC=  602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b0000001010101010; // vC=  682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000001011110101; // vC=  757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b0000001011011010; // vC=  730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001110; // iC= 1678 
vC = 14'b0000001011110100; // vC=  756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110101; // iC= 1781 
vC = 14'b0000001011101100; // vC=  748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b0000001010001001; // vC=  649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001000; // iC= 1672 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b0000001011111001; // vC=  761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000110; // iC= 1670 
vC = 14'b0000001100011111; // vC=  799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110100; // iC= 1652 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101110; // iC= 1646 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111100; // iC= 1788 
vC = 14'b0000001100100011; // vC=  803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101101; // iC= 1709 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b0000001100011101; // vC=  797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011110; // iC= 1630 
vC = 14'b0000001100001100; // vC=  780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101001; // iC= 1641 
vC = 14'b0000001011001101; // vC=  717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100110; // iC= 1766 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000001; // iC= 1665 
vC = 14'b0000001011010001; // vC=  721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110111; // iC= 1655 
vC = 14'b0000001100010111; // vC=  791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b0000001100010111; // vC=  791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111100; // iC= 1596 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b0000001011111110; // vC=  766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b0000001101111111; // vC=  895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b0000001100011110; // vC=  798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001100000001; // vC=  769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b0000001110000011; // vC=  899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101011; // iC= 1579 
vC = 14'b0000001101101100; // vC=  876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b0000001110000001; // vC=  897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b0000001101111101; // vC=  893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b0000001100111111; // vC=  831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111100; // iC= 1596 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010010; // iC= 1618 
vC = 14'b0000001100011011; // vC=  795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011111; // iC= 1695 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110100; // iC= 1652 
vC = 14'b0000001110010110; // vC=  918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010010; // iC= 1554 
vC = 14'b0000001110010000; // vC=  912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111011; // iC= 1659 
vC = 14'b0000001110000110; // vC=  902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b0000001110010101; // vC=  917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001101000101; // vC=  837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001110101111; // vC=  943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111000; // iC= 1528 
vC = 14'b0000001101110100; // vC=  884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110111; // iC= 1527 
vC = 14'b0000001110010001; // vC=  913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011011; // iC= 1499 
vC = 14'b0000001110001110; // vC=  910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100111; // iC= 1639 
vC = 14'b0000001110111100; // vC=  956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010100; // iC= 1492 
vC = 14'b0000001111101001; // vC= 1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110101; // iC= 1525 
vC = 14'b0000001111010010; // vC=  978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110111; // iC= 1591 
vC = 14'b0000001111100110; // vC=  998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010110; // iC= 1494 
vC = 14'b0000001110010010; // vC=  914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101010; // iC= 1514 
vC = 14'b0000001110111111; // vC=  959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001110; // iC= 1486 
vC = 14'b0000001111011000; // vC=  984 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000010; // iC= 1474 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001110; // iC= 1550 
vC = 14'b0000001111011000; // vC=  984 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110101; // iC= 1525 
vC = 14'b0000001111000001; // vC=  961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000110; // iC= 1542 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010100; // iC= 1492 
vC = 14'b0000001111110110; // vC= 1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100110; // iC= 1446 
vC = 14'b0000010000110110; // vC= 1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010110; // iC= 1494 
vC = 14'b0000010000100011; // vC= 1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110001; // iC= 1457 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010011; // iC= 1555 
vC = 14'b0000001111001001; // vC=  969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010101; // iC= 1429 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001111; // iC= 1423 
vC = 14'b0000010000011010; // vC= 1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000010; // iC= 1538 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000010; // iC= 1538 
vC = 14'b0000001111000001; // vC=  961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001110; // iC= 1422 
vC = 14'b0000010001011111; // vC= 1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110110; // iC= 1462 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011111; // iC= 1503 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111110; // iC= 1406 
vC = 14'b0000001111101101; // vC= 1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000010; // iC= 1474 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011001; // iC= 1497 
vC = 14'b0000010001111111; // vC= 1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001110; // iC= 1486 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101110; // iC= 1390 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100100; // iC= 1444 
vC = 14'b0000010010001001; // vC= 1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000111; // iC= 1479 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000110; // iC= 1414 
vC = 14'b0000010010000011; // vC= 1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100101; // iC= 1445 
vC = 14'b0000010010010011; // vC= 1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111110; // iC= 1470 
vC = 14'b0000010010100001; // vC= 1185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001010; // iC= 1418 
vC = 14'b0000010010001101; // vC= 1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100111; // iC= 1383 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000000; // iC= 1472 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000100; // iC= 1476 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000100; // iC= 1412 
vC = 14'b0000010010110011; // vC= 1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001111; // iC= 1423 
vC = 14'b0000010010000001; // vC= 1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010000; // iC= 1424 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111110; // iC= 1406 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100010; // iC= 1314 
vC = 14'b0000010010001011; // vC= 1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001100; // iC= 1356 
vC = 14'b0000010001101101; // vC= 1133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011000; // iC= 1432 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000111; // iC= 1415 
vC = 14'b0000010001100000; // vC= 1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000100; // iC= 1412 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100100; // iC= 1380 
vC = 14'b0000010010101111; // vC= 1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010001; // iC= 1425 
vC = 14'b0000010011000100; // vC= 1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110101; // iC= 1333 
vC = 14'b0000010011011001; // vC= 1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101010; // iC= 1322 
vC = 14'b0000010011101100; // vC= 1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001101; // iC= 1357 
vC = 14'b0000010010111111; // vC= 1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111110; // iC= 1342 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111000; // iC= 1336 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010100; // iC= 1300 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011110; // iC= 1246 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110101; // iC= 1269 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111100; // iC= 1276 
vC = 14'b0000010011101010; // vC= 1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000000; // iC= 1344 
vC = 14'b0000010011101001; // vC= 1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100100; // iC= 1252 
vC = 14'b0000010010000010; // vC= 1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011100; // iC= 1244 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111101; // iC= 1277 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001010; // iC= 1290 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100111; // iC= 1255 
vC = 14'b0000010100000101; // vC= 1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100101; // iC= 1253 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110111; // iC= 1207 
vC = 14'b0000010100100100; // vC= 1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111000; // iC= 1336 
vC = 14'b0000010011100111; // vC= 1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110110; // iC= 1206 
vC = 14'b0000010100111101; // vC= 1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001000; // iC= 1224 
vC = 14'b0000010100101010; // vC= 1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110011; // iC= 1331 
vC = 14'b0000010100000111; // vC= 1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001110; // iC= 1294 
vC = 14'b0000010100011101; // vC= 1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011111; // iC= 1247 
vC = 14'b0000010101000011; // vC= 1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001000; // iC= 1224 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010000; // iC= 1168 
vC = 14'b0000010100010110; // vC= 1302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011010; // iC= 1306 
vC = 14'b0000010101001010; // vC= 1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110110; // iC= 1206 
vC = 14'b0000010101010100; // vC= 1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000001; // iC= 1217 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110001; // iC= 1137 
vC = 14'b0000010100010000; // vC= 1296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000011; // iC= 1155 
vC = 14'b0000010011001110; // vC= 1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101110; // iC= 1262 
vC = 14'b0000010101101011; // vC= 1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111100; // iC= 1148 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010010; // iC= 1234 
vC = 14'b0000010100101101; // vC= 1325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110000; // iC= 1136 
vC = 14'b0000010011010110; // vC= 1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010001; // iC= 1169 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110001; // iC= 1137 
vC = 14'b0000010101101010; // vC= 1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011010; // iC= 1242 
vC = 14'b0000010011101100; // vC= 1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b0000010100101010; // vC= 1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000110; // iC= 1222 
vC = 14'b0000010100001110; // vC= 1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000000; // iC= 1088 
vC = 14'b0000010100111010; // vC= 1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011100; // iC= 1116 
vC = 14'b0000010101010011; // vC= 1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000010011110010; // vC= 1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000011; // iC= 1155 
vC = 14'b0000010100000111; // vC= 1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000010011110111; // vC= 1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111011; // iC= 1211 
vC = 14'b0000010101101010; // vC= 1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010100; // iC= 1044 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110001; // iC= 1201 
vC = 14'b0000010110000101; // vC= 1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011100; // iC= 1052 
vC = 14'b0000010110011110; // vC= 1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111001; // iC= 1081 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011101; // iC= 1117 
vC = 14'b0000010101111011; // vC= 1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011101; // iC= 1053 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001101; // iC= 1037 
vC = 14'b0000010110001010; // vC= 1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010001; // iC= 1041 
vC = 14'b0000010101111000; // vC= 1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010010; // iC= 1042 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111110; // iC= 1150 
vC = 14'b0000010101110101; // vC= 1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100110; // iC=  998 
vC = 14'b0000010101000011; // vC= 1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110100; // iC= 1140 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101100; // iC= 1004 
vC = 14'b0000010100111010; // vC= 1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110111; // iC= 1079 
vC = 14'b0000010100111111; // vC= 1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111011; // iC= 1019 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101101; // iC= 1069 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110111; // iC= 1079 
vC = 14'b0000010101000100; // vC= 1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001100; // iC= 1036 
vC = 14'b0000010110111000; // vC= 1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011100; // iC=  988 
vC = 14'b0000010111010000; // vC= 1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011001; // iC=  985 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011001; // iC=  985 
vC = 14'b0000010101100101; // vC= 1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001011; // iC= 1035 
vC = 14'b0000010110010011; // vC= 1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000011; // iC=  963 
vC = 14'b0000010111011001; // vC= 1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110011; // iC=  947 
vC = 14'b0000010111101010; // vC= 1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001100; // iC=  972 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010010; // iC=  978 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011101; // iC=  989 
vC = 14'b0000010110000010; // vC= 1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011110; // iC=  990 
vC = 14'b0000010110100101; // vC= 1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100100; // iC=  932 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010100; // iC=  916 
vC = 14'b0000010110010000; // vC= 1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101010; // iC= 1002 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001100; // iC=  972 
vC = 14'b0000010111100100; // vC= 1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101101; // iC=  941 
vC = 14'b0000010110110000; // vC= 1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010001; // iC=  977 
vC = 14'b0000010111000010; // vC= 1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100000; // iC=  928 
vC = 14'b0000010111100111; // vC= 1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010010; // iC=  914 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001111; // iC=  911 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010000; // iC=  976 
vC = 14'b0000010110110110; // vC= 1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010011; // iC=  979 
vC = 14'b0000010111011110; // vC= 1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010110; // iC=  918 
vC = 14'b0000010111001000; // vC= 1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100010; // iC=  866 
vC = 14'b0000010111000011; // vC= 1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010001; // iC=  977 
vC = 14'b0000010111011011; // vC= 1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110011; // iC=  883 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010011; // iC=  851 
vC = 14'b0000010111001101; // vC= 1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101100; // iC=  940 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110111; // iC=  887 
vC = 14'b0000010110110111; // vC= 1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100000; // iC=  864 
vC = 14'b0000010110001110; // vC= 1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110001; // iC=  945 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010011; // iC=  851 
vC = 14'b0000010111001110; // vC= 1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111000; // iC=  824 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000010; // iC=  834 
vC = 14'b0000011000101011; // vC= 1579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111100; // iC=  892 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001001; // iC=  905 
vC = 14'b0000010111001010; // vC= 1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111011; // iC=  891 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000010; // iC=  898 
vC = 14'b0000010111100100; // vC= 1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001111; // iC=  847 
vC = 14'b0000010111010010; // vC= 1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111011; // iC=  891 
vC = 14'b0000010111100111; // vC= 1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110100; // iC=  756 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110010; // iC=  818 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101111; // iC=  879 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100110; // iC=  806 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011101; // iC=  861 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000011; // iC=  707 
vC = 14'b0000010111100101; // vC= 1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000010; // iC=  834 
vC = 14'b0000011000010011; // vC= 1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100100; // iC=  740 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110100; // iC=  692 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100001; // iC=  801 
vC = 14'b0000010110111001; // vC= 1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010100; // iC=  788 
vC = 14'b0000010111000010; // vC= 1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110101; // iC=  757 
vC = 14'b0000011001001101; // vC= 1613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100010; // iC=  674 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100111; // iC=  807 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001001; // iC=  649 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010101; // iC=  789 
vC = 14'b0000010111101011; // vC= 1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001110; // iC=  718 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000000; // iC=  640 
vC = 14'b0000011000110001; // vC= 1585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010000; // iC=  656 
vC = 14'b0000011000110110; // vC= 1590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000001; // iC=  769 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010000; // iC=  656 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110010; // iC=  690 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010010; // iC=  722 
vC = 14'b0000011001100111; // vC= 1639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000001; // iC=  641 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011101; // iC=  605 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011100; // iC=  668 
vC = 14'b0000011001001100; // vC= 1612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011111; // iC=  671 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001110; // iC=  590 
vC = 14'b0000011001001110; // vC= 1614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100010; // iC=  674 
vC = 14'b0000010111110111; // vC= 1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001110; // iC=  654 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000110; // iC=  646 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110001; // iC=  561 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111010; // iC=  698 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010011; // iC=  659 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001100; // iC=  588 
vC = 14'b0000010111110011; // vC= 1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110100; // iC=  628 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111000; // iC=  568 
vC = 14'b0000011001000101; // vC= 1605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111110; // iC=  574 
vC = 14'b0000010111111000; // vC= 1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101000; // iC=  552 
vC = 14'b0000011010001001; // vC= 1673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100100; // iC=  612 
vC = 14'b0000011001111100; // vC= 1660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110001; // iC=  497 
vC = 14'b0000011001010110; // vC= 1622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011010; // iC=  538 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000100; // iC=  516 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100001; // iC=  481 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110100; // iC=  500 
vC = 14'b0000011001010001; // vC= 1617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000011; // iC=  579 
vC = 14'b0000011001010110; // vC= 1622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001110; // iC=  462 
vC = 14'b0000011001101110; // vC= 1646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100011; // iC=  547 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101110; // iC=  494 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001000; // iC=  456 
vC = 14'b0000011000110001; // vC= 1585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011111; // iC=  479 
vC = 14'b0000011001000110; // vC= 1606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101111; // iC=  559 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110100; // iC=  564 
vC = 14'b0000011010011001; // vC= 1689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000100; // iC=  580 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100111; // iC=  423 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001000; // iC=  520 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010001; // iC=  401 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001001; // iC=  457 
vC = 14'b0000011001000110; // vC= 1606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110011; // iC=  435 
vC = 14'b0000011001111101; // vC= 1661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110000; // iC=  432 
vC = 14'b0000011001011011; // vC= 1627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000010; // iC=  514 
vC = 14'b0000011010010111; // vC= 1687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000001; // iC=  449 
vC = 14'b0000011001001110; // vC= 1614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000000; // iC=  384 
vC = 14'b0000011010000101; // vC= 1669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110011; // iC=  435 
vC = 14'b0000011010100000; // vC= 1696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111101; // iC=  317 
vC = 14'b0000011001101110; // vC= 1646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010011; // iC=  339 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010101; // iC=  405 
vC = 14'b0000011001111100; // vC= 1660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101011; // iC=  427 
vC = 14'b0000011010010011; // vC= 1683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011101; // iC=  413 
vC = 14'b0000011010001001; // vC= 1673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000101; // iC=  261 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001000; // iC=  392 
vC = 14'b0000011001000110; // vC= 1606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110001; // iC=  241 
vC = 14'b0000011010100010; // vC= 1698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010010; // iC=  338 
vC = 14'b0000011010011110; // vC= 1694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011101; // iC=  349 
vC = 14'b0000011010011011; // vC= 1691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010001; // iC=  209 
vC = 14'b0000011000101010; // vC= 1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100111; // iC=  167 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010011; // iC=  147 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000111; // iC=  263 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100000; // iC=  160 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010100; // iC=  148 
vC = 14'b0000011001000110; // vC= 1606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000011; // iC=  131 
vC = 14'b0000011000111101; // vC= 1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001100; // iC=  204 
vC = 14'b0000011010100111; // vC= 1703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000001; // iC=  129 
vC = 14'b0000011010011100; // vC= 1692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000111; // iC=  199 
vC = 14'b0000011010010101; // vC= 1685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011100; // iC=  156 
vC = 14'b0000011010011100; // vC= 1692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000111; // iC=   71 
vC = 14'b0000011001111011; // vC= 1659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010011; // iC=  147 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101100; // iC=   44 
vC = 14'b0000011000011101; // vC= 1565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000111; // iC=   71 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010110; // iC=   22 
vC = 14'b0000011001101010; // vC= 1642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101101; // iC=  -19 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000000; // iC=   64 
vC = 14'b0000011010011111; // vC= 1695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111101; // iC=   -3 
vC = 14'b0000011001011011; // vC= 1627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111001; // iC= -135 
vC = 14'b0000011010010111; // vC= 1687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111001; // iC=   -7 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101111; // iC= -145 
vC = 14'b0000011000101011; // vC= 1579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010101; // iC= -107 
vC = 14'b0000011000001001; // vC= 1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111011; // iC=  -69 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001110; // iC= -242 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000001; // iC= -127 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110000; // iC= -208 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011001; // iC= -231 
vC = 14'b0000011010010011; // vC= 1683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001110; // iC= -306 
vC = 14'b0000011001100101; // vC= 1637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111110; // iC= -194 
vC = 14'b0000011001101000; // vC= 1640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110010; // iC= -270 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101101; // iC= -275 
vC = 14'b0000011010011100; // vC= 1692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001101; // iC= -371 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100100; // iC= -348 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111110; // iC= -322 
vC = 14'b0000011010001001; // vC= 1673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100100; // iC= -412 
vC = 14'b0000011010000110; // vC= 1670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000110; // iC= -442 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000110; // iC= -442 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100000; // iC= -544 
vC = 14'b0000011001011101; // vC= 1629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000101; // iC= -507 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001011; // iC= -565 
vC = 14'b0000011001000101; // vC= 1605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101101; // iC= -595 
vC = 14'b0000010111111110; // vC= 1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001000; // iC= -504 
vC = 14'b0000010111111001; // vC= 1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011010; // iC= -614 
vC = 14'b0000011001110011; // vC= 1651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010111; // iC= -617 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000011; // iC= -701 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010001; // iC= -623 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011101; // iC= -739 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111111; // iC= -641 
vC = 14'b0000011000011101; // vC= 1565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011101; // iC= -739 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010101; // iC= -683 
vC = 14'b0000010111110101; // vC= 1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001101; // iC= -691 
vC = 14'b0000011001101001; // vC= 1641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011011; // iC= -741 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100100; // iC= -860 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011001; // iC= -807 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101110; // iC= -850 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100101; // iC= -923 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011110; // iC= -802 
vC = 14'b0000010111000100; // vC= 1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111111; // iC= -961 
vC = 14'b0000010111100100; // vC= 1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100010; // iC= -862 
vC = 14'b0000011001001110; // vC= 1614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010110; // iC= -874 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111010; // iC= -902 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101010; // iC= -918 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001000; // iC=-1080 
vC = 14'b0000010110111110; // vC= 1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110101; // iC=-1099 
vC = 14'b0000010110011000; // vC= 1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110100; // iC= -972 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111111; // iC=-1153 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100001; // iC=-1119 
vC = 14'b0000010110110100; // vC= 1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011111; // iC=-1185 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b0000010110101001; // vC= 1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110101; // iC=-1099 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011100; // iC=-1188 
vC = 14'b0000010110001000; // vC= 1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001001; // iC=-1207 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000001; // iC=-1151 
vC = 14'b0000010111001000; // vC= 1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100100; // iC=-1180 
vC = 14'b0000010111101100; // vC= 1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101001; // iC=-1239 
vC = 14'b0000010101100010; // vC= 1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110010; // iC=-1230 
vC = 14'b0000010111100101; // vC= 1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b0000010111011100; // vC= 1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111111; // iC=-1345 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101000; // iC=-1304 
vC = 14'b0000010111000001; // vC= 1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b0000010111010110; // vC= 1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011111; // iC=-1313 
vC = 14'b0000010101011010; // vC= 1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b0000010101101111; // vC= 1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010100; // iC=-1260 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001111; // iC=-1393 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b0000010101010101; // vC= 1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011110; // iC=-1378 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011000; // iC=-1320 
vC = 14'b0000010100101011; // vC= 1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110100; // iC=-1420 
vC = 14'b0000010101010010; // vC= 1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011111; // iC=-1377 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100011; // iC=-1437 
vC = 14'b0000010100001111; // vC= 1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010010; // iC=-1454 
vC = 14'b0000010101111100; // vC= 1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000110; // iC=-1402 
vC = 14'b0000010110010001; // vC= 1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b0000010100011000; // vC= 1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b0000010110011011; // vC= 1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000111; // iC=-1529 
vC = 14'b0000010101110101; // vC= 1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b0000010100101110; // vC= 1326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b0000010100111000; // vC= 1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b0000010100011101; // vC= 1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110100; // iC=-1548 
vC = 14'b0000010011110000; // vC= 1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b0000010100101100; // vC= 1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b0000010100100011; // vC= 1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000010011110111; // vC= 1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010010; // iC=-1582 
vC = 14'b0000010101001101; // vC= 1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101101; // iC=-1555 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000010011111101; // vC= 1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b0000010011011000; // vC= 1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110110; // iC=-1674 
vC = 14'b0000010100100000; // vC= 1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010001; // iC=-1583 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b0000010011111011; // vC= 1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b0000010010110010; // vC= 1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100110; // iC=-1562 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111101; // iC=-1603 
vC = 14'b0000010001110111; // vC= 1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011000; // iC=-1704 
vC = 14'b0000010010110001; // vC= 1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101101; // iC=-1619 
vC = 14'b0000010001110010; // vC= 1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010011; // iC=-1581 
vC = 14'b0000010010111000; // vC= 1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011100; // iC=-1636 
vC = 14'b0000010010100010; // vC= 1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101001; // iC=-1623 
vC = 14'b0000010001000010; // vC= 1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000010000111010; // vC= 1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b0000010000101100; // vC= 1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b0000010001100000; // vC= 1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b0000010000111100; // vC= 1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b0000010000010111; // vC= 1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b0000010001010011; // vC= 1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000010000010000; // vC= 1040 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000001111110011; // vC= 1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011101; // iC=-1699 
vC = 14'b0000010001011111; // vC= 1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b0000001111100101; // vC=  997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110110; // iC=-1674 
vC = 14'b0000001111111000; // vC= 1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101000; // iC=-1688 
vC = 14'b0000010000011010; // vC= 1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001101; // iC=-1651 
vC = 14'b0000001110111110; // vC=  958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000010000110101; // vC= 1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b0000010000100000; // vC= 1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000001111100001; // vC=  993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110111; // iC=-1673 
vC = 14'b0000001110100111; // vC=  935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b0000010000101000; // vC= 1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001111011000; // vC=  984 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000001111100001; // vC=  993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b0000001111110110; // vC= 1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b0000001111010000; // vC=  976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000001111000100; // vC=  964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110111; // iC=-1673 
vC = 14'b0000001111100011; // vC=  995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b0000001101100101; // vC=  869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000001101110010; // vC=  882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000001111001111; // vC=  975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110011; // iC=-1741 
vC = 14'b0000001101101110; // vC=  878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000001111011111; // vC=  991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000001111010001; // vC=  977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001101010000; // vC=  848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b0000001110110000; // vC=  944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110000; // iC=-1680 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b0000001100100000; // vC=  800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000001110101011; // vC=  939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000001101011100; // vC=  860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000001101110001; // vC=  881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001101011110; // vC=  862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000001100010101; // vC=  789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000001100001000; // vC=  776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001011; // iC=-1845 
vC = 14'b0000001011110111; // vC=  759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000001101100101; // vC=  869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000001011011100; // vC=  732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000001011011100; // vC=  732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100000; // iC=-1760 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b0000001011110100; // vC=  756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000001100001000; // vC=  776 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000001101001000; // vC=  840 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000001101001101; // vC=  845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000001011011100; // vC=  732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000001100000011; // vC=  771 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010011; // iC=-1837 
vC = 14'b0000001010011011; // vC=  667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b0000001100011001; // vC=  793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000001100101011; // vC=  811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000001011101011; // vC=  747 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111100; // iC=-1860 
vC = 14'b0000001010110011; // vC=  691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000001100001101; // vC=  781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000001010010011; // vC=  659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110010; // iC=-1806 
vC = 14'b0000001011110111; // vC=  759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b0000001010100111; // vC=  679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000001010010001; // vC=  657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000001001101001; // vC=  617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000001001010001; // vC=  593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110011; // iC=-1741 
vC = 14'b0000001011001001; // vC=  713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100000; // iC=-1760 
vC = 14'b0000001001001101; // vC=  589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000001010110010; // vC=  690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000001011000110; // vC=  710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000001010101111; // vC=  687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010000; // iC=-1840 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000001000100100; // vC=  548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010011; // iC=-1837 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111011; // iC=-1797 
vC = 14'b0000001001101101; // vC=  621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000001010101011; // vC=  683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000001000111111; // vC=  575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000001000001000; // vC=  520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000001000000101; // vC=  517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000001010000000; // vC=  640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111011; // iC=-1861 
vC = 14'b0000001001001110; // vC=  590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000001000011001; // vC=  537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110010; // iC=-1870 
vC = 14'b0000001001111000; // vC=  632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b0000001000101100; // vC=  556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000001000011010; // vC=  538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000000111101111; // vC=  495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000001001011100; // vC=  604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b0000001000101011; // vC=  555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000001000001100; // vC=  524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110001; // iC=-1871 
vC = 14'b0000001000101000; // vC=  552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000001000101100; // vC=  556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000111; // iC=-1849 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000001000110010; // vC=  562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000000111101010; // vC=  490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b0000000110100101; // vC=  421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000000111000000; // vC=  448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000000111100011; // vC=  483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000000110000100; // vC=  388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000010; // iC=-1854 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b0000000101011101; // vC=  349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000000101100101; // vC=  357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000000110011000; // vC=  408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000000110110100; // vC=  436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000000101000100; // vC=  324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000000101111110; // vC=  382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000000110101111; // vC=  431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001111; // iC=-1841 
vC = 14'b0000000101011000; // vC=  344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000000101001100; // vC=  332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000000110110001; // vC=  433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000000100101111; // vC=  303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000101000001; // vC=  321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000000110011111; // vC=  415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000000110011010; // vC=  410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000000101111001; // vC=  377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111101; // iC=-1859 
vC = 14'b0000000101011011; // vC=  347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100111; // iC=-1881 
vC = 14'b0000000100001010; // vC=  266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000000011111111; // vC=  255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011110; // iC=-1890 
vC = 14'b0000000011111110; // vC=  254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000000100101010; // vC=  298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000000011101111; // vC=  239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000000011111010; // vC=  250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110001; // iC=-1871 
vC = 14'b0000000011001111; // vC=  207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100000; // iC=-1888 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b0000000011011100; // vC=  220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000100000100; // vC=  260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000000010111000; // vC=  184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000000100001110; // vC=  270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000000011101010; // vC=  234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000000100100001; // vC=  289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000000011110011; // vC=  243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000000011100100; // vC=  228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000000011100101; // vC=  229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b0000000010010110; // vC=  150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001011; // iC=-1845 
vC = 14'b0000000100000011; // vC=  259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110110; // iC=-1866 
vC = 14'b0000000001111010; // vC=  122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000000011011100; // vC=  220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000000010011101; // vC=  157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b0000000001101001; // vC=  105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111011; // iC=-1797 
vC = 14'b0000000000011100; // vC=   28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000000010010011; // vC=  147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b0000000001010110; // vC=   86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010000; // iC=-1840 
vC = 14'b0000000000101010; // vC=   42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001110; // iC=-1842 
vC = 14'b0000000001110100; // vC=  116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b1111111111110111; // vC=   -9 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b0000000001011101; // vC=   93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b1111111111101011; // vC=  -21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b1111111111011000; // vC=  -40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000000001010010; // vC=   82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000000000100100; // vC=   36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010000; // iC=-1840 
vC = 14'b0000000000011011; // vC=   27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000000000011001; // vC=   25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001110; // iC=-1842 
vC = 14'b0000000000001011; // vC=   11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000000000100001; // vC=   33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b1111111111000111; // vC=  -57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b1111111111010011; // vC=  -45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b1111111111000010; // vC=  -62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000000; // iC=-1792 
vC = 14'b1111111110111111; // vC=  -65 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b1111111111101000; // vC=  -24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b1111111111111100; // vC=   -4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b1111111111101110; // vC=  -18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b1111111110010000; // vC= -112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b1111111101100010; // vC= -158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b1111111110010001; // vC= -111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b1111111110111011; // vC=  -69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b1111111111010010; // vC=  -46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b1111111101011010; // vC= -166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101000; // iC=-1688 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111010; // iC=-1798 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b1111111100110011; // vC= -205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b1111111111001011; // vC=  -53 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b1111111101001111; // vC= -177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b1111111100100111; // vC= -217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b1111111110001110; // vC= -114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b1111111110001101; // vC= -115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b1111111101101001; // vC= -151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b1111111110011010; // vC= -102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011101; // iC=-1699 
vC = 14'b1111111100100011; // vC= -221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111100; // iC=-1668 
vC = 14'b1111111100000110; // vC= -250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b1111111101010111; // vC= -169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000100; // iC=-1724 
vC = 14'b1111111101100011; // vC= -157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b1111111101011111; // vC= -161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b1111111101001010; // vC= -182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b1111111011101010; // vC= -278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b1111111011100111; // vC= -281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b1111111011001101; // vC= -307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b1111111011011000; // vC= -296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b1111111100011101; // vC= -227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010000; // iC=-1648 
vC = 14'b1111111010101100; // vC= -340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b1111111100011010; // vC= -230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010010; // iC=-1646 
vC = 14'b1111111011010100; // vC= -300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b1111111010101100; // vC= -340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101011; // iC=-1621 
vC = 14'b1111111010100101; // vC= -347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b1111111011110001; // vC= -271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100011; // iC=-1629 
vC = 14'b1111111010001011; // vC= -373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b1111111010000101; // vC= -379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b1111111011101000; // vC= -280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b1111111010111010; // vC= -326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b1111111011000111; // vC= -313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b1111111010010101; // vC= -363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b1111111010111111; // vC= -321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000001; // iC=-1663 
vC = 14'b1111111010010011; // vC= -365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100100; // iC=-1692 
vC = 14'b1111111010010001; // vC= -367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b1111111001001000; // vC= -440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100011; // iC=-1629 
vC = 14'b1111111000111111; // vC= -449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b1111111000111000; // vC= -456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b1111111001000011; // vC= -445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011001; // iC=-1639 
vC = 14'b1111111010110000; // vC= -336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b1111111001101111; // vC= -401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010000; // iC=-1648 
vC = 14'b1111111001100000; // vC= -416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111001; // iC=-1607 
vC = 14'b1111111000011101; // vC= -483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b1111111001010100; // vC= -428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b1111111000010101; // vC= -491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b1111111000111000; // vC= -456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b1111111000000101; // vC= -507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b1111111000001111; // vC= -497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b1111111001011000; // vC= -424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b1111111010001100; // vC= -372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b1111111001001100; // vC= -436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101101; // iC=-1619 
vC = 14'b1111111000100101; // vC= -475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b1111111010000000; // vC= -384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100101; // iC=-1691 
vC = 14'b1111111000010000; // vC= -496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110110; // iC=-1610 
vC = 14'b1111111000111110; // vC= -450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b1111111000100000; // vC= -480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b1111111000001101; // vC= -499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110001; // iC=-1551 
vC = 14'b1111110111100101; // vC= -539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100100; // iC=-1628 
vC = 14'b1111111000001100; // vC= -500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010001; // iC=-1583 
vC = 14'b1111110111011100; // vC= -548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111001; // iC=-1607 
vC = 14'b1111111000000000; // vC= -512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100000; // iC=-1632 
vC = 14'b1111110111001100; // vC= -564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001100; // iC=-1588 
vC = 14'b1111111000110110; // vC= -458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100100; // iC=-1564 
vC = 14'b1111111000000010; // vC= -510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111111; // iC=-1665 
vC = 14'b1111110110011111; // vC= -609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b1111111000011010; // vC= -486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111001; // iC=-1607 
vC = 14'b1111110110100000; // vC= -608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111100; // iC=-1540 
vC = 14'b1111111000011010; // vC= -486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b1111110111001110; // vC= -562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b1111110110110101; // vC= -587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b1111111000001110; // vC= -498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011101; // iC=-1507 
vC = 14'b1111110111010110; // vC= -554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100011; // iC=-1565 
vC = 14'b1111110111101010; // vC= -534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101101; // iC=-1555 
vC = 14'b1111110111000110; // vC= -570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b1111110101111111; // vC= -641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000111; // iC=-1529 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b1111110110110010; // vC= -590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b1111110101011100; // vC= -676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b1111110111010011; // vC= -557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010010; // iC=-1582 
vC = 14'b1111110111000101; // vC= -571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b1111110110000010; // vC= -638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b1111110110100110; // vC= -602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100110; // iC=-1562 
vC = 14'b1111110101000001; // vC= -703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b1111110101010000; // vC= -688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b1111110100101010; // vC= -726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b1111110101100110; // vC= -666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b1111110110100101; // vC= -603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b1111110100010100; // vC= -748 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110000; // iC=-1552 
vC = 14'b1111110101111100; // vC= -644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101011; // iC=-1429 
vC = 14'b1111110110001000; // vC= -632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b1111110101010000; // vC= -688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b1111110011111010; // vC= -774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b1111110100110011; // vC= -717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b1111110101101011; // vC= -661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010111; // iC=-1513 
vC = 14'b1111110100101100; // vC= -724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101111; // iC=-1553 
vC = 14'b1111110100010001; // vC= -751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b1111110100001110; // vC= -754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010101; // iC=-1451 
vC = 14'b1111110101110010; // vC= -654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b1111110011111110; // vC= -770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b1111110011110001; // vC= -783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110110; // iC=-1418 
vC = 14'b1111110101011000; // vC= -680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001100; // iC=-1524 
vC = 14'b1111110011110111; // vC= -777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b1111110011100111; // vC= -793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010010; // iC=-1390 
vC = 14'b1111110011001011; // vC= -821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000001; // iC=-1407 
vC = 14'b1111110100110101; // vC= -715 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111110011001100; // vC= -820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011000; // iC=-1448 
vC = 14'b1111110011000110; // vC= -826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110111; // iC=-1481 
vC = 14'b1111110011010110; // vC= -810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110001; // iC=-1359 
vC = 14'b1111110011011101; // vC= -803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111011; // iC=-1413 
vC = 14'b1111110010011111; // vC= -865 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011111; // iC=-1441 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001110; // iC=-1458 
vC = 14'b1111110010001110; // vC= -882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001010; // iC=-1398 
vC = 14'b1111110100000101; // vC= -763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111111; // iC=-1473 
vC = 14'b1111110010011110; // vC= -866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b1111110011000011; // vC= -829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b1111110011001100; // vC= -820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010101; // iC=-1323 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110100; // iC=-1356 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011111; // iC=-1377 
vC = 14'b1111110011001100; // vC= -820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011100; // iC=-1444 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b1111110011001100; // vC= -820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110101; // iC=-1419 
vC = 14'b1111110010101110; // vC= -850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111000; // iC=-1416 
vC = 14'b1111110011000101; // vC= -827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100010; // iC=-1374 
vC = 14'b1111110010101000; // vC= -856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010111; // iC=-1385 
vC = 14'b1111110001111110; // vC= -898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b1111110010001100; // vC= -884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010010; // iC=-1390 
vC = 14'b1111110000101001; // vC= -983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101001; // iC=-1303 
vC = 14'b1111110001011101; // vC= -931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111111; // iC=-1345 
vC = 14'b1111110010011001; // vC= -871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000011; // iC=-1341 
vC = 14'b1111110001111100; // vC= -900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b1111110001111101; // vC= -899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101101; // iC=-1299 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000010; // iC=-1278 
vC = 14'b1111110000001000; // vC=-1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100000; // iC=-1376 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110011; // iC=-1357 
vC = 14'b1111110001111101; // vC= -899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101001; // iC=-1303 
vC = 14'b1111110010000001; // vC= -895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101000; // iC=-1368 
vC = 14'b1111110000011111; // vC= -993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110001; // iC=-1295 
vC = 14'b1111110001110100; // vC= -908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101000; // iC=-1368 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110010; // iC=-1294 
vC = 14'b1111110001010110; // vC= -938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000000; // iC=-1344 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110100; // iC=-1228 
vC = 14'b1111101111101011; // vC=-1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111101111110001; // vC=-1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110101; // iC=-1355 
vC = 14'b1111110000100010; // vC= -990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010010; // iC=-1198 
vC = 14'b1111110000011000; // vC=-1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010101; // iC=-1323 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000111; // iC=-1273 
vC = 14'b1111101111100010; // vC=-1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b1111110000111101; // vC= -963 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000100; // iC=-1212 
vC = 14'b1111110001011100; // vC= -932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111101; // iC=-1219 
vC = 14'b1111110000001111; // vC=-1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101110; // iC=-1170 
vC = 14'b1111101111101001; // vC=-1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100110; // iC=-1242 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110111; // iC=-1289 
vC = 14'b1111101110110001; // vC=-1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111111; // iC=-1217 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101001; // iC=-1175 
vC = 14'b1111101111101010; // vC=-1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100100; // iC=-1244 
vC = 14'b1111101111011100; // vC=-1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b1111101111011111; // vC=-1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101101; // iC=-1171 
vC = 14'b1111101110110100; // vC=-1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110110; // iC=-1226 
vC = 14'b1111110000100001; // vC= -991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001101; // iC=-1139 
vC = 14'b1111101111000100; // vC=-1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011001; // iC=-1191 
vC = 14'b1111101111001111; // vC=-1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101010; // iC=-1238 
vC = 14'b1111101110011011; // vC=-1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011101; // iC=-1187 
vC = 14'b1111101110101111; // vC=-1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010110; // iC=-1258 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100100; // iC=-1244 
vC = 14'b1111101110100110; // vC=-1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011010; // iC=-1190 
vC = 14'b1111101111101000; // vC=-1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010000; // iC=-1136 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111000; // iC=-1096 
vC = 14'b1111101110010010; // vC=-1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000100; // iC=-1212 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000110; // iC=-1082 
vC = 14'b1111101110001101; // vC=-1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100110; // iC=-1178 
vC = 14'b1111101110110111; // vC=-1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111111; // iC=-1217 
vC = 14'b1111101110111001; // vC=-1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000111; // iC=-1209 
vC = 14'b1111101111000101; // vC=-1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011100; // iC=-1188 
vC = 14'b1111101111000011; // vC=-1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111011; // iC=-1157 
vC = 14'b1111101101101101; // vC=-1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100011; // iC=-1181 
vC = 14'b1111101110111000; // vC=-1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001010; // iC=-1206 
vC = 14'b1111101110110001; // vC=-1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000010; // iC=-1086 
vC = 14'b1111101111010111; // vC=-1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111110; // iC=-1154 
vC = 14'b1111101101111000; // vC=-1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100111; // iC=-1177 
vC = 14'b1111101110011010; // vC=-1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101100; // iC=-1108 
vC = 14'b1111101101010010; // vC=-1198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011000; // iC=-1128 
vC = 14'b1111101101101111; // vC=-1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001001; // iC=-1079 
vC = 14'b1111101110101101; // vC=-1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010111; // iC=-1065 
vC = 14'b1111101110100101; // vC=-1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000100; // iC=-1020 
vC = 14'b1111101110101100; // vC=-1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111111; // iC=-1153 
vC = 14'b1111101110111000; // vC=-1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010010; // iC=-1006 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100111; // iC=-1113 
vC = 14'b1111101101100011; // vC=-1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100000; // iC=-1120 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100100; // iC= -988 
vC = 14'b1111101101111000; // vC=-1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001001; // iC=-1079 
vC = 14'b1111101101110011; // vC=-1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110010; // iC=-1102 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011100; // iC=-1124 
vC = 14'b1111101100101000; // vC=-1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110000; // iC= -976 
vC = 14'b1111101100101110; // vC=-1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000010; // iC=-1022 
vC = 14'b1111101100000011; // vC=-1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000010; // iC=-1022 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001010; // iC=-1078 
vC = 14'b1111101100000101; // vC=-1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100001; // iC=-1055 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100111; // iC=-1049 
vC = 14'b1111101101000101; // vC=-1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111101101100011; // vC=-1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111000; // iC= -968 
vC = 14'b1111101011110101; // vC=-1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011111; // iC= -929 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100010; // iC=-1054 
vC = 14'b1111101011100101; // vC=-1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101110; // iC=-1042 
vC = 14'b1111101101000011; // vC=-1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001101; // iC= -947 
vC = 14'b1111101100011011; // vC=-1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111000; // iC= -904 
vC = 14'b1111101101000000; // vC=-1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011011; // iC= -997 
vC = 14'b1111101101011000; // vC=-1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001100; // iC=-1012 
vC = 14'b1111101100101100; // vC=-1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001010; // iC= -886 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010000; // iC= -944 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010011; // iC= -877 
vC = 14'b1111101100011011; // vC=-1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010001; // iC=-1007 
vC = 14'b1111101100101100; // vC=-1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000001; // iC=-1023 
vC = 14'b1111101101010000; // vC=-1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110101; // iC= -971 
vC = 14'b1111101011011011; // vC=-1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000011; // iC= -893 
vC = 14'b1111101100111100; // vC=-1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000100; // iC= -892 
vC = 14'b1111101011111011; // vC=-1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001000; // iC= -888 
vC = 14'b1111101100110011; // vC=-1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010111; // iC= -873 
vC = 14'b1111101100111000; // vC=-1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011000; // iC= -936 
vC = 14'b1111101100111000; // vC=-1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111000; // iC= -904 
vC = 14'b1111101010110011; // vC=-1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111111; // iC= -961 
vC = 14'b1111101100111101; // vC=-1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111111; // iC= -897 
vC = 14'b1111101010101010; // vC=-1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101101; // iC= -915 
vC = 14'b1111101100111101; // vC=-1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110100; // iC= -908 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010010; // iC= -814 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100101; // iC= -859 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100101; // iC= -795 
vC = 14'b1111101011011100; // vC=-1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010111; // iC= -809 
vC = 14'b1111101011001111; // vC=-1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010100; // iC= -876 
vC = 14'b1111101010110001; // vC=-1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111101011111110; // vC=-1282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010111; // iC= -809 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100011; // iC= -861 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111110; // iC= -770 
vC = 14'b1111101011100111; // vC=-1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111011; // iC= -773 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110001; // iC= -783 
vC = 14'b1111101100001110; // vC=-1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001110; // iC= -818 
vC = 14'b1111101011001001; // vC=-1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101000; // iC= -792 
vC = 14'b1111101010101111; // vC=-1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101001; // iC= -855 
vC = 14'b1111101010100111; // vC=-1369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000111; // iC= -825 
vC = 14'b1111101011011000; // vC=-1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001011; // iC= -821 
vC = 14'b1111101011010111; // vC=-1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001000; // iC= -824 
vC = 14'b1111101001101110; // vC=-1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110001; // iC= -719 
vC = 14'b1111101010011101; // vC=-1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110000; // iC= -720 
vC = 14'b1111101010000010; // vC=-1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101011; // iC= -725 
vC = 14'b1111101010000000; // vC=-1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111101011001001; // vC=-1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001100; // iC= -820 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111101; // iC= -707 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000000; // iC= -704 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010110; // iC= -746 
vC = 14'b1111101001101110; // vC=-1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010100; // iC= -812 
vC = 14'b1111101011101001; // vC=-1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100010; // iC= -798 
vC = 14'b1111101011011100; // vC=-1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010011; // iC= -685 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010001; // iC= -687 
vC = 14'b1111101001001000; // vC=-1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110101; // iC= -651 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001111; // iC= -753 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101100; // iC= -788 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100111; // iC= -729 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011010; // iC= -678 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010001; // iC= -751 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010100; // iC= -684 
vC = 14'b1111101010100101; // vC=-1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110101; // iC= -651 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010111; // iC= -745 
vC = 14'b1111101011001101; // vC=-1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111010; // iC= -646 
vC = 14'b1111101010110111; // vC=-1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111010; // iC= -710 
vC = 14'b1111101010111110; // vC=-1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110100; // iC= -716 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000010; // iC= -702 
vC = 14'b1111101010010100; // vC=-1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100100; // iC= -732 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110111; // iC= -585 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001101; // iC= -627 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110111; // iC= -713 
vC = 14'b1111101000101111; // vC=-1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011000; // iC= -552 
vC = 14'b1111101010110011; // vC=-1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010100; // iC= -684 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101100; // iC= -596 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010011; // iC= -621 
vC = 14'b1111101010010101; // vC=-1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101110; // iC= -530 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010111; // iC= -617 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110111; // iC= -521 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111010; // iC= -646 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010001; // iC= -559 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110111; // iC= -585 
vC = 14'b1111101001000100; // vC=-1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000101; // iC= -507 
vC = 14'b1111101000010000; // vC=-1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001101; // iC= -499 
vC = 14'b1111101001101001; // vC=-1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011011; // iC= -485 
vC = 14'b1111101000110011; // vC=-1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001010; // iC= -502 
vC = 14'b1111101010100001; // vC=-1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111100; // iC= -516 
vC = 14'b1111101000100101; // vC=-1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011110; // iC= -546 
vC = 14'b1111101001010001; // vC=-1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000000; // iC= -512 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000110; // iC= -506 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001010; // iC= -502 
vC = 14'b1111101000111100; // vC=-1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100110; // iC= -538 
vC = 14'b1111101010010010; // vC=-1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100001; // iC= -543 
vC = 14'b1111101000101111; // vC=-1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100111; // iC= -537 
vC = 14'b1111100111110001; // vC=-1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100110; // iC= -538 
vC = 14'b1111101001100111; // vC=-1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011001; // iC= -551 
vC = 14'b1111101000001000; // vC=-1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001011; // iC= -565 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111101; // iC= -451 
vC = 14'b1111101001000110; // vC=-1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000010; // iC= -446 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011001; // iC= -487 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111000; // iC= -392 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000100; // iC= -508 
vC = 14'b1111101001011111; // vC=-1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000001; // iC= -383 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000001; // iC= -447 
vC = 14'b1111100111110100; // vC=-1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000000; // iC= -448 
vC = 14'b1111101000110011; // vC=-1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010001; // iC= -431 
vC = 14'b1111101001000110; // vC=-1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101101; // iC= -467 
vC = 14'b1111101001111011; // vC=-1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110011; // iC= -397 
vC = 14'b1111101000100110; // vC=-1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001010; // iC= -374 
vC = 14'b1111101000001011; // vC=-1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111011; // iC= -325 
vC = 14'b1111101001001111; // vC=-1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011011; // iC= -421 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111000; // iC= -328 
vC = 14'b1111101000000010; // vC=-1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000000; // iC= -384 
vC = 14'b1111101000001110; // vC=-1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101111; // iC= -273 
vC = 14'b1111100111110111; // vC=-1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111001; // iC= -263 
vC = 14'b1111101001101001; // vC=-1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010110; // iC= -234 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000010; // iC= -254 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100010; // iC= -222 
vC = 14'b1111101001101100; // vC=-1428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111001; // iC= -199 
vC = 14'b1111100111110011; // vC=-1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011001; // iC= -167 
vC = 14'b1111100111100011; // vC=-1565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101111; // iC= -273 
vC = 14'b1111100111111001; // vC=-1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000111; // iC= -185 
vC = 14'b1111101000100110; // vC=-1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110101; // iC= -203 
vC = 14'b1111101001001101; // vC=-1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011101; // iC=  -99 
vC = 14'b1111101000000011; // vC=-1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011100; // iC= -164 
vC = 14'b1111100111101001; // vC=-1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101010; // iC=  -86 
vC = 14'b1111100111100001; // vC=-1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000010; // iC= -190 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011110; // iC= -162 
vC = 14'b1111100111010001; // vC=-1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000001; // iC= -127 
vC = 14'b1111101000000111; // vC=-1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011001; // iC= -103 
vC = 14'b1111101000010111; // vC=-1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111010010; // iC=  -46 
vC = 14'b1111100111111001; // vC=-1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101001; // iC=  -23 
vC = 14'b1111101000110110; // vC=-1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010010; // iC= -110 
vC = 14'b1111101000010000; // vC=-1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000100; // iC=   68 
vC = 14'b1111100111101000; // vC=-1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010111; // iC=   87 
vC = 14'b1111100111100010; // vC=-1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100010; // iC=   98 
vC = 14'b1111100111100101; // vC=-1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000110; // iC=   70 
vC = 14'b1111101000000111; // vC=-1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000000; // iC=   64 
vC = 14'b1111101000010011; // vC=-1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001001; // iC=  137 
vC = 14'b1111100111100000; // vC=-1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001110; // iC=  142 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101010; // iC=  170 
vC = 14'b1111101000010100; // vC=-1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110101; // iC=  181 
vC = 14'b1111101001101000; // vC=-1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001101; // iC=  141 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011000; // iC=  216 
vC = 14'b1111101000010001; // vC=-1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000101; // iC=  197 
vC = 14'b1111101000010000; // vC=-1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010110; // iC=  278 
vC = 14'b1111101000000110; // vC=-1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000100; // iC=  196 
vC = 14'b1111101000001101; // vC=-1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011000; // iC=  280 
vC = 14'b1111101000010101; // vC=-1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000010; // iC=  386 
vC = 14'b1111101000000110; // vC=-1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011111; // iC=  287 
vC = 14'b1111101001011111; // vC=-1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001001; // iC=  329 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000101; // iC=  389 
vC = 14'b1111101001110101; // vC=-1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000011; // iC=  323 
vC = 14'b1111101001010100; // vC=-1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011111; // iC=  351 
vC = 14'b1111100111101001; // vC=-1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101011; // iC=  427 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010010; // iC=  530 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100010; // iC=  482 
vC = 14'b1111101000111111; // vC=-1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010000; // iC=  592 
vC = 14'b1111101001111100; // vC=-1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111111; // iC=  511 
vC = 14'b1111101000001001; // vC=-1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001011; // iC=  523 
vC = 14'b1111101000000110; // vC=-1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111000; // iC=  568 
vC = 14'b1111101000001100; // vC=-1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010010; // iC=  594 
vC = 14'b1111101000011011; // vC=-1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000010; // iC=  578 
vC = 14'b1111101000111001; // vC=-1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000011; // iC=  707 
vC = 14'b1111100111101111; // vC=-1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010110; // iC=  662 
vC = 14'b1111101010001011; // vC=-1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111010; // iC=  698 
vC = 14'b1111101001111101; // vC=-1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000101; // iC=  773 
vC = 14'b1111101000010011; // vC=-1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000110; // iC=  774 
vC = 14'b1111101000111111; // vC=-1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101111; // iC=  815 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111001; // iC=  761 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101111; // iC=  815 
vC = 14'b1111101001111011; // vC=-1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100101; // iC=  805 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000101; // iC=  901 
vC = 14'b1111101001111011; // vC=-1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010100; // iC=  852 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111111; // iC=  895 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100010; // iC=  994 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010000; // iC=  912 
vC = 14'b1111101000011000; // vC=-1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111000; // iC= 1016 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101000; // iC=  936 
vC = 14'b1111101010101110; // vC=-1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101110; // iC= 1006 
vC = 14'b1111101001111101; // vC=-1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100000; // iC= 1056 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101000; // iC= 1128 
vC = 14'b1111101010110000; // vC=-1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000010; // iC= 1026 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011001; // iC= 1113 
vC = 14'b1111101010111110; // vC=-1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001110; // iC= 1102 
vC = 14'b1111101001101110; // vC=-1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100000; // iC= 1120 
vC = 14'b1111101011010000; // vC=-1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010111; // iC= 1111 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101011; // iC= 1131 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010101; // iC= 1237 
vC = 14'b1111101001001001; // vC=-1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101000; // iC= 1256 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101000; // iC= 1192 
vC = 14'b1111101010110001; // vC=-1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110110; // iC= 1334 
vC = 14'b1111101001011001; // vC=-1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110010; // iC= 1266 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110110; // iC= 1334 
vC = 14'b1111101010011101; // vC=-1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011011; // iC= 1307 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001100; // iC= 1420 
vC = 14'b1111101010110101; // vC=-1355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010100; // iC= 1428 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010111; // iC= 1367 
vC = 14'b1111101100000010; // vC=-1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011111; // iC= 1439 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001001; // iC= 1417 
vC = 14'b1111101011011011; // vC=-1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110111; // iC= 1399 
vC = 14'b1111101010100100; // vC=-1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010001; // iC= 1425 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110001; // iC= 1457 
vC = 14'b1111101100010011; // vC=-1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100000; // iC= 1440 
vC = 14'b1111101011101110; // vC=-1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010001; // iC= 1489 
vC = 14'b1111101010101110; // vC=-1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001111; // iC= 1551 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001010; // iC= 1482 
vC = 14'b1111101011010101; // vC=-1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110010; // iC= 1522 
vC = 14'b1111101011110010; // vC=-1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000110; // iC= 1542 
vC = 14'b1111101100101000; // vC=-1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101010; // iC= 1578 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b1111101011010011; // vC=-1325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001110; // iC= 1614 
vC = 14'b1111101101010010; // vC=-1198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101110; // iC= 1582 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010011; // iC= 1747 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001010; // iC= 1738 
vC = 14'b1111101101111011; // vC=-1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011011; // iC= 1627 
vC = 14'b1111101100011011; // vC=-1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b1111101100011101; // vC=-1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101111; // iC= 1711 
vC = 14'b1111101100000100; // vC=-1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101000; // iC= 1704 
vC = 14'b1111101100111000; // vC=-1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101100; // iC= 1772 
vC = 14'b1111101101100101; // vC=-1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000110; // iC= 1798 
vC = 14'b1111101110101001; // vC=-1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101101; // iC= 1709 
vC = 14'b1111101110001111; // vC=-1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b1111101110100010; // vC=-1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b1111101101111001; // vC=-1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000000; // iC= 1792 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b1111101101110101; // vC=-1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b1111101101101010; // vC=-1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001101; // iC= 1869 
vC = 14'b1111101110011011; // vC=-1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101000; // iC= 1832 
vC = 14'b1111101111000101; // vC=-1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000100; // iC= 1796 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001000; // iC= 1864 
vC = 14'b1111101101110100; // vC=-1164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010100; // iC= 1876 
vC = 14'b1111101110111100; // vC=-1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111101110010001; // vC=-1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b1111101111011010; // vC=-1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b1111101110001101; // vC=-1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111101110111111; // vC=-1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b1111101110010110; // vC=-1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001010; // iC= 1866 
vC = 14'b1111101111000111; // vC=-1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111101110011110; // vC=-1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b1111101111101100; // vC=-1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111101111001001; // vC=-1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b1111101111001000; // vC=-1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000101; // iC= 1861 
vC = 14'b1111101111110111; // vC=-1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b1111101111010001; // vC=-1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111101111111000; // vC=-1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111110000010001; // vC=-1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b1111110001110010; // vC= -910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110010; // iC= 1906 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111110000110011; // vC= -973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111110001010100; // vC= -940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011001; // iC= 1881 
vC = 14'b1111110001000000; // vC= -960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111110000011011; // vC= -997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111110010001011; // vC= -885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101100; // iC= 1964 
vC = 14'b1111110010001110; // vC= -882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b1111110001110011; // vC= -909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111110010101011; // vC= -853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001010; // iC= 1866 
vC = 14'b1111110001010001; // vC= -943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001011; // iC= 1867 
vC = 14'b1111110011010001; // vC= -815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b1111110010100011; // vC= -861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110100; // iC= 1972 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111110010011100; // vC= -868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111110100000101; // vC= -763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111110011101110; // vC= -786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b1111110010001110; // vC= -882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b1111110010100101; // vC= -859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111110100011110; // vC= -738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b1111110010011001; // vC= -871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b1111110100000111; // vC= -761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111110100111011; // vC= -709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111110100000011; // vC= -765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111110100001011; // vC= -757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b1111110011000111; // vC= -825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100001; // iC= 2017 
vC = 14'b1111110101011011; // vC= -677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110100; // iC= 1972 
vC = 14'b1111110100000010; // vC= -766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111110100110010; // vC= -718 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b1111110100001011; // vC= -757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111110011110101; // vC= -779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111110100100011; // vC= -733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111110101100000; // vC= -672 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100010; // iC= 2018 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111111; // iC= 2047 
vC = 14'b1111110100101110; // vC= -722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111110100111011; // vC= -709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111110110010001; // vC= -623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000000; // iC= 2048 
vC = 14'b1111110101110101; // vC= -651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b1111110100111011; // vC= -709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110101011000; // vC= -680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111000; // iC= 2040 
vC = 14'b1111110101101000; // vC= -664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110101011000; // vC= -680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101100; // iC= 1964 
vC = 14'b1111110110100111; // vC= -601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111110110011010; // vC= -614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b1111110101111101; // vC= -643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011101; // iC= 2077 
vC = 14'b1111110111011011; // vC= -549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111110110001010; // vC= -630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101101; // iC= 2029 
vC = 14'b1111110110111001; // vC= -583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b1111110111000001; // vC= -575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111110110001100; // vC= -628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111000010111; // vC= -489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111110111001101; // vC= -563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111111000110110; // vC= -458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111110110111000; // vC= -584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b1111111000001100; // vC= -500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111000011011; // vC= -485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111110111111110; // vC= -514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111111001011010; // vC= -422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111111000101010; // vC= -470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011100; // iC= 1948 
vC = 14'b1111111001001101; // vC= -435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b1111111001011000; // vC= -424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111111000000100; // vC= -508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b1111111000101110; // vC= -466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111110; // iC= 1982 
vC = 14'b1111111000000001; // vC= -511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b1111111010001001; // vC= -375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111110111110010; // vC= -526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001100; // iC= 2060 
vC = 14'b1111110111111010; // vC= -518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b1111111010010011; // vC= -365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b1111111001000100; // vC= -444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001001; // iC= 2057 
vC = 14'b1111111001100110; // vC= -410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111010011011; // vC= -357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111111001000101; // vC= -443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b1111111001011110; // vC= -418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b1111111010010111; // vC= -361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000101000; // iC= 2088 
vC = 14'b1111111011000010; // vC= -318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b1111111001011110; // vC= -418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111111010101100; // vC= -340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000100; // iC= 2052 
vC = 14'b1111111011101101; // vC= -275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111111001101000; // vC= -408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111111011001010; // vC= -310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010011; // iC= 2067 
vC = 14'b1111111010110111; // vC= -329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b1111111010011101; // vC= -355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010001; // iC= 2065 
vC = 14'b1111111011001010; // vC= -310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111010010110; // vC= -362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111111010001111; // vC= -369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111010101000; // vC= -344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100011; // iC= 2083 
vC = 14'b1111111011101000; // vC= -280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111111011111110; // vC= -258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111111011101101; // vC= -275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111100100110; // vC= -218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b1111111100101010; // vC= -214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111111100011101; // vC= -227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100001; // iC= 2081 
vC = 14'b1111111101000011; // vC= -189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000101; // iC= 2053 
vC = 14'b1111111101001111; // vC= -177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111111011101101; // vC= -275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011101; // iC= 2077 
vC = 14'b1111111011010101; // vC= -299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111111101100000; // vC= -160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111111101011110; // vC= -162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111101; // iC= 2045 
vC = 14'b1111111101001010; // vC= -182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111011101111; // vC= -273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100001; // iC= 2017 
vC = 14'b1111111100101101; // vC= -211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111111100100000; // vC= -224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001100; // iC= 2060 
vC = 14'b1111111101101110; // vC= -146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b1111111101000011; // vC= -189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000011; // iC= 2051 
vC = 14'b1111111100110010; // vC= -206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111111110101110; // vC=  -82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010110; // iC= 2070 
vC = 14'b1111111110001100; // vC= -116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010101; // iC= 2069 
vC = 14'b1111111101111101; // vC= -131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011000; // iC= 2072 
vC = 14'b1111111100110111; // vC= -201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111111101010101; // vC= -171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111111101001010; // vC= -182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b1111111111001001; // vC=  -55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b1111111101101010; // vC= -150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b1111111111001000; // vC=  -56 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010001; // iC= 2065 
vC = 14'b1111111110000011; // vC= -125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b1111111110111000; // vC=  -72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111111110011110; // vC=  -98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111111101111101; // vC= -131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111111110111101; // vC=  -67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111111110010110; // vC= -106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b1111111111011110; // vC=  -34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b1111111111111010; // vC=   -6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101111; // iC= 2031 
vC = 14'b0000000000100100; // vC=   36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b0000000000000111; // vC=    7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111111111001010; // vC=  -54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b1111111111000100; // vC=  -60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b1111111111111100; // vC=   -4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111111111111110; // vC=   -2 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b0000000001101111; // vC=  111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b0000000000111001; // vC=   57 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b0000000000010001; // vC=   17 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b0000000000100010; // vC=   34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b0000000001011010; // vC=   90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b0000000010001110; // vC=  142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b0000000000011111; // vC=   31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101011; // iC= 2027 
vC = 14'b0000000000010010; // vC=   18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000000110100; // vC=   52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b0000000010011000; // vC=  152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100011; // iC= 2019 
vC = 14'b0000000001011010; // vC=   90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000000; // iC= 1984 
vC = 14'b0000000001111011; // vC=  123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b0000000001111001; // vC=  121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b0000000010001111; // vC=  143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b0000000011111001; // vC=  249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b0000000001101011; // vC=  107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b0000000011000101; // vC=  197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b0000000011011100; // vC=  220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b0000000011000100; // vC=  196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b0000000100000001; // vC=  257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b0000000010001111; // vC=  143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b0000000010100111; // vC=  167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b0000000100101011; // vC=  299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b0000000010101100; // vC=  172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b0000000011010111; // vC=  215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001010; // iC= 1994 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b0000000011001010; // vC=  202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b0000000011001011; // vC=  203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b0000000011011100; // vC=  220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b0000000100001111; // vC=  271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b0000000100010111; // vC=  279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b0000000100101101; // vC=  301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110000; // iC= 1840 
vC = 14'b0000000011101110; // vC=  238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b0000000101000000; // vC=  320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b0000000011110010; // vC=  242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b0000000110010111; // vC=  407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000010; // iC= 1858 
vC = 14'b0000000100000000; // vC=  256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b0000000101010000; // vC=  336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b0000000101001011; // vC=  331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b0000000110011000; // vC=  408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b0000000100100000; // vC=  288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b0000000110100001; // vC=  417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b0000000100110110; // vC=  310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b0000000110111011; // vC=  443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b0000000100111111; // vC=  319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b0000000101000000; // vC=  320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011100; // iC= 1884 
vC = 14'b0000000101011001; // vC=  345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000101; // iC= 1797 
vC = 14'b0000000101101101; // vC=  365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000000110001100; // vC=  396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001000; // iC= 1864 
vC = 14'b0000000110010111; // vC=  407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b0000000101010111; // vC=  343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110101; // iC= 1781 
vC = 14'b0000000110110100; // vC=  436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b0000000111011111; // vC=  479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110110; // iC= 1846 
vC = 14'b0000000101110100; // vC=  372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101010; // iC= 1898 
vC = 14'b0000000111011010; // vC=  474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b0000000111000100; // vC=  452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b0000000111000100; // vC=  452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111110; // iC= 1790 
vC = 14'b0000000111010100; // vC=  468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000000111101011; // vC=  491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b0000001000111001; // vC=  569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010000; // iC= 1808 
vC = 14'b0000000111111000; // vC=  504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b0000000111000011; // vC=  451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100010; // iC= 1826 
vC = 14'b0000001000001110; // vC=  526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000000111111001; // vC=  505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101011; // iC= 1835 
vC = 14'b0000001000111001; // vC=  569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b0000001001000000; // vC=  576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b0000000111100001; // vC=  481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001100; // iC= 1804 
vC = 14'b0000000111111000; // vC=  504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001011; // iC= 1739 
vC = 14'b0000001001010110; // vC=  598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b0000001000111110; // vC=  574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b0000001001010101; // vC=  597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000001000011100; // vC=  540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b0000001000100000; // vC=  544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b0000001000001101; // vC=  525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b0000001000101101; // vC=  557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b0000001001000100; // vC=  580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000011; // iC= 1795 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100001; // iC= 1697 
vC = 14'b0000001010111010; // vC=  698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101110; // iC= 1838 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b0000001010111100; // vC=  700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110101; // iC= 1717 
vC = 14'b0000001010011001; // vC=  665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100011; // iC= 1699 
vC = 14'b0000001001110100; // vC=  628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b0000001001110010; // vC=  626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b0000001010111101; // vC=  701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010101; // iC= 1685 
vC = 14'b0000001011000010; // vC=  706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010101; // iC= 1685 
vC = 14'b0000001011100101; // vC=  741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111110; // iC= 1790 
vC = 14'b0000001001110010; // vC=  626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111110; // iC= 1662 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111110; // iC= 1790 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b0000001100000001; // vC=  769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b0000001011010101; // vC=  725 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111110; // iC= 1726 
vC = 14'b0000001010101110; // vC=  686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b0000001010100101; // vC=  677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b0000001100010110; // vC=  790 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001000; // iC= 1672 
vC = 14'b0000001100011110; // vC=  798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b0000001010010110; // vC=  662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b0000001011000110; // vC=  710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011000; // iC= 1688 
vC = 14'b0000001010101101; // vC=  685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001010; // iC= 1738 
vC = 14'b0000001011100011; // vC=  739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110011; // iC= 1651 
vC = 14'b0000001011010110; // vC=  726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011101; // iC= 1693 
vC = 14'b0000001100111110; // vC=  830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100111; // iC= 1703 
vC = 14'b0000001011111001; // vC=  761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b0000001011100110; // vC=  742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b0000001011110110; // vC=  758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011011; // iC= 1627 
vC = 14'b0000001011010010; // vC=  722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111111; // iC= 1599 
vC = 14'b0000001100111110; // vC=  830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001100; // iC= 1612 
vC = 14'b0000001100100000; // vC=  800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b0000001101001011; // vC=  843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100101; // iC= 1637 
vC = 14'b0000001011101000; // vC=  744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b0000001100100001; // vC=  801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110101; // iC= 1589 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000000; // iC= 1664 
vC = 14'b0000001100101111; // vC=  815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111110; // iC= 1662 
vC = 14'b0000001100111010; // vC=  826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b0000001100111100; // vC=  828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000111; // iC= 1671 
vC = 14'b0000001100000110; // vC=  774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010000; // iC= 1616 
vC = 14'b0000001101000011; // vC=  835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011100; // iC= 1564 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011001; // iC= 1561 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b0000001101101011; // vC=  875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001101; // iC= 1677 
vC = 14'b0000001100011011; // vC=  795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011011; // iC= 1627 
vC = 14'b0000001101001100; // vC=  844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111011; // iC= 1659 
vC = 14'b0000001101110100; // vC=  884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b0000001100111110; // vC=  830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111001; // iC= 1657 
vC = 14'b0000001111001001; // vC=  969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b0000001100111111; // vC=  831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000110; // iC= 1606 
vC = 14'b0000001110100000; // vC=  928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001010; // iC= 1610 
vC = 14'b0000001101101111; // vC=  879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111111; // iC= 1535 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000001; // iC= 1665 
vC = 14'b0000001110000011; // vC=  899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001110011001; // vC=  921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101000; // iC= 1576 
vC = 14'b0000001110101011; // vC=  939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110100; // iC= 1652 
vC = 14'b0000001110111001; // vC=  953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011100; // iC= 1564 
vC = 14'b0000001110011111; // vC=  927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100101; // iC= 1637 
vC = 14'b0000001110110010; // vC=  946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011011; // iC= 1563 
vC = 14'b0000001111000100; // vC=  964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b0000001110000110; // vC=  902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010000; // iC= 1488 
vC = 14'b0000001110001011; // vC=  907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010010; // iC= 1554 
vC = 14'b0000001110110001; // vC=  945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111001; // iC= 1465 
vC = 14'b0000010000000100; // vC= 1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011110; // iC= 1566 
vC = 14'b0000001110100111; // vC=  935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110101; // iC= 1589 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111100; // iC= 1532 
vC = 14'b0000010000001000; // vC= 1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000000; // iC= 1472 
vC = 14'b0000001111001111; // vC=  975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b0000010000000110; // vC= 1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001110; // iC= 1550 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001101; // iC= 1485 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001000; // iC= 1480 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011110; // iC= 1502 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110101; // iC= 1525 
vC = 14'b0000001111011111; // vC=  991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110101; // iC= 1461 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110011; // iC= 1459 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b0000001111000011; // vC=  963 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000000; // iC= 1472 
vC = 14'b0000010000110101; // vC= 1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001011; // iC= 1483 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010110; // iC= 1430 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000011; // iC= 1539 
vC = 14'b0000010001000110; // vC= 1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011100; // iC= 1500 
vC = 14'b0000010001110010; // vC= 1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101011; // iC= 1387 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011110; // iC= 1502 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001111; // iC= 1487 
vC = 14'b0000010001000010; // vC= 1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110110; // iC= 1526 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011100; // iC= 1372 
vC = 14'b0000010010000100; // vC= 1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101100; // iC= 1452 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110110; // iC= 1398 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111010; // iC= 1402 
vC = 14'b0000010000000001; // vC= 1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001101; // iC= 1357 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110110; // iC= 1462 
vC = 14'b0000010000000111; // vC= 1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001001; // iC= 1481 
vC = 14'b0000010001101011; // vC= 1131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001110; // iC= 1422 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011010; // iC= 1370 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111000; // iC= 1400 
vC = 14'b0000010001010100; // vC= 1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101010; // iC= 1386 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001110; // iC= 1422 
vC = 14'b0000010001000111; // vC= 1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110001; // iC= 1393 
vC = 14'b0000010000100011; // vC= 1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101101; // iC= 1453 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111000; // iC= 1464 
vC = 14'b0000010010111000; // vC= 1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011101; // iC= 1309 
vC = 14'b0000010010100100; // vC= 1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010011; // iC= 1427 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101100; // iC= 1388 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011100; // iC= 1308 
vC = 14'b0000010010111000; // vC= 1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001101; // iC= 1421 
vC = 14'b0000010010010111; // vC= 1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011001; // iC= 1433 
vC = 14'b0000010001100101; // vC= 1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111101; // iC= 1341 
vC = 14'b0000010011001100; // vC= 1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010000; // iC= 1360 
vC = 14'b0000010011010000; // vC= 1232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100001; // iC= 1377 
vC = 14'b0000010011011001; // vC= 1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111100; // iC= 1340 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001001; // iC= 1289 
vC = 14'b0000010011110101; // vC= 1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101010; // iC= 1258 
vC = 14'b0000010001011111; // vC= 1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100011; // iC= 1315 
vC = 14'b0000010100000101; // vC= 1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100110; // iC= 1382 
vC = 14'b0000010001101110; // vC= 1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000111; // iC= 1351 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110101; // iC= 1333 
vC = 14'b0000010100000111; // vC= 1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001001; // iC= 1225 
vC = 14'b0000010011000010; // vC= 1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010000; // iC= 1360 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001111; // iC= 1231 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111100; // iC= 1276 
vC = 14'b0000010011110011; // vC= 1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000111; // iC= 1287 
vC = 14'b0000010100100011; // vC= 1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001111; // iC= 1295 
vC = 14'b0000010100000001; // vC= 1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110000; // iC= 1328 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011010; // iC= 1306 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000011; // iC= 1219 
vC = 14'b0000010010110111; // vC= 1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111110; // iC= 1214 
vC = 14'b0000010100100000; // vC= 1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000010; // iC= 1282 
vC = 14'b0000010100010101; // vC= 1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110101; // iC= 1269 
vC = 14'b0000010011111010; // vC= 1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001111; // iC= 1231 
vC = 14'b0000010011010101; // vC= 1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101111; // iC= 1263 
vC = 14'b0000010011110100; // vC= 1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101000; // iC= 1192 
vC = 14'b0000010011101111; // vC= 1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011100; // iC= 1308 
vC = 14'b0000010101001111; // vC= 1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000000; // iC= 1280 
vC = 14'b0000010100011000; // vC= 1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110110; // iC= 1270 
vC = 14'b0000010011011000; // vC= 1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101010; // iC= 1194 
vC = 14'b0000010011010001; // vC= 1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000110; // iC= 1158 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110001; // iC= 1265 
vC = 14'b0000010011110110; // vC= 1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001110; // iC= 1230 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001111; // iC= 1231 
vC = 14'b0000010011110111; // vC= 1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100010; // iC= 1250 
vC = 14'b0000010100001010; // vC= 1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000010101101001; // vC= 1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111010; // iC= 1210 
vC = 14'b0000010011101001; // vC= 1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000010; // iC= 1218 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000011; // iC= 1219 
vC = 14'b0000010101100110; // vC= 1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010011; // iC= 1171 
vC = 14'b0000010011100011; // vC= 1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101101; // iC= 1133 
vC = 14'b0000010101111001; // vC= 1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011010; // iC= 1114 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100111; // iC= 1127 
vC = 14'b0000010101111000; // vC= 1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011111; // iC= 1183 
vC = 14'b0000010011111100; // vC= 1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010101; // iC= 1173 
vC = 14'b0000010101111101; // vC= 1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111001; // iC= 1145 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000000; // iC= 1152 
vC = 14'b0000010100000010; // vC= 1282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001011; // iC= 1099 
vC = 14'b0000010100000110; // vC= 1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110000; // iC= 1072 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000110; // iC= 1158 
vC = 14'b0000010101110101; // vC= 1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110010; // iC= 1138 
vC = 14'b0000010100100001; // vC= 1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101000; // iC= 1128 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011011; // iC= 1051 
vC = 14'b0000010101100111; // vC= 1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010100; // iC= 1108 
vC = 14'b0000010101101111; // vC= 1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100010; // iC= 1122 
vC = 14'b0000010100100101; // vC= 1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001101; // iC= 1101 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010011; // iC= 1043 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110101; // iC= 1077 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010011; // iC= 1107 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000111; // iC= 1095 
vC = 14'b0000010100110110; // vC= 1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010011; // iC= 1107 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010000; // iC= 1040 
vC = 14'b0000010101101110; // vC= 1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001000; // iC= 1096 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111111; // iC=  959 
vC = 14'b0000010111001000; // vC= 1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100001; // iC=  993 
vC = 14'b0000010101111000; // vC= 1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101101; // iC= 1005 
vC = 14'b0000010101001001; // vC= 1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110000; // iC=  944 
vC = 14'b0000010111010100; // vC= 1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011101; // iC= 1053 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100010; // iC=  994 
vC = 14'b0000010110010110; // vC= 1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100011; // iC=  995 
vC = 14'b0000010101100010; // vC= 1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100101; // iC= 1061 
vC = 14'b0000010110011001; // vC= 1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000100; // iC= 1028 
vC = 14'b0000010101010101; // vC= 1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100010; // iC= 1058 
vC = 14'b0000010101100101; // vC= 1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001110; // iC= 1038 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011111; // iC= 1055 
vC = 14'b0000010110011111; // vC= 1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110101; // iC= 1013 
vC = 14'b0000010110011111; // vC= 1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001111; // iC=  975 
vC = 14'b0000010111101001; // vC= 1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111101; // iC=  957 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110101; // iC=  949 
vC = 14'b0000010111111000; // vC= 1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000100; // iC= 1028 
vC = 14'b0000010110010101; // vC= 1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110010; // iC=  882 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b0000010111000010; // vC= 1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001000; // iC=  968 
vC = 14'b0000010101101010; // vC= 1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111011; // iC=  955 
vC = 14'b0000010110011011; // vC= 1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111000; // iC=  888 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100000; // iC=  992 
vC = 14'b0000010110001110; // vC= 1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001000; // iC=  968 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111001; // iC=  825 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110000; // iC=  880 
vC = 14'b0000010110111101; // vC= 1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110100; // iC=  884 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111110; // iC=  894 
vC = 14'b0000010111000001; // vC= 1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111100; // iC=  956 
vC = 14'b0000010110100010; // vC= 1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000111; // iC=  839 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010010; // iC=  914 
vC = 14'b0000010111110001; // vC= 1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100000; // iC=  928 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111100; // iC=  828 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010111; // iC=  791 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100000; // iC=  928 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000111; // iC=  903 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010010; // iC=  850 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001101; // iC=  909 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001000; // iC=  904 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010011; // iC=  787 
vC = 14'b0000010111001001; // vC= 1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100000; // iC=  736 
vC = 14'b0000010111010101; // vC= 1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010010; // iC=  850 
vC = 14'b0000010111010100; // vC= 1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100010; // iC=  866 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011011; // iC=  731 
vC = 14'b0000010110100011; // vC= 1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101110; // iC=  814 
vC = 14'b0000010111000100; // vC= 1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101111; // iC=  751 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000011; // iC=  771 
vC = 14'b0000011000101011; // vC= 1579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001010; // iC=  842 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101101; // iC=  749 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100010; // iC=  738 
vC = 14'b0000010111100100; // vC= 1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110011; // iC=  691 
vC = 14'b0000010111010100; // vC= 1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111100; // iC=  700 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110011; // iC=  691 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110011; // iC=  819 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010010; // iC=  786 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001011; // iC=  715 
vC = 14'b0000010111000001; // vC= 1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100001; // iC=  801 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110001; // iC=  753 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010101; // iC=  725 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100100; // iC=  676 
vC = 14'b0000010111110111; // vC= 1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101000; // iC=  744 
vC = 14'b0000011000001001; // vC= 1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110011; // iC=  755 
vC = 14'b0000011000110100; // vC= 1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000001; // iC=  641 
vC = 14'b0000011000101111; // vC= 1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100001; // iC=  673 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110100; // iC=  692 
vC = 14'b0000011000110010; // vC= 1586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110011; // iC=  691 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101000; // iC=  616 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000011; // iC=  643 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111011; // iC=  635 
vC = 14'b0000011001001110; // vC= 1614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001100; // iC=  652 
vC = 14'b0000011001000000; // vC= 1600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000110; // iC=  646 
vC = 14'b0000011000101011; // vC= 1579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011100; // iC=  668 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000100; // iC=  644 
vC = 14'b0000011001110010; // vC= 1650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101110; // iC=  558 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101001; // iC=  617 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101101; // iC=  685 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001101; // iC=  525 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101101; // iC=  621 
vC = 14'b0000011010000101; // vC= 1669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110011; // iC=  563 
vC = 14'b0000010111110100; // vC= 1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010110; // iC=  598 
vC = 14'b0000011001101100; // vC= 1644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111101; // iC=  573 
vC = 14'b0000010111111111; // vC= 1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000110; // iC=  582 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000001; // iC=  577 
vC = 14'b0000010111101100; // vC= 1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010100; // iC=  596 
vC = 14'b0000011001111100; // vC= 1660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011000; // iC=  536 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110000; // iC=  624 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000010; // iC=  514 
vC = 14'b0000011010000100; // vC= 1668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011111; // iC=  479 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100001; // iC=  609 
vC = 14'b0000011001100101; // vC= 1637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000100; // iC=  580 
vC = 14'b0000011001110110; // vC= 1654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011011; // iC=  539 
vC = 14'b0000011001000010; // vC= 1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011110; // iC=  542 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000011; // iC=  451 
vC = 14'b0000011001101110; // vC= 1646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101011; // iC=  427 
vC = 14'b0000011010000110; // vC= 1670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011111; // iC=  543 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110101; // iC=  501 
vC = 14'b0000011000110010; // vC= 1586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100100; // iC=  420 
vC = 14'b0000011010010011; // vC= 1683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110110; // iC=  438 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000100; // iC=  516 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111001; // iC=  441 
vC = 14'b0000011001010001; // vC= 1617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111101; // iC=  445 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011111; // iC=  479 
vC = 14'b0000011010010010; // vC= 1682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100011; // iC=  419 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100011; // iC=  419 
vC = 14'b0000011000101000; // vC= 1576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010011; // iC=  403 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001110; // iC=  398 
vC = 14'b0000011001110101; // vC= 1653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110111; // iC=  311 
vC = 14'b0000011010000110; // vC= 1670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010010; // iC=  402 
vC = 14'b0000011010011011; // vC= 1691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000010; // iC=  322 
vC = 14'b0000011010100100; // vC= 1700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100011; // iC=  355 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110101; // iC=  309 
vC = 14'b0000011010100010; // vC= 1698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010100; // iC=  276 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100101; // iC=  293 
vC = 14'b0000011000101011; // vC= 1579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111111; // iC=  319 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101110; // iC=  174 
vC = 14'b0000011001100111; // vC= 1639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001011; // iC=  267 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001000; // iC=  136 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000110; // iC=  134 
vC = 14'b0000011010010000; // vC= 1680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101111; // iC=  239 
vC = 14'b0000011010100010; // vC= 1698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100110; // iC=  166 
vC = 14'b0000011001010010; // vC= 1618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010111; // iC=   87 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001000; // iC=   72 
vC = 14'b0000011000101000; // vC= 1576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001011; // iC=  203 
vC = 14'b0000011001110011; // vC= 1651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010011; // iC=  147 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101111; // iC=  111 
vC = 14'b0000011001101000; // vC= 1640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001001; // iC=   73 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001100; // iC=   12 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010110; // iC=   22 
vC = 14'b0000011000110001; // vC= 1585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111000; // iC=   56 
vC = 14'b0000011010000000; // vC= 1664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001110; // iC=   78 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000111; // iC=    7 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100011; // iC=   35 
vC = 14'b0000011000010111; // vC= 1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000111; // iC=  -57 
vC = 14'b0000011000001001; // vC= 1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011010; // iC=  -38 
vC = 14'b0000011010010000; // vC= 1680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000100; // iC= -124 
vC = 14'b0000011001010010; // vC= 1618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100001; // iC= -159 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101010; // iC= -150 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001101; // iC= -115 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110011; // iC= -141 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010100; // iC= -172 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010001; // iC= -239 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110010; // iC= -206 
vC = 14'b0000011000111101; // vC= 1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101000; // iC= -280 
vC = 14'b0000011010001101; // vC= 1677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110110; // iC= -266 
vC = 14'b0000011001010111; // vC= 1623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101000; // iC= -280 
vC = 14'b0000011010010110; // vC= 1686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100011; // iC= -349 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011101; // iC= -291 
vC = 14'b0000011000101101; // vC= 1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001001; // iC= -311 
vC = 14'b0000011010010000; // vC= 1680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101011; // iC= -341 
vC = 14'b0000011000111101; // vC= 1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001010; // iC= -374 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001011; // iC= -373 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010000; // iC= -368 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001010; // iC= -502 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001011; // iC= -501 
vC = 14'b0000011000001101; // vC= 1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101011; // iC= -469 
vC = 14'b0000011000101000; // vC= 1576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000110; // iC= -442 
vC = 14'b0000010111100011; // vC= 1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000001; // iC= -575 
vC = 14'b0000011001101000; // vC= 1640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010011; // iC= -493 
vC = 14'b0000010111101011; // vC= 1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100110; // iC= -602 
vC = 14'b0000011001011100; // vC= 1628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110010; // iC= -526 
vC = 14'b0000011001011110; // vC= 1630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101101; // iC= -659 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b0000011001011101; // vC= 1629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111010; // iC= -710 
vC = 14'b0000011000110101; // vC= 1589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110000; // iC= -656 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001000; // iC= -696 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b0000011000101000; // vC= 1576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110101; // iC= -779 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111111; // iC= -769 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111110; // iC= -770 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001011; // iC= -885 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011101; // iC= -867 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011110; // iC= -802 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001001; // iC= -823 
vC = 14'b0000011000001101; // vC= 1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001001; // iC= -951 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101110; // iC= -914 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100011; // iC= -925 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001110; // iC= -882 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111111; // iC=-1025 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011110; // iC=-1058 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111101; // iC= -963 
vC = 14'b0000010111011110; // vC= 1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000001; // iC= -959 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110011; // iC= -973 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010010; // iC=-1134 
vC = 14'b0000010111010110; // vC= 1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011010; // iC=-1126 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100000; // iC=-1120 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011111; // iC=-1121 
vC = 14'b0000010111101010; // vC= 1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010010; // iC=-1198 
vC = 14'b0000010110011011; // vC= 1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101001; // iC=-1111 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101000; // iC=-1176 
vC = 14'b0000011000000001; // vC= 1537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111010; // iC=-1222 
vC = 14'b0000010110011011; // vC= 1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b0000010101100110; // vC= 1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100011; // iC=-1181 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000010; // iC=-1278 
vC = 14'b0000010111111000; // vC= 1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011100; // iC=-1188 
vC = 14'b0000010110001010; // vC= 1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011000; // iC=-1256 
vC = 14'b0000010110111101; // vC= 1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111111; // iC=-1345 
vC = 14'b0000010111011001; // vC= 1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000111; // iC=-1209 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000000; // iC=-1344 
vC = 14'b0000010110001101; // vC= 1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110111; // iC=-1289 
vC = 14'b0000010101001110; // vC= 1358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010111; // iC=-1385 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001000; // iC=-1272 
vC = 14'b0000010101001001; // vC= 1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000010; // iC=-1278 
vC = 14'b0000010101111100; // vC= 1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110101; // iC=-1419 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110100; // iC=-1292 
vC = 14'b0000010100111111; // vC= 1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011010; // iC=-1318 
vC = 14'b0000010100100000; // vC= 1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111101; // iC=-1411 
vC = 14'b0000010110110100; // vC= 1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b0000010101100110; // vC= 1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100110; // iC=-1434 
vC = 14'b0000010110011111; // vC= 1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010010; // iC=-1390 
vC = 14'b0000010011111101; // vC= 1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110011; // iC=-1421 
vC = 14'b0000010101110111; // vC= 1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b0000010101010111; // vC= 1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b0000010101111000; // vC= 1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b0000010100100010; // vC= 1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010010; // iC=-1518 
vC = 14'b0000010100111101; // vC= 1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011101; // iC=-1571 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b0000010101100111; // vC= 1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101101; // iC=-1555 
vC = 14'b0000010011110110; // vC= 1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111101; // iC=-1603 
vC = 14'b0000010011111101; // vC= 1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b0000010101010110; // vC= 1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110001; // iC=-1487 
vC = 14'b0000010010111111; // vC= 1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b0000010100010011; // vC= 1299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000010011111100; // vC= 1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b0000010100010100; // vC= 1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b0000010100100010; // vC= 1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011010; // iC=-1574 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b0000010010111111; // vC= 1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111101; // iC=-1539 
vC = 14'b0000010010110111; // vC= 1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b0000010010011010; // vC= 1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000010011101010; // vC= 1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b0000010010101001; // vC= 1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b0000010001111001; // vC= 1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000010010011110; // vC= 1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011001; // iC=-1639 
vC = 14'b0000010010101011; // vC= 1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010100; // iC=-1644 
vC = 14'b0000010010101111; // vC= 1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100101; // iC=-1627 
vC = 14'b0000010001100011; // vC= 1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011111; // iC=-1633 
vC = 14'b0000010000100000; // vC= 1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000010010011000; // vC= 1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b0000010010100001; // vC= 1185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b0000010010000100; // vC= 1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b0000010001110010; // vC= 1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000010001101001; // vC= 1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110110; // iC=-1674 
vC = 14'b0000001111011111; // vC=  991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000010000010100; // vC= 1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b0000010000111010; // vC= 1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b0000001111011101; // vC=  989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000010000010001; // vC= 1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b0000010000001100; // vC= 1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000010; // iC=-1662 
vC = 14'b0000010000111011; // vC= 1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000001111110111; // vC= 1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111100; // iC=-1668 
vC = 14'b0000010000010001; // vC= 1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b0000001110010110; // vC=  918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000010000001001; // vC= 1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000010000000010; // vC= 1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000010000000001; // vC= 1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b0000001110101100; // vC=  940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b0000001110000101; // vC=  901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b0000001110110110; // vC=  950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000001110011011; // vC=  923 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000001110011100; // vC=  924 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b0000001101010111; // vC=  855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000001101000111; // vC=  839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000001110001001; // vC=  905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101010; // iC=-1686 
vC = 14'b0000001101011100; // vC=  860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111100; // iC=-1668 
vC = 14'b0000001101001100; // vC=  844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000001110101001; // vC=  937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000001110000001; // vC=  897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b0000001110001101; // vC=  909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001110011010; // vC=  922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001110011111; // vC=  927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000001100001110; // vC=  782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b0000001110010011; // vC=  915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000001101000000; // vC=  832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000001110000000; // vC=  896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000001100010000; // vC=  784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000001011110000; // vC=  752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000001011100110; // vC=  742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000001011110000; // vC=  752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b0000001011000010; // vC=  706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001100011111; // vC=  799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010000; // iC=-1840 
vC = 14'b0000001100000110; // vC=  774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000001011100111; // vC=  743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b0000001100110110; // vC=  822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000001010011001; // vC=  665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000001010111001; // vC=  697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000001010000000; // vC=  640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000001010011011; // vC=  667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000001011010111; // vC=  727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000001011010110; // vC=  726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000001011100000; // vC=  736 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000001001100110; // vC=  614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b0000001011000101; // vC=  709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001010110111; // vC=  695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000001010011100; // vC=  668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000001010110011; // vC=  691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110100; // iC=-1868 
vC = 14'b0000001001110010; // vC=  626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000001001010110; // vC=  598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001010010011; // vC=  659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000001001110010; // vC=  626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000001010101110; // vC=  686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000001001000101; // vC=  581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110000; // iC=-1872 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001001010000; // vC=  592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000001001001101; // vC=  589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000001000011000; // vC=  536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000001001000001; // vC=  577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001111; // iC=-1841 
vC = 14'b0000001000001000; // vC=  520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b0000000111101000; // vC=  488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b0000001000001000; // vC=  520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000001000001100; // vC=  524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110001; // iC=-1871 
vC = 14'b0000001001011100; // vC=  604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101010; // iC=-1878 
vC = 14'b0000000111110011; // vC=  499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000001000001011; // vC=  523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000001001001110; // vC=  590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111000; // iC=-1864 
vC = 14'b0000000111111010; // vC=  506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000001000001100; // vC=  524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000001000011111; // vC=  543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000001000001000; // vC=  520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000001000011001; // vC=  537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000000111101010; // vC=  490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b0000000111010111; // vC=  471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000000111101100; // vC=  492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000000110111111; // vC=  447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000001000000000; // vC=  512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101000; // iC=-1880 
vC = 14'b0000000110001001; // vC=  393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b0000000111010101; // vC=  469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000000101000111; // vC=  327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000101101110; // vC=  366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110010; // iC=-1870 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000000110110011; // vC=  435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000000110000101; // vC=  389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101001; // iC=-1815 
vC = 14'b0000000101111101; // vC=  381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000000100111001; // vC=  313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b0000000110001100; // vC=  396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000000110000100; // vC=  388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000000100010000; // vC=  272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000000110001000; // vC=  392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000000110001001; // vC=  393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110011; // iC=-1741 
vC = 14'b0000000101101111; // vC=  367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b0000000101111000; // vC=  376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000000101000100; // vC=  324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101110; // iC=-1874 
vC = 14'b0000000011110110; // vC=  246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000000011110000; // vC=  240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101101; // iC=-1875 
vC = 14'b0000000100011100; // vC=  284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111010; // iC=-1862 
vC = 14'b0000000011100010; // vC=  226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000000101010101; // vC=  341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000000011000000; // vC=  192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000000011100111; // vC=  231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000000100100111; // vC=  295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000000100101111; // vC=  303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b0000000100011001; // vC=  281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000000100000000; // vC=  256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000111; // iC=-1849 
vC = 14'b0000000010100100; // vC=  164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110000; // iC=-1872 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000000011011001; // vC=  217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000000100010101; // vC=  277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000000100010011; // vC=  275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111101; // iC=-1859 
vC = 14'b0000000011000011; // vC=  195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000000011111011; // vC=  251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111111; // iC=-1857 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111011; // iC=-1797 
vC = 14'b0000000001010101; // vC=   85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b0000000010111110; // vC=  190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110110; // iC=-1866 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000000010110101; // vC=  181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111101; // iC=-1859 
vC = 14'b0000000010100111; // vC=  167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111100; // iC=-1860 
vC = 14'b0000000010110001; // vC=  177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000000010100101; // vC=  165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000000000100110; // vC=   38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b0000000010111000; // vC=  184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000000000010101; // vC=   21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b1111111111110110; // vC=  -10 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000000000100101; // vC=   37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b1111111111111111; // vC=   -1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000000001101000; // vC=  104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b1111111110111100; // vC=  -68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b1111111111011100; // vC=  -36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000000001001111; // vC=   79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b1111111111111100; // vC=   -4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b1111111111010111; // vC=  -41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b1111111111110010; // vC=  -14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000000100100; // vC=   36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b1111111111100101; // vC=  -27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b1111111110010111; // vC= -105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b1111111110010111; // vC= -105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b1111111111110011; // vC=  -13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101010; // iC=-1686 
vC = 14'b1111111111000010; // vC=  -62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b1111111111111010; // vC=   -6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b1111111101101010; // vC= -150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b1111111111000101; // vC=  -59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b1111111111000100; // vC=  -60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b1111111110001011; // vC= -117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b1111111101101001; // vC= -151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b1111111101110110; // vC= -138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b1111111110010100; // vC= -108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b1111111110100111; // vC=  -89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b1111111101111010; // vC= -134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b1111111101011010; // vC= -166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b1111111101110001; // vC= -143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b1111111101011000; // vC= -168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b1111111101110000; // vC= -144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b1111111110011110; // vC=  -98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101010; // iC=-1686 
vC = 14'b1111111100001010; // vC= -246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b1111111101100001; // vC= -159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b1111111101001001; // vC= -183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b1111111100010011; // vC= -237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b1111111011101000; // vC= -280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b1111111100001010; // vC= -246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b1111111100001101; // vC= -243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b1111111101110000; // vC= -144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b1111111101011101; // vC= -163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b1111111100110001; // vC= -207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b1111111100100000; // vC= -224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000001; // iC=-1663 
vC = 14'b1111111100100010; // vC= -222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b1111111100110110; // vC= -202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b1111111011000000; // vC= -320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100101; // iC=-1691 
vC = 14'b1111111011101010; // vC= -278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b1111111010010110; // vC= -362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b1111111010100100; // vC= -348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011000; // iC=-1704 
vC = 14'b1111111100001010; // vC= -246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000100; // iC=-1724 
vC = 14'b1111111011010010; // vC= -302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b1111111010110010; // vC= -334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b1111111010000111; // vC= -377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b1111111011110011; // vC= -269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b1111111010100101; // vC= -347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b1111111010010001; // vC= -367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b1111111010110110; // vC= -330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b1111111010100101; // vC= -347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b1111111011101111; // vC= -273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110110; // iC=-1610 
vC = 14'b1111111010010101; // vC= -363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b1111111001001110; // vC= -434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b1111111010010101; // vC= -363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b1111111010001001; // vC= -375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b1111111011001100; // vC= -308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b1111111001011011; // vC= -421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111001; // iC=-1607 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100100; // iC=-1628 
vC = 14'b1111111010101100; // vC= -340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b1111111000011000; // vC= -488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101010; // iC=-1558 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b1111111001110110; // vC= -394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b1111111010000111; // vC= -377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b1111111001010111; // vC= -425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b1111111001000010; // vC= -446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b1111111000110000; // vC= -464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b1111111000000100; // vC= -508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b1111111000011000; // vC= -488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b1111110111111110; // vC= -514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101000; // iC=-1688 
vC = 14'b1111110111011110; // vC= -546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b1111110111101010; // vC= -534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010100; // iC=-1644 
vC = 14'b1111111001001010; // vC= -438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b1111110111011100; // vC= -548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000000; // iC=-1536 
vC = 14'b1111110111011011; // vC= -549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110111; // iC=-1609 
vC = 14'b1111111000000001; // vC= -511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010011; // iC=-1517 
vC = 14'b1111110111011000; // vC= -552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b1111110111111000; // vC= -520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001111; // iC=-1521 
vC = 14'b1111111000100100; // vC= -476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101011; // iC=-1557 
vC = 14'b1111110110110111; // vC= -585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b1111111000100001; // vC= -479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b1111110111011100; // vC= -548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b1111110110110110; // vC= -586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b1111110110010011; // vC= -621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b1111110111100001; // vC= -543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101110; // iC=-1618 
vC = 14'b1111110111011010; // vC= -550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b1111110110010000; // vC= -624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b1111110101111001; // vC= -647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b1111110110010101; // vC= -619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101111; // iC=-1553 
vC = 14'b1111110111111101; // vC= -515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001100; // iC=-1588 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000011; // iC=-1533 
vC = 14'b1111110111000110; // vC= -570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001010; // iC=-1526 
vC = 14'b1111110111001010; // vC= -566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b1111110111010101; // vC= -555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b1111110110000010; // vC= -638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b1111110110111010; // vC= -582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101101; // iC=-1555 
vC = 14'b1111110110010111; // vC= -617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110000; // iC=-1488 
vC = 14'b1111110110110101; // vC= -587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101010; // iC=-1558 
vC = 14'b1111110101110110; // vC= -650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b1111110100110110; // vC= -714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b1111110101011000; // vC= -680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110111; // iC=-1481 
vC = 14'b1111110100101001; // vC= -727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111101; // iC=-1539 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b1111110110011010; // vC= -614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b1111110101000100; // vC= -700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100010; // iC=-1502 
vC = 14'b1111110100101111; // vC= -721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b1111110101111010; // vC= -646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000011; // iC=-1533 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100100; // iC=-1500 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110101; // iC=-1483 
vC = 14'b1111110110000010; // vC= -638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000110; // iC=-1402 
vC = 14'b1111110100100010; // vC= -734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b1111110101010100; // vC= -684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111110; // iC=-1538 
vC = 14'b1111110011100110; // vC= -794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b1111110101110100; // vC= -652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b1111110011110110; // vC= -778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110000; // iC=-1488 
vC = 14'b1111110011101100; // vC= -788 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111011; // iC=-1541 
vC = 14'b1111110100010000; // vC= -752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111101; // iC=-1411 
vC = 14'b1111110100100011; // vC= -733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110100; // iC=-1484 
vC = 14'b1111110100010000; // vC= -752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b1111110100000000; // vC= -768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b1111110011011001; // vC= -807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010101; // iC=-1451 
vC = 14'b1111110011110000; // vC= -784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111101; // iC=-1411 
vC = 14'b1111110011110100; // vC= -780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101011; // iC=-1493 
vC = 14'b1111110100011111; // vC= -737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b1111110100001111; // vC= -753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010010; // iC=-1454 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000100; // iC=-1404 
vC = 14'b1111110010101011; // vC= -853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b1111110010010101; // vC= -875 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110000; // iC=-1488 
vC = 14'b1111110011010111; // vC= -809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000101; // iC=-1339 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b1111110011010010; // vC= -814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001100; // iC=-1332 
vC = 14'b1111110010100111; // vC= -857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b1111110010100111; // vC= -857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b1111110010001110; // vC= -882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b1111110010110001; // vC= -847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111000; // iC=-1352 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100011; // iC=-1309 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111010; // iC=-1350 
vC = 14'b1111110001111101; // vC= -899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101101; // iC=-1363 
vC = 14'b1111110001100101; // vC= -923 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110001; // iC=-1295 
vC = 14'b1111110010001111; // vC= -881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110101; // iC=-1291 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010101; // iC=-1323 
vC = 14'b1111110010100000; // vC= -864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101010; // iC=-1366 
vC = 14'b1111110010001011; // vC= -885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b1111110011000011; // vC= -829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000111; // iC=-1337 
vC = 14'b1111110011011001; // vC= -807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001000; // iC=-1272 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011101; // iC=-1315 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010100; // iC=-1324 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001011; // iC=-1333 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000101; // iC=-1275 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111011; // iC=-1285 
vC = 14'b1111110010100110; // vC= -858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101001; // iC=-1367 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011100; // iC=-1316 
vC = 14'b1111110001110110; // vC= -906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001110; // iC=-1394 
vC = 14'b1111110000010011; // vC=-1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110000; // iC=-1232 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101001; // iC=-1239 
vC = 14'b1111110000011010; // vC= -998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100011; // iC=-1309 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b1111110010000100; // vC= -892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101001; // iC=-1303 
vC = 14'b1111110001000111; // vC= -953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111001; // iC=-1223 
vC = 14'b1111110000001000; // vC=-1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000111; // iC=-1273 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110011; // iC=-1357 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111111; // iC=-1345 
vC = 14'b1111101111110011; // vC=-1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111110; // iC=-1218 
vC = 14'b1111110000110010; // vC= -974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010000; // iC=-1200 
vC = 14'b1111110000101001; // vC= -983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011001; // iC=-1319 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011110; // iC=-1314 
vC = 14'b1111110000110111; // vC= -969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b1111110001000110; // vC= -954 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011100; // iC=-1188 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011011; // iC=-1189 
vC = 14'b1111110000101101; // vC= -979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000100; // iC=-1276 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101110; // iC=-1234 
vC = 14'b1111101111101100; // vC=-1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100010; // iC=-1310 
vC = 14'b1111101111001011; // vC=-1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111101; // iC=-1283 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b1111110000110111; // vC= -969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001011; // iC=-1141 
vC = 14'b1111101110101000; // vC=-1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100011; // iC=-1181 
vC = 14'b1111101111110011; // vC=-1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100001; // iC=-1247 
vC = 14'b1111101110101011; // vC=-1109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100011; // iC=-1181 
vC = 14'b1111101111110110; // vC=-1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010100; // iC=-1196 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111110; // iC=-1154 
vC = 14'b1111110000011000; // vC=-1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110101; // iC=-1163 
vC = 14'b1111101111000000; // vC=-1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010001; // iC=-1199 
vC = 14'b1111101111010011; // vC=-1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b1111101111100110; // vC=-1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100000; // iC=-1184 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111001; // iC=-1095 
vC = 14'b1111101110111101; // vC=-1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010100; // iC=-1196 
vC = 14'b1111101110110000; // vC=-1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000000; // iC=-1152 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000001; // iC=-1151 
vC = 14'b1111101110001100; // vC=-1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000111; // iC=-1209 
vC = 14'b1111101110011110; // vC=-1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010111; // iC=-1065 
vC = 14'b1111101110000000; // vC=-1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100000; // iC=-1120 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000101; // iC=-1147 
vC = 14'b1111101111001000; // vC=-1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011101; // iC=-1123 
vC = 14'b1111101101011000; // vC=-1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011000; // iC=-1064 
vC = 14'b1111101101110001; // vC=-1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000001; // iC=-1087 
vC = 14'b1111101101010101; // vC=-1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001000; // iC=-1144 
vC = 14'b1111101110110101; // vC=-1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110101; // iC=-1035 
vC = 14'b1111101110110111; // vC=-1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001000; // iC=-1080 
vC = 14'b1111101101001010; // vC=-1206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000000; // iC=-1152 
vC = 14'b1111101110111010; // vC=-1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001000; // iC=-1080 
vC = 14'b1111101110110101; // vC=-1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101100; // iC=-1172 
vC = 14'b1111101101011110; // vC=-1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110000; // iC=-1040 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011101; // iC=-1059 
vC = 14'b1111101101011101; // vC=-1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011001; // iC=-1127 
vC = 14'b1111101110110100; // vC=-1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010000; // iC=-1008 
vC = 14'b1111101100110101; // vC=-1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001011; // iC=-1141 
vC = 14'b1111101100110001; // vC=-1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100000; // iC=-1056 
vC = 14'b1111101110000000; // vC=-1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111001; // iC=-1031 
vC = 14'b1111101110010111; // vC=-1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011011; // iC=-1061 
vC = 14'b1111101100111110; // vC=-1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011110; // iC=-1122 
vC = 14'b1111101100110100; // vC=-1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100001; // iC= -991 
vC = 14'b1111101110100111; // vC=-1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011101; // iC=-1059 
vC = 14'b1111101101000101; // vC=-1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000000; // iC= -960 
vC = 14'b1111101110101000; // vC=-1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111011; // iC=-1029 
vC = 14'b1111101110010000; // vC=-1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001001; // iC= -951 
vC = 14'b1111101101110110; // vC=-1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011010; // iC=-1062 
vC = 14'b1111101101110100; // vC=-1164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011110; // iC=-1058 
vC = 14'b1111101100000101; // vC=-1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001000; // iC=-1080 
vC = 14'b1111101100010010; // vC=-1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010111; // iC= -937 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001010; // iC=-1014 
vC = 14'b1111101100111010; // vC=-1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000000; // iC= -960 
vC = 14'b1111101101101000; // vC=-1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111100; // iC=-1028 
vC = 14'b1111101101101000; // vC=-1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100101; // iC=-1051 
vC = 14'b1111101100001101; // vC=-1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110000; // iC=-1040 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110101; // iC= -971 
vC = 14'b1111101101111001; // vC=-1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111111; // iC=-1025 
vC = 14'b1111101100011110; // vC=-1250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001110; // iC= -882 
vC = 14'b1111101011101110; // vC=-1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111100; // iC= -964 
vC = 14'b1111101101010011; // vC=-1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110001; // iC= -975 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110001; // iC= -975 
vC = 14'b1111101011011110; // vC=-1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010111; // iC= -937 
vC = 14'b1111101100100101; // vC=-1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000111; // iC= -889 
vC = 14'b1111101101001011; // vC=-1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101010; // iC= -918 
vC = 14'b1111101100000011; // vC=-1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110000; // iC= -976 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001011; // iC= -949 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000000; // iC= -832 
vC = 14'b1111101100100111; // vC=-1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b1111101101000110; // vC=-1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100111; // iC= -921 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000000; // iC= -832 
vC = 14'b1111101100011001; // vC=-1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000101; // iC= -891 
vC = 14'b1111101100001000; // vC=-1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100001; // iC= -863 
vC = 14'b1111101100010100; // vC=-1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000000; // iC= -960 
vC = 14'b1111101100001000; // vC=-1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101010; // iC= -918 
vC = 14'b1111101011110101; // vC=-1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010001; // iC= -943 
vC = 14'b1111101100101011; // vC=-1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111011; // iC= -901 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101011; // iC= -853 
vC = 14'b1111101100000100; // vC=-1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110001; // iC= -783 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010110; // iC= -874 
vC = 14'b1111101100101010; // vC=-1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011110; // iC= -802 
vC = 14'b1111101100101011; // vC=-1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110110; // iC= -842 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011011; // iC= -869 
vC = 14'b1111101010001010; // vC=-1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010100; // iC= -876 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100100; // iC= -796 
vC = 14'b1111101011011000; // vC=-1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011011; // iC= -805 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101000; // iC= -856 
vC = 14'b1111101011011110; // vC=-1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001011; // iC= -885 
vC = 14'b1111101100000011; // vC=-1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001100; // iC= -820 
vC = 14'b1111101011010101; // vC=-1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010110; // iC= -810 
vC = 14'b1111101001111100; // vC=-1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101101; // iC= -723 
vC = 14'b1111101011111000; // vC=-1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001101; // iC= -819 
vC = 14'b1111101010101110; // vC=-1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000011; // iC= -765 
vC = 14'b1111101011110001; // vC=-1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001101; // iC= -819 
vC = 14'b1111101001111011; // vC=-1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001110; // iC= -818 
vC = 14'b1111101010001001; // vC=-1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010011; // iC= -685 
vC = 14'b1111101011001000; // vC=-1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110100; // iC= -780 
vC = 14'b1111101011111010; // vC=-1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101010; // iC= -790 
vC = 14'b1111101011100101; // vC=-1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001010; // iC= -694 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010001; // iC= -815 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111111; // iC= -769 
vC = 14'b1111101010010101; // vC=-1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000000; // iC= -768 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001111; // iC= -689 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011011; // iC= -741 
vC = 14'b1111101010000010; // vC=-1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001001; // iC= -759 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010001; // iC= -751 
vC = 14'b1111101001011010; // vC=-1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011111; // iC= -673 
vC = 14'b1111101011100010; // vC=-1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011110; // iC= -610 
vC = 14'b1111101011010010; // vC=-1326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101010; // iC= -726 
vC = 14'b1111101001110100; // vC=-1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110110; // iC= -650 
vC = 14'b1111101011001011; // vC=-1333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010000; // iC= -752 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111000; // iC= -712 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100101; // iC= -731 
vC = 14'b1111101010000110; // vC=-1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111001; // iC= -711 
vC = 14'b1111101011010001; // vC=-1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101111; // iC= -593 
vC = 14'b1111101010111010; // vC=-1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000100; // iC= -700 
vC = 14'b1111101010100100; // vC=-1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111000; // iC= -712 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111101; // iC= -707 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001000; // iC= -696 
vC = 14'b1111101001001101; // vC=-1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101011; // iC= -661 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011100; // iC= -612 
vC = 14'b1111101001110101; // vC=-1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010110; // iC= -618 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011110; // iC= -674 
vC = 14'b1111101010000011; // vC=-1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101101; // iC= -595 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011111; // iC= -545 
vC = 14'b1111101001100100; // vC=-1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110111; // iC= -585 
vC = 14'b1111101000011100; // vC=-1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101010; // iC= -534 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000000; // iC= -640 
vC = 14'b1111101010001000; // vC=-1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110001; // iC= -527 
vC = 14'b1111101001101101; // vC=-1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010011; // iC= -621 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b1111101000110100; // vC=-1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000101; // iC= -507 
vC = 14'b1111101000001011; // vC=-1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101100; // iC= -596 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111110; // iC= -578 
vC = 14'b1111101010000010; // vC=-1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101110; // iC= -466 
vC = 14'b1111101000110100; // vC=-1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100110; // iC= -538 
vC = 14'b1111101000010110; // vC=-1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111111; // iC= -449 
vC = 14'b1111101001011001; // vC=-1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101010; // iC= -470 
vC = 14'b1111101000111001; // vC=-1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011100; // iC= -484 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101011; // iC= -533 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011110; // iC= -482 
vC = 14'b1111101000000000; // vC=-1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000010; // iC= -446 
vC = 14'b1111101001001001; // vC=-1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110011; // iC= -461 
vC = 14'b1111101000100101; // vC=-1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000111; // iC= -441 
vC = 14'b1111100111110110; // vC=-1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111101; // iC= -451 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011011; // iC= -485 
vC = 14'b1111101010000110; // vC=-1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100110; // iC= -410 
vC = 14'b1111101001010001; // vC=-1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001000; // iC= -504 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110011; // iC= -461 
vC = 14'b1111101000010001; // vC=-1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001010; // iC= -502 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001001; // iC= -503 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111110; // iC= -386 
vC = 14'b1111101010000011; // vC=-1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000110; // iC= -378 
vC = 14'b1111100111110111; // vC=-1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010010; // iC= -430 
vC = 14'b1111101001001111; // vC=-1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101110; // iC= -402 
vC = 14'b1111100111101111; // vC=-1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000101; // iC= -315 
vC = 14'b1111101001001101; // vC=-1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010101; // iC= -363 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100101; // iC= -411 
vC = 14'b1111101001001000; // vC=-1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100111; // iC= -409 
vC = 14'b1111101001101110; // vC=-1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000001; // iC= -255 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111001; // iC= -391 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000110; // iC= -378 
vC = 14'b1111101000110111; // vC=-1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101010; // iC= -342 
vC = 14'b1111101001000011; // vC=-1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111100; // iC= -260 
vC = 14'b1111101001010100; // vC=-1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011110; // iC= -226 
vC = 14'b1111101001001000; // vC=-1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100111; // iC= -281 
vC = 14'b1111100111011110; // vC=-1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010111; // iC= -297 
vC = 14'b1111101000110110; // vC=-1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001000; // iC= -184 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000010; // iC= -254 
vC = 14'b1111100111100101; // vC=-1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001000; // iC= -248 
vC = 14'b1111100111110010; // vC=-1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110011; // iC= -141 
vC = 14'b1111100111101001; // vC=-1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111001; // iC= -199 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101110; // iC=  -82 
vC = 14'b1111101001110010; // vC=-1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101111; // iC= -145 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101110; // iC=  -82 
vC = 14'b1111101000001011; // vC=-1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101010; // iC=  -86 
vC = 14'b1111101000110011; // vC=-1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001010; // iC=  -54 
vC = 14'b1111100111010001; // vC=-1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011101; // iC=  -35 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110011; // iC=  -13 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000100110; // iC=   38 
vC = 14'b1111100111111011; // vC=-1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101101; // iC=  -19 
vC = 14'b1111101001011000; // vC=-1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011100; // iC=  -36 
vC = 14'b1111100111110010; // vC=-1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101111; // iC=  -17 
vC = 14'b1111101000000010; // vC=-1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010000; // iC=   80 
vC = 14'b1111101001101100; // vC=-1428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101111; // iC=   47 
vC = 14'b1111101000011010; // vC=-1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000010; // iC=   66 
vC = 14'b1111101000000100; // vC=-1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100100; // iC=  100 
vC = 14'b1111101000000111; // vC=-1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000000; // iC=  128 
vC = 14'b1111101000100000; // vC=-1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110001; // iC=  177 
vC = 14'b1111101001100111; // vC=-1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000001; // iC=  129 
vC = 14'b1111100111110010; // vC=-1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000111; // iC=  135 
vC = 14'b1111101000101100; // vC=-1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010101; // iC=  277 
vC = 14'b1111101000011101; // vC=-1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010111; // iC=  215 
vC = 14'b1111100111010110; // vC=-1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111101; // iC=  189 
vC = 14'b1111101001001001; // vC=-1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001110; // iC=  206 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101011; // iC=  363 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100111; // iC=  295 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001100; // iC=  268 
vC = 14'b1111100111110111; // vC=-1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011011; // iC=  411 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000000; // iC=  448 
vC = 14'b1111100111110011; // vC=-1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001111; // iC=  399 
vC = 14'b1111101000111110; // vC=-1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101111; // iC=  367 
vC = 14'b1111101001110110; // vC=-1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001110; // iC=  462 
vC = 14'b1111100111110111; // vC=-1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111111; // iC=  447 
vC = 14'b1111100111101100; // vC=-1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001101; // iC=  461 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001100; // iC=  460 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110101; // iC=  629 
vC = 14'b1111101001110000; // vC=-1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110101; // iC=  565 
vC = 14'b1111100111111001; // vC=-1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001101; // iC=  589 
vC = 14'b1111101000000111; // vC=-1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101110; // iC=  558 
vC = 14'b1111101000000001; // vC=-1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000110; // iC=  646 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010001; // iC=  593 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101100; // iC=  684 
vC = 14'b1111101001100110; // vC=-1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111110; // iC=  766 
vC = 14'b1111101010010000; // vC=-1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101001; // iC=  681 
vC = 14'b1111101000111100; // vC=-1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101111; // iC=  687 
vC = 14'b1111101000010010; // vC=-1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010110; // iC=  854 
vC = 14'b1111101001110110; // vC=-1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011010; // iC=  794 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010100; // iC=  788 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001000; // iC=  840 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001010; // iC=  906 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b1111101001001110; // vC=-1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111110; // iC=  830 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100110; // iC=  934 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110111; // iC= 1015 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101001; // iC=  937 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110010; // iC= 1010 
vC = 14'b1111101000110111; // vC=-1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001010; // iC= 1034 
vC = 14'b1111101011000011; // vC=-1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001001; // iC= 1097 
vC = 14'b1111101001011010; // vC=-1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101001; // iC= 1129 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111100; // iC= 1084 
vC = 14'b1111101010011101; // vC=-1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011000; // iC= 1048 
vC = 14'b1111101001001001; // vC=-1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011101; // iC= 1117 
vC = 14'b1111101001000110; // vC=-1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100111; // iC= 1127 
vC = 14'b1111101011010101; // vC=-1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001011; // iC= 1099 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000001; // iC= 1153 
vC = 14'b1111101011000011; // vC=-1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011010; // iC= 1114 
vC = 14'b1111101010111100; // vC=-1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111110; // iC= 1214 
vC = 14'b1111101011000001; // vC=-1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010111; // iC= 1239 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110100; // iC= 1268 
vC = 14'b1111101010010111; // vC=-1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100001; // iC= 1313 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b1111101001100110; // vC=-1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100001; // iC= 1377 
vC = 14'b1111101100000001; // vC=-1279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010100; // iC= 1300 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010001; // iC= 1361 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011110; // iC= 1374 
vC = 14'b1111101011100100; // vC=-1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110001; // iC= 1393 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100101; // iC= 1445 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111110; // iC= 1406 
vC = 14'b1111101011111001; // vC=-1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011000; // iC= 1496 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011011; // iC= 1371 
vC = 14'b1111101011011110; // vC=-1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011111; // iC= 1503 
vC = 14'b1111101100011011; // vC=-1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111110; // iC= 1534 
vC = 14'b1111101011110101; // vC=-1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100000; // iC= 1504 
vC = 14'b1111101100000111; // vC=-1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110111; // iC= 1463 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111011; // iC= 1467 
vC = 14'b1111101011001011; // vC=-1333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110110; // iC= 1526 
vC = 14'b1111101100001100; // vC=-1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001111; // iC= 1615 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101100; // iC= 1580 
vC = 14'b1111101101000011; // vC=-1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101110; // iC= 1646 
vC = 14'b1111101100101000; // vC=-1240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001110; // iC= 1550 
vC = 14'b1111101100010110; // vC=-1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101111; // iC= 1519 
vC = 14'b1111101011101001; // vC=-1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100110; // iC= 1574 
vC = 14'b1111101100111010; // vC=-1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011001; // iC= 1561 
vC = 14'b1111101100010010; // vC=-1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100101; // iC= 1701 
vC = 14'b1111101100011001; // vC=-1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110110; // iC= 1654 
vC = 14'b1111101100000101; // vC=-1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001001; // iC= 1737 
vC = 14'b1111101100001101; // vC=-1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010000; // iC= 1616 
vC = 14'b1111101100000001; // vC=-1279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101101; // iC= 1709 
vC = 14'b1111101100111101; // vC=-1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b1111101110001011; // vC=-1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111111; // iC= 1663 
vC = 14'b1111101110001101; // vC=-1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110111; // iC= 1655 
vC = 14'b1111101101000000; // vC=-1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001001; // iC= 1737 
vC = 14'b1111101101100010; // vC=-1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000010; // iC= 1794 
vC = 14'b1111101101000000; // vC=-1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b1111101101100101; // vC=-1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b1111101100101111; // vC=-1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111010; // iC= 1786 
vC = 14'b1111101110001000; // vC=-1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001011; // iC= 1739 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011100; // iC= 1820 
vC = 14'b1111101101010000; // vC=-1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b1111101101100011; // vC=-1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b1111101101010100; // vC=-1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b1111101110110111; // vC=-1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000100; // iC= 1732 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b1111101110010101; // vC=-1131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100100; // iC= 1764 
vC = 14'b1111101110111110; // vC=-1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b1111101111101101; // vC=-1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111101110100101; // vC=-1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b1111101111010011; // vC=-1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b1111110000000011; // vC=-1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b1111101111100110; // vC=-1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111110000010100; // vC=-1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b1111101110011001; // vC=-1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b1111101110101100; // vC=-1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101010; // iC= 1898 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b1111101111101110; // vC=-1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b1111110000000100; // vC=-1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010011; // iC= 1811 
vC = 14'b1111101111110001; // vC=-1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b1111101111111010; // vC=-1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111101; // iC= 1853 
vC = 14'b1111110000100000; // vC= -992 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b1111110000111110; // vC= -962 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b1111101111011100; // vC=-1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b1111110000111100; // vC= -964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b1111101111101000; // vC=-1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b1111101111111010; // vC=-1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b1111110000101100; // vC= -980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b1111101111111011; // vC=-1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b1111110001111110; // vC= -898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011100; // iC= 1884 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111110010010110; // vC= -874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000010; // iC= 1858 
vC = 14'b1111110010101111; // vC= -849 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111110010011111; // vC= -865 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110001000011; // vC= -957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111110010001100; // vC= -884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111110011001100; // vC= -820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b1111110011011001; // vC= -807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111110011101110; // vC= -786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111110010011100; // vC= -868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001010; // iC= 1866 
vC = 14'b1111110010000000; // vC= -896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b1111110011100010; // vC= -798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000111; // iC= 1863 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111110011000110; // vC= -826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b1111110100000000; // vC= -768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b1111110100101010; // vC= -726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b1111110011001101; // vC= -819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b1111110011010101; // vC= -811 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b1111110100000100; // vC= -764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101100; // iC= 1964 
vC = 14'b1111110011001110; // vC= -818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b1111110101011111; // vC= -673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010100; // iC= 2004 
vC = 14'b1111110100011110; // vC= -738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111110101001110; // vC= -690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111110100110000; // vC= -720 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111110100101101; // vC= -723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111110100111000; // vC= -712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110100001100; // vC= -756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b1111110100100101; // vC= -731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111110110010110; // vC= -618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111110100110101; // vC= -715 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111110110010101; // vC= -619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101110; // iC= 2030 
vC = 14'b1111110110011110; // vC= -610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111110111001111; // vC= -561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110101000101; // vC= -699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111110101001011; // vC= -693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111110110101000; // vC= -600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111111; // iC= 2047 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111110110111011; // vC= -581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111110110011101; // vC= -611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111110111110011; // vC= -525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111110110011110; // vC= -610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110010; // iC= 2034 
vC = 14'b1111110111110011; // vC= -525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110111; // iC= 1975 
vC = 14'b1111111000010011; // vC= -493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101110; // iC= 2030 
vC = 14'b1111110110100011; // vC= -605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101110; // iC= 2030 
vC = 14'b1111110111111101; // vC= -515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111110110100111; // vC= -601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b1111110111010100; // vC= -556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010000; // iC= 2064 
vC = 14'b1111110111111000; // vC= -520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111110111111001; // vC= -519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111110110101111; // vC= -593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111110110110010; // vC= -590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111001; // iC= 2041 
vC = 14'b1111110111100000; // vC= -544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111111000100010; // vC= -478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000100; // iC= 2052 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b1111110111010001; // vC= -559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b1111110111110000; // vC= -528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111110111111101; // vC= -515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111110111100000; // vC= -544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b1111111000011001; // vC= -487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111111000101000; // vC= -472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011101; // iC= 2013 
vC = 14'b1111111001111101; // vC= -387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111111001110100; // vC= -396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b1111110111111011; // vC= -517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b1111111000110110; // vC= -458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b1111111001100110; // vC= -410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011000; // iC= 2072 
vC = 14'b1111111000010101; // vC= -491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b1111111000110011; // vC= -461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111010100000; // vC= -352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111111001011101; // vC= -419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001101; // iC= 2061 
vC = 14'b1111111001100111; // vC= -409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000100; // iC= 2052 
vC = 14'b1111111010111000; // vC= -328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111111001011101; // vC= -419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001100; // iC= 2060 
vC = 14'b1111111010000110; // vC= -378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111111011100010; // vC= -286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111010110001; // vC= -335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000000; // iC= 1984 
vC = 14'b1111111011011001; // vC= -295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111111001110001; // vC= -399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111111010001010; // vC= -374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b1111111010100110; // vC= -346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010110; // iC= 2070 
vC = 14'b1111111011001000; // vC= -312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010111; // iC= 2071 
vC = 14'b1111111011111001; // vC= -263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000101; // iC= 2053 
vC = 14'b1111111010111010; // vC= -326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b1111111100011001; // vC= -231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101110; // iC= 2030 
vC = 14'b1111111011001101; // vC= -307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111111100111101; // vC= -195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011011; // iC= 2011 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b1111111100110001; // vC= -207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111111011011100; // vC= -292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111110; // iC= 1982 
vC = 14'b1111111101011110; // vC= -162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101011; // iC= 2027 
vC = 14'b1111111011111111; // vC= -257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b1111111100110110; // vC= -202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111111100000000; // vC= -256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111111101000001; // vC= -191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b1111111101111010; // vC= -134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111111101110100; // vC= -140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111111101101101; // vC= -147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111111100101110; // vC= -210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100010; // iC= 2018 
vC = 14'b1111111100000111; // vC= -249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111111100111010; // vC= -198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111111110100100; // vC=  -92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100011; // iC= 2019 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111111101111101; // vC= -131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001101; // iC= 2061 
vC = 14'b1111111110010011; // vC= -109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111101000001; // vC= -191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111101110010; // vC= -142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111111101100100; // vC= -156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111111000100; // vC=  -60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111111110010001; // vC= -111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b1111111110011111; // vC=  -97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110111; // iC= 1975 
vC = 14'b1111111101111010; // vC= -134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b1111111110101101; // vC=  -83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b1111111101100001; // vC= -159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b1111111111000001; // vC=  -63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111111111111111; // vC=   -1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100101; // iC= 2021 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b1111111111111101; // vC=   -3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b0000000000010001; // vC=   17 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b1111111111101001; // vC=  -23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b0000000000010010; // vC=   18 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111111111000010; // vC=  -62 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111111111100101; // vC=  -27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b0000000000100111; // vC=   39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111111111001111; // vC=  -49 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001010; // iC= 1994 
vC = 14'b0000000000110111; // vC=   55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111110110110; // vC=  -74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b1111111110111001; // vC=  -71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b0000000000101111; // vC=   47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110111; // iC= 1975 
vC = 14'b1111111111001010; // vC=  -54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111111111001101; // vC=  -51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b0000000000011011; // vC=   27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011001; // iC= 1881 
vC = 14'b0000000000000101; // vC=    5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100010; // iC= 2018 
vC = 14'b0000000000101110; // vC=   46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b0000000010001001; // vC=  137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011110; // iC= 1886 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b0000000000001110; // vC=   14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101100; // iC= 1964 
vC = 14'b0000000000110101; // vC=   53 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b0000000010000110; // vC=  134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b0000000010100011; // vC=  163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b0000000010110111; // vC=  183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b0000000001110110; // vC=  118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b0000000001101010; // vC=  106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b0000000010001001; // vC=  137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b0000000011011100; // vC=  220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b0000000011110000; // vC=  240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b0000000010000011; // vC=  131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b0000000010100110; // vC=  166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b0000000100101011; // vC=  299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b0000000010101101; // vC=  173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001010; // iC= 1866 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b0000000010111100; // vC=  188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b0000000011100100; // vC=  228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b0000000011100000; // vC=  224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b0000000100011101; // vC=  285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b0000000101000100; // vC=  324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000011; // iC= 1859 
vC = 14'b0000000011101010; // vC=  234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b0000000011101001; // vC=  233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000000011101000; // vC=  232 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b0000000101000010; // vC=  322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b0000000101011100; // vC=  348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b0000000100101101; // vC=  301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110010; // iC= 1906 
vC = 14'b0000000100010010; // vC=  274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b0000000101000100; // vC=  324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b0000000110000001; // vC=  385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b0000000100010100; // vC=  276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b0000000100101010; // vC=  298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b0000000101100000; // vC=  352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000000110010111; // vC=  407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b0000000101101100; // vC=  364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b0000000110111110; // vC=  446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b0000000110011101; // vC=  413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b0000000111100000; // vC=  480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101110; // iC= 1838 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110010; // iC= 1778 
vC = 14'b0000000110000100; // vC=  388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100011; // iC= 1827 
vC = 14'b0000000101011101; // vC=  349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b0000000111010000; // vC=  464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b0000000101101010; // vC=  362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b0000000110011111; // vC=  415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b0000000111110111; // vC=  503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100110; // iC= 1830 
vC = 14'b0000000111100011; // vC=  483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b0000000110010000; // vC=  400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b0000001000000000; // vC=  512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b0000000110011101; // vC=  413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b0000000110011011; // vC=  411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b0000000110101011; // vC=  427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110101; // iC= 1781 
vC = 14'b0000001000101011; // vC=  555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b0000001000011110; // vC=  542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010011; // iC= 1747 
vC = 14'b0000001000100000; // vC=  544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b0000000111101111; // vC=  495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001000; // iC= 1864 
vC = 14'b0000000111000000; // vC=  448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b0000001000011100; // vC=  540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b0000001000101000; // vC=  552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b0000001000111101; // vC=  573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000110; // iC= 1734 
vC = 14'b0000000111010111; // vC=  471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b0000001001011110; // vC=  606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b0000001001100110; // vC=  614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111001; // iC= 1849 
vC = 14'b0000001010000001; // vC=  641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000001000001111; // vC=  527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101110; // iC= 1710 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000001001011100; // vC=  604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b0000001001101010; // vC=  618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b0000001001101110; // vC=  622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b0000001001001110; // vC=  590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b0000001001010011; // vC=  595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111110; // iC= 1726 
vC = 14'b0000001001011101; // vC=  605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b0000001000101100; // vC=  556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b0000001010100110; // vC=  678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011111; // iC= 1759 
vC = 14'b0000001010111010; // vC=  698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011011; // iC= 1755 
vC = 14'b0000001001001010; // vC=  586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b0000001010011000; // vC=  664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b0000001010110000; // vC=  688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011000; // iC= 1688 
vC = 14'b0000001011000101; // vC=  709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b0000001001111011; // vC=  635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000000; // iC= 1664 
vC = 14'b0000001001101001; // vC=  617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000001011111011; // vC=  763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001110; // iC= 1678 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b0000001011110101; // vC=  757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b0000001010100101; // vC=  677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b0000001011011111; // vC=  735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b0000001010011111; // vC=  671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b0000001010101111; // vC=  687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b0000001100010101; // vC=  789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b0000001010101100; // vC=  684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b0000001010111101; // vC=  701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100111; // iC= 1639 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b0000001010110001; // vC=  689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b0000001100111100; // vC=  828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010100; // iC= 1620 
vC = 14'b0000001010110111; // vC=  695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000111; // iC= 1607 
vC = 14'b0000001100101010; // vC=  810 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101110; // iC= 1710 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b0000001100100010; // vC=  802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b0000001100000010; // vC=  770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010010; // iC= 1618 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101100; // iC= 1580 
vC = 14'b0000001101001110; // vC=  846 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101001; // iC= 1705 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b0000001110000000; // vC=  896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b0000001101101111; // vC=  879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b0000001100111010; // vC=  826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101010; // iC= 1578 
vC = 14'b0000001101011010; // vC=  858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b0000001101011111; // vC=  863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b0000001100110111; // vC=  823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b0000001100001111; // vC=  783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b0000001110010111; // vC=  919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110101; // iC= 1653 
vC = 14'b0000001110101010; // vC=  938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b0000001100111111; // vC=  831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011110; // iC= 1566 
vC = 14'b0000001110100000; // vC=  928 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100111; // iC= 1639 
vC = 14'b0000001101011111; // vC=  863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101101; // iC= 1645 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100100; // iC= 1636 
vC = 14'b0000001110101001; // vC=  937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111000; // iC= 1592 
vC = 14'b0000001101100010; // vC=  866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010000; // iC= 1552 
vC = 14'b0000001101011110; // vC=  862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100011; // iC= 1507 
vC = 14'b0000001101011010; // vC=  858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111110; // iC= 1534 
vC = 14'b0000001110000000; // vC=  896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b0000001110000110; // vC=  902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101011; // iC= 1515 
vC = 14'b0000001110001101; // vC=  909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101100; // iC= 1580 
vC = 14'b0000001101010010; // vC=  850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011010; // iC= 1626 
vC = 14'b0000001110000010; // vC=  898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101010; // iC= 1642 
vC = 14'b0000001111000101; // vC=  965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011010; // iC= 1562 
vC = 14'b0000001110011001; // vC=  921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011010; // iC= 1498 
vC = 14'b0000001110000010; // vC=  898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001001; // iC= 1609 
vC = 14'b0000001111111110; // vC= 1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011001; // iC= 1497 
vC = 14'b0000001111100101; // vC=  997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110001; // iC= 1585 
vC = 14'b0000001111010111; // vC=  983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110100; // iC= 1460 
vC = 14'b0000010000010100; // vC= 1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000001110001101; // vC=  909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110111; // iC= 1527 
vC = 14'b0000010000000010; // vC= 1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101111; // iC= 1455 
vC = 14'b0000001110101101; // vC=  941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000001; // iC= 1473 
vC = 14'b0000010000001001; // vC= 1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100110; // iC= 1574 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101010; // iC= 1578 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110000; // iC= 1584 
vC = 14'b0000010000010001; // vC= 1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011010; // iC= 1498 
vC = 14'b0000001111010011; // vC=  979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011010; // iC= 1562 
vC = 14'b0000001110101111; // vC=  943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000001111000010; // vC=  962 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011010; // iC= 1498 
vC = 14'b0000001111111010; // vC= 1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111111; // iC= 1407 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100010; // iC= 1506 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000010000111011; // vC= 1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110100; // iC= 1396 
vC = 14'b0000001111010100; // vC=  980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000111; // iC= 1479 
vC = 14'b0000010001011111; // vC= 1119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100101; // iC= 1445 
vC = 14'b0000001111100010; // vC=  994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011111; // iC= 1439 
vC = 14'b0000010000100001; // vC= 1057 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000011; // iC= 1411 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000101; // iC= 1477 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b0000001111101011; // vC= 1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101100; // iC= 1388 
vC = 14'b0000010001011100; // vC= 1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100010; // iC= 1442 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000010; // iC= 1474 
vC = 14'b0000001111110101; // vC= 1013 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110101; // iC= 1397 
vC = 14'b0000001111110110; // vC= 1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000111; // iC= 1351 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000010; // iC= 1474 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010001; // iC= 1361 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b0000010010000001; // vC= 1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010010; // iC= 1426 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001100; // iC= 1356 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000011; // iC= 1347 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010001; // iC= 1425 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001001; // iC= 1353 
vC = 14'b0000010010101001; // vC= 1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100010; // iC= 1378 
vC = 14'b0000010000111001; // vC= 1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000000; // iC= 1408 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011111; // iC= 1311 
vC = 14'b0000010010010101; // vC= 1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111010; // iC= 1338 
vC = 14'b0000010000101011; // vC= 1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011100; // iC= 1372 
vC = 14'b0000010011000011; // vC= 1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101001; // iC= 1321 
vC = 14'b0000010010111111; // vC= 1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110110; // iC= 1334 
vC = 14'b0000010010101000; // vC= 1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111100; // iC= 1404 
vC = 14'b0000010001101110; // vC= 1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100100; // iC= 1316 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101001; // iC= 1385 
vC = 14'b0000010010001011; // vC= 1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001010; // iC= 1418 
vC = 14'b0000010001010001; // vC= 1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110001; // iC= 1393 
vC = 14'b0000010011101000; // vC= 1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111110; // iC= 1342 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010111; // iC= 1367 
vC = 14'b0000010011000000; // vC= 1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001111; // iC= 1359 
vC = 14'b0000010011010111; // vC= 1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010011; // iC= 1363 
vC = 14'b0000010010101001; // vC= 1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010100; // iC= 1364 
vC = 14'b0000010010100001; // vC= 1185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000100; // iC= 1348 
vC = 14'b0000010011001001; // vC= 1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011000; // iC= 1368 
vC = 14'b0000010010011001; // vC= 1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010010; // iC= 1234 
vC = 14'b0000010010111000; // vC= 1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001111; // iC= 1295 
vC = 14'b0000010011011100; // vC= 1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110000; // iC= 1264 
vC = 14'b0000010010100000; // vC= 1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111010; // iC= 1274 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000010100000011; // vC= 1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100011; // iC= 1251 
vC = 14'b0000010011000000; // vC= 1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001111; // iC= 1295 
vC = 14'b0000010010001101; // vC= 1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001011; // iC= 1291 
vC = 14'b0000010100100010; // vC= 1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110010; // iC= 1266 
vC = 14'b0000010100101101; // vC= 1325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111111; // iC= 1279 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000010011001111; // vC= 1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100011; // iC= 1187 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010001; // iC= 1169 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001010; // iC= 1226 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011000; // iC= 1176 
vC = 14'b0000010011100011; // vC= 1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110111; // iC= 1271 
vC = 14'b0000010011100110; // vC= 1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010110; // iC= 1302 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111001; // iC= 1145 
vC = 14'b0000010011010100; // vC= 1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000010; // iC= 1282 
vC = 14'b0000010101001001; // vC= 1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001110; // iC= 1230 
vC = 14'b0000010100000101; // vC= 1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001011; // iC= 1163 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111000; // iC= 1208 
vC = 14'b0000010100111111; // vC= 1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011101; // iC= 1117 
vC = 14'b0000010100011110; // vC= 1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010110; // iC= 1110 
vC = 14'b0000010011010010; // vC= 1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100101; // iC= 1125 
vC = 14'b0000010100001111; // vC= 1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111011; // iC= 1147 
vC = 14'b0000010101101101; // vC= 1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110010; // iC= 1202 
vC = 14'b0000010101001101; // vC= 1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001010; // iC= 1162 
vC = 14'b0000010100100100; // vC= 1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111000; // iC= 1144 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100101; // iC= 1189 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001111; // iC= 1103 
vC = 14'b0000010100110010; // vC= 1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010100; // iC= 1172 
vC = 14'b0000010011101100; // vC= 1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011111; // iC= 1183 
vC = 14'b0000010011101010; // vC= 1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111010; // iC= 1146 
vC = 14'b0000010100101101; // vC= 1325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100001; // iC= 1185 
vC = 14'b0000010100001010; // vC= 1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111010; // iC= 1082 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001111; // iC= 1039 
vC = 14'b0000010100110011; // vC= 1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101001; // iC= 1065 
vC = 14'b0000010100001111; // vC= 1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001010; // iC= 1034 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010000; // iC= 1040 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010001; // iC= 1105 
vC = 14'b0000010101001110; // vC= 1358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110001; // iC= 1137 
vC = 14'b0000010100000101; // vC= 1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000101; // iC= 1093 
vC = 14'b0000010100110110; // vC= 1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110010; // iC= 1074 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101000; // iC= 1064 
vC = 14'b0000010110011010; // vC= 1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100110; // iC=  998 
vC = 14'b0000010100011101; // vC= 1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111010; // iC= 1082 
vC = 14'b0000010100110010; // vC= 1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101111; // iC= 1007 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111001; // iC= 1017 
vC = 14'b0000010100011100; // vC= 1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010100; // iC= 1044 
vC = 14'b0000010100101010; // vC= 1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101100; // iC= 1068 
vC = 14'b0000010110011110; // vC= 1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010110; // iC=  982 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111000; // iC= 1080 
vC = 14'b0000010101001001; // vC= 1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000010; // iC= 1090 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011010; // iC=  986 
vC = 14'b0000010101010001; // vC= 1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000111; // iC= 1031 
vC = 14'b0000010110001010; // vC= 1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001100; // iC= 1036 
vC = 14'b0000010101111101; // vC= 1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110111; // iC= 1079 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111010; // iC=  954 
vC = 14'b0000010110011110; // vC= 1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011110; // iC=  990 
vC = 14'b0000010101101011; // vC= 1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010000; // iC=  976 
vC = 14'b0000010111011000; // vC= 1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100001; // iC=  993 
vC = 14'b0000010110111111; // vC= 1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001111; // iC=  911 
vC = 14'b0000010111010000; // vC= 1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100000; // iC=  992 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101010; // iC=  938 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101001; // iC= 1001 
vC = 14'b0000010110010001; // vC= 1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001010; // iC=  906 
vC = 14'b0000010111011011; // vC= 1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001111; // iC=  911 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011010; // iC=  986 
vC = 14'b0000010110101001; // vC= 1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000001; // iC= 1025 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100000; // iC=  992 
vC = 14'b0000010111011101; // vC= 1501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110011; // iC=  947 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111011; // iC=  891 
vC = 14'b0000010110010110; // vC= 1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010010; // iC=  978 
vC = 14'b0000010110100101; // vC= 1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110110; // iC=  886 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000110; // iC=  966 
vC = 14'b0000010111001011; // vC= 1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011101; // iC=  861 
vC = 14'b0000010110001000; // vC= 1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001100; // iC=  972 
vC = 14'b0000010110000101; // vC= 1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010000; // iC=  912 
vC = 14'b0000010111000100; // vC= 1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111010; // iC=  954 
vC = 14'b0000010110111010; // vC= 1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000011; // iC=  963 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100011; // iC=  867 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000010; // iC=  834 
vC = 14'b0000011000001001; // vC= 1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000011; // iC=  835 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111100; // iC=  892 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011111; // iC=  863 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110010; // iC=  818 
vC = 14'b0000010111100111; // vC= 1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010011; // iC=  915 
vC = 14'b0000010111001010; // vC= 1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001010; // iC=  778 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111100; // iC=  764 
vC = 14'b0000010110011010; // vC= 1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110010; // iC=  818 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110000; // iC=  880 
vC = 14'b0000010111000011; // vC= 1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110000; // iC=  880 
vC = 14'b0000010110010111; // vC= 1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011011; // iC=  795 
vC = 14'b0000010110111101; // vC= 1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110101; // iC=  757 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110000; // iC=  880 
vC = 14'b0000010111010000; // vC= 1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111010; // iC=  762 
vC = 14'b0000011000111101; // vC= 1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110001; // iC=  817 
vC = 14'b0000011000101010; // vC= 1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100011; // iC=  739 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000111; // iC=  711 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010010; // iC=  786 
vC = 14'b0000010111110101; // vC= 1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000110; // iC=  774 
vC = 14'b0000010111101100; // vC= 1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001001; // iC=  777 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000111; // iC=  775 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100001; // iC=  673 
vC = 14'b0000011001000000; // vC= 1600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010010; // iC=  786 
vC = 14'b0000010111001111; // vC= 1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100001; // iC=  673 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011000; // iC=  728 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101111; // iC=  687 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001101; // iC=  653 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000000; // iC=  768 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010111; // iC=  663 
vC = 14'b0000010111010110; // vC= 1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011001; // iC=  729 
vC = 14'b0000010111000010; // vC= 1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110110; // iC=  758 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000111; // iC=  647 
vC = 14'b0000010111111110; // vC= 1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000000; // iC=  640 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011011; // iC=  603 
vC = 14'b0000011001011101; // vC= 1629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000100; // iC=  708 
vC = 14'b0000011000101000; // vC= 1576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010001; // iC=  593 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010011; // iC=  723 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101111; // iC=  623 
vC = 14'b0000011001011000; // vC= 1624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100001; // iC=  673 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011100; // iC=  604 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001000; // iC=  648 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001011; // iC=  587 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111011; // iC=  571 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100010; // iC=  546 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100011; // iC=  611 
vC = 14'b0000011000101111; // vC= 1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111111; // iC=  639 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110111; // iC=  567 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111110; // iC=  574 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110000; // iC=  560 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110000; // iC=  624 
vC = 14'b0000011000010010; // vC= 1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111111; // iC=  511 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101000; // iC=  552 
vC = 14'b0000011000101111; // vC= 1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001110; // iC=  526 
vC = 14'b0000011010000000; // vC= 1664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100101; // iC=  485 
vC = 14'b0000011001000000; // vC= 1600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101000; // iC=  616 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110111; // iC=  567 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010011; // iC=  531 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110000; // iC=  560 
vC = 14'b0000011001100111; // vC= 1639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110011; // iC=  563 
vC = 14'b0000011001111100; // vC= 1660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100001; // iC=  481 
vC = 14'b0000011001100110; // vC= 1638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001101; // iC=  461 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100011; // iC=  547 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101111; // iC=  495 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001110; // iC=  526 
vC = 14'b0000011000011001; // vC= 1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011100; // iC=  412 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110000; // iC=  432 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101110; // iC=  494 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001100; // iC=  460 
vC = 14'b0000011001001110; // vC= 1614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100101; // iC=  357 
vC = 14'b0000011010000000; // vC= 1664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000010; // iC=  450 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001111; // iC=  335 
vC = 14'b0000011010010111; // vC= 1687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010011; // iC=  467 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110111; // iC=  311 
vC = 14'b0000011001100111; // vC= 1639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100000; // iC=  352 
vC = 14'b0000011001111010; // vC= 1658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001100; // iC=  332 
vC = 14'b0000011000010011; // vC= 1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010111; // iC=  279 
vC = 14'b0000011010001110; // vC= 1678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101000; // iC=  360 
vC = 14'b0000011001111111; // vC= 1663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000000; // iC=  320 
vC = 14'b0000011001111100; // vC= 1660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101100; // iC=  300 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001010; // iC=  330 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100001; // iC=  353 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110100; // iC=  244 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010011; // iC=  275 
vC = 14'b0000011010001101; // vC= 1677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010111; // iC=  215 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101010; // iC=  170 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010101111; // iC=  175 
vC = 14'b0000011010000001; // vC= 1665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110101; // iC=  181 
vC = 14'b0000011000001101; // vC= 1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000011; // iC=  195 
vC = 14'b0000011001111011; // vC= 1659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001110; // iC=   78 
vC = 14'b0000011000110001; // vC= 1585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001101; // iC=   77 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000011; // iC=  131 
vC = 14'b0000011010000100; // vC= 1668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111111; // iC=   63 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111100; // iC=   60 
vC = 14'b0000011010000001; // vC= 1665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100111; // iC=  103 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110011; // iC=  -13 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011010; // iC=   90 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100101; // iC=  -27 
vC = 14'b0000011001111011; // vC= 1659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110010; // iC=  -14 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011110; // iC=   30 
vC = 14'b0000011010000101; // vC= 1669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100110; // iC=  -90 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110000; // iC= -144 
vC = 14'b0000011000111110; // vC= 1598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100011; // iC=  -93 
vC = 14'b0000011010010011; // vC= 1683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011110; // iC= -162 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111100; // iC=  -68 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110100; // iC= -140 
vC = 14'b0000010111111110; // vC= 1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000011; // iC= -125 
vC = 14'b0000011001110110; // vC= 1654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111110; // iC= -194 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110100; // iC= -204 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001011; // iC= -309 
vC = 14'b0000011000110110; // vC= 1590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000110; // iC= -314 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000101; // iC= -315 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111100; // iC= -260 
vC = 14'b0000011010001011; // vC= 1675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001110; // iC= -370 
vC = 14'b0000011010000010; // vC= 1666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101101; // iC= -403 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001010; // iC= -310 
vC = 14'b0000011001101111; // vC= 1647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011001; // iC= -423 
vC = 14'b0000011001110110; // vC= 1654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011000; // iC= -360 
vC = 14'b0000010111100110; // vC= 1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010100; // iC= -492 
vC = 14'b0000010111101010; // vC= 1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110000; // iC= -528 
vC = 14'b0000011001101010; // vC= 1642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010010; // iC= -430 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111001; // iC= -519 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101010; // iC= -470 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111100; // iC= -580 
vC = 14'b0000010111111101; // vC= 1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110010; // iC= -526 
vC = 14'b0000010111110100; // vC= 1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100100; // iC= -604 
vC = 14'b0000010111101011; // vC= 1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011110; // iC= -546 
vC = 14'b0000011000011001; // vC= 1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101101; // iC= -659 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011111; // iC= -737 
vC = 14'b0000010111110101; // vC= 1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010011; // iC= -685 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100101; // iC= -731 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110010; // iC= -654 
vC = 14'b0000010111111111; // vC= 1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011000; // iC= -744 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000100; // iC= -700 
vC = 14'b0000011001010001; // vC= 1617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010000; // iC= -816 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001111; // iC= -753 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110111; // iC= -905 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101010; // iC= -790 
vC = 14'b0000010111100110; // vC= 1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100110; // iC= -794 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000100; // iC= -892 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011000; // iC= -872 
vC = 14'b0000010110111101; // vC= 1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101100; // iC= -980 
vC = 14'b0000010110110011; // vC= 1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111101; // iC= -899 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001010; // iC= -950 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b0000011000101010; // vC= 1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101011; // iC= -981 
vC = 14'b0000010110001111; // vC= 1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111010; // iC= -966 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011111; // iC=-1121 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010010; // iC=-1070 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010010; // iC=-1006 
vC = 14'b0000010110010010; // vC= 1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001001; // iC=-1143 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101000; // iC=-1176 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010100; // iC=-1196 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001010; // iC=-1078 
vC = 14'b0000010101111000; // vC= 1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100111; // iC=-1177 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101000; // iC=-1240 
vC = 14'b0000010110000001; // vC= 1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001010; // iC=-1206 
vC = 14'b0000010111001111; // vC= 1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010010; // iC=-1198 
vC = 14'b0000010111101010; // vC= 1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110111; // iC=-1289 
vC = 14'b0000010111000010; // vC= 1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000110; // iC=-1210 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b0000010110000101; // vC= 1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100010; // iC=-1246 
vC = 14'b0000010101110010; // vC= 1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110110; // iC=-1290 
vC = 14'b0000010100111111; // vC= 1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101001; // iC=-1239 
vC = 14'b0000010101010001; // vC= 1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011000; // iC=-1320 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110110; // iC=-1354 
vC = 14'b0000010111000011; // vC= 1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010001; // iC=-1327 
vC = 14'b0000010101100000; // vC= 1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000111; // iC=-1401 
vC = 14'b0000010101111100; // vC= 1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110011; // iC=-1421 
vC = 14'b0000010100111111; // vC= 1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101001; // iC=-1367 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b0000010101010011; // vC= 1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101011; // iC=-1365 
vC = 14'b0000010101110010; // vC= 1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000010100111111; // vC= 1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b0000010110011000; // vC= 1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001011; // iC=-1461 
vC = 14'b0000010100111011; // vC= 1339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011001; // iC=-1511 
vC = 14'b0000010101110010; // vC= 1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b0000010101110001; // vC= 1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b0000010100011101; // vC= 1309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110010; // iC=-1486 
vC = 14'b0000010011111111; // vC= 1279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b0000010101011001; // vC= 1369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000010; // iC=-1470 
vC = 14'b0000010100000001; // vC= 1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000010100011110; // vC= 1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110010; // iC=-1486 
vC = 14'b0000010100101001; // vC= 1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b0000010011011001; // vC= 1241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010111; // iC=-1513 
vC = 14'b0000010011101000; // vC= 1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001101; // iC=-1587 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110100; // iC=-1548 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b0000010011101100; // vC= 1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b0000010010110110; // vC= 1206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001101; // iC=-1587 
vC = 14'b0000010010110111; // vC= 1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b0000010011100110; // vC= 1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000010010110110; // vC= 1206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011110; // iC=-1698 
vC = 14'b0000010011010010; // vC= 1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b0000010011000111; // vC= 1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b0000010010000011; // vC= 1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b0000010011100101; // vC= 1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000010010001001; // vC= 1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011010; // iC=-1702 
vC = 14'b0000010010011001; // vC= 1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b0000010000101111; // vC= 1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000010010000010; // vC= 1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001010; // iC=-1654 
vC = 14'b0000010001011010; // vC= 1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000010010010011; // vC= 1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b0000010000101010; // vC= 1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100101; // iC=-1627 
vC = 14'b0000010010000100; // vC= 1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000001111111100; // vC= 1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b0000010001111000; // vC= 1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001111; // iC=-1649 
vC = 14'b0000001111111011; // vC= 1019 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b0000010000100000; // vC= 1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000001110111100; // vC=  956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010010; // iC=-1646 
vC = 14'b0000001111101100; // vC= 1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001111100110; // vC=  998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100101; // iC=-1691 
vC = 14'b0000010000000000; // vC= 1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b0000001111010111; // vC=  983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000001111001001; // vC=  969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b0000001110110011; // vC=  947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000001110100001; // vC=  929 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b0000001111100100; // vC=  996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000010000000000; // vC= 1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b0000001110010000; // vC=  912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b0000001111010100; // vC=  980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100101; // iC=-1691 
vC = 14'b0000001110010101; // vC=  917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000001101011101; // vC=  861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000001111010101; // vC=  981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000001101100000; // vC=  864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b0000001101011000; // vC=  856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000001100111011; // vC=  827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000001110110101; // vC=  949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110010; // iC=-1806 
vC = 14'b0000001110111001; // vC=  953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b0000001101111011; // vC=  891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100000; // iC=-1824 
vC = 14'b0000001100110110; // vC=  822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000001110010100; // vC=  916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b0000001100001111; // vC=  783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000001101011111; // vC=  863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000001101110111; // vC=  887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000001101110010; // vC=  882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000001101011111; // vC=  863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000001011100011; // vC=  739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000001100000101; // vC=  773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000001100001110; // vC=  782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000001100101001; // vC=  809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b0000001100000101; // vC=  773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000001011111010; // vC=  762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b0000001100010100; // vC=  788 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b0000001100101001; // vC=  809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011010; // iC=-1830 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000001100001001; // vC=  777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001100011010; // vC=  794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000001100011010; // vC=  794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111011; // iC=-1797 
vC = 14'b0000001011101001; // vC=  745 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000001011101101; // vC=  749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b0000001001111010; // vC=  634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000001010010011; // vC=  659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000001001101101; // vC=  621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000001011010110; // vC=  726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000001010101101; // vC=  685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001010010010; // vC=  658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000001000111100; // vC=  572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101000; // iC=-1880 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000001001000001; // vC=  577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000001010110001; // vC=  689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000001000111101; // vC=  573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000001000110000; // vC=  560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111011; // iC=-1797 
vC = 14'b0000001001010101; // vC=  597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000001000111101; // vC=  573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b0000001000000000; // vC=  512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110100; // iC=-1868 
vC = 14'b0000001001110110; // vC=  630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100101; // iC=-1883 
vC = 14'b0000001001011111; // vC=  607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000001001100000; // vC=  608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000001000010101; // vC=  533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b0000001001010110; // vC=  598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011010; // iC=-1830 
vC = 14'b0000001001011110; // vC=  606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000001001100101; // vC=  613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100000; // iC=-1888 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000000111010101; // vC=  469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000000111101110; // vC=  494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b0000001001001000; // vC=  584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000000111000001; // vC=  449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000001000100100; // vC=  548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110000; // iC=-1872 
vC = 14'b0000000110110111; // vC=  439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000000111000101; // vC=  453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000000111100010; // vC=  482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110100; // iC=-1868 
vC = 14'b0000000110101101; // vC=  429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110010; // iC=-1806 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000000111111111; // vC=  511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000011; // iC=-1853 
vC = 14'b0000000111011000; // vC=  472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b0000000110000110; // vC=  390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b0000000110010101; // vC=  405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000000101100111; // vC=  359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b0000000101001001; // vC=  329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b0000000111000101; // vC=  453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001111; // iC=-1841 
vC = 14'b0000000101100110; // vC=  358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000000101001101; // vC=  333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000000101100111; // vC=  359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100110; // iC=-1882 
vC = 14'b0000000101011010; // vC=  346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000000100111110; // vC=  318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000000100100010; // vC=  290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000000100111000; // vC=  312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b0000000101111001; // vC=  377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000000101000110; // vC=  326 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111101; // iC=-1859 
vC = 14'b0000000101000010; // vC=  322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101100; // iC=-1876 
vC = 14'b0000000100101101; // vC=  301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111001; // iC=-1863 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000000101001101; // vC=  333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000000101101101; // vC=  365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000000100100101; // vC=  293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101011; // iC=-1877 
vC = 14'b0000000011011111; // vC=  223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b0000000101001010; // vC=  330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111010; // iC=-1862 
vC = 14'b0000000100010001; // vC=  273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b0000000100000000; // vC=  256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000000011011111; // vC=  223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000000100000011; // vC=  259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010000; // iC=-1840 
vC = 14'b0000000101000011; // vC=  323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b0000000010110000; // vC=  176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000000010110111; // vC=  183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101110; // iC=-1874 
vC = 14'b0000000011101110; // vC=  238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000000100100001; // vC=  289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000000100000011; // vC=  259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000000011010111; // vC=  215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000000001100101; // vC=  101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101011; // iC=-1877 
vC = 14'b0000000011001111; // vC=  207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b0000000011001100; // vC=  204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000000010101001; // vC=  169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000010001001; // vC=  137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000000001011000; // vC=   88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010000; // iC=-1840 
vC = 14'b0000000010001100; // vC=  140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000000; // iC=-1792 
vC = 14'b0000000001101011; // vC=  107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000000010100110; // vC=  166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000000001101010; // vC=  106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b0000000010100000; // vC=  160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000010001110; // vC=  142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b0000000010001011; // vC=  139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000000000111111; // vC=   63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010011; // iC=-1837 
vC = 14'b0000000000101001; // vC=   41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100110; // iC=-1754 
vC = 14'b0000000000100010; // vC=   34 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b1111111111011101; // vC=  -35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b1111111111000110; // vC=  -58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000000001010111; // vC=   87 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b1111111111100011; // vC=  -29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001011; // iC=-1845 
vC = 14'b1111111111111111; // vC=   -1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b0000000000001000; // vC=    8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b0000000000011110; // vC=   30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b1111111110101011; // vC=  -85 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b1111111110011011; // vC= -101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b1111111110110001; // vC=  -79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b1111111111010101; // vC=  -43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b1111111110010011; // vC= -109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b1111111110111110; // vC=  -66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011010; // iC=-1702 
vC = 14'b1111111110101101; // vC=  -83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b1111111111111111; // vC=   -1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b1111111110001001; // vC= -119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b1111111101111001; // vC= -135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110000; // iC=-1680 
vC = 14'b1111111110010000; // vC= -112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b1111111110110001; // vC=  -79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b1111111111100011; // vC=  -29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b1111111101001110; // vC= -178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b1111111110000001; // vC= -127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b1111111110001011; // vC= -117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b1111111110011101; // vC=  -99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b1111111110110000; // vC=  -80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b1111111111000001; // vC=  -63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111010; // iC=-1798 
vC = 14'b1111111100110101; // vC= -203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b1111111110001110; // vC= -114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b1111111101010010; // vC= -174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111111; // iC=-1665 
vC = 14'b1111111101010101; // vC= -171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b1111111101100110; // vC= -154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110011; // iC=-1741 
vC = 14'b1111111100101000; // vC= -216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b1111111100111001; // vC= -199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b1111111100001101; // vC= -243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b1111111011111010; // vC= -262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b1111111101001010; // vC= -182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b1111111100001000; // vC= -248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100100; // iC=-1692 
vC = 14'b1111111100111001; // vC= -199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b1111111101011011; // vC= -165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b1111111011000001; // vC= -319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b1111111100110110; // vC= -202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b1111111100100101; // vC= -219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b1111111100010010; // vC= -238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b1111111011001101; // vC= -307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b1111111101000010; // vC= -190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100101; // iC=-1627 
vC = 14'b1111111011010000; // vC= -304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b1111111011010110; // vC= -298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b1111111011110110; // vC= -266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b1111111100001000; // vC= -248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b1111111010000110; // vC= -378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b1111111011101001; // vC= -279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110111; // iC=-1609 
vC = 14'b1111111010000011; // vC= -381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b1111111010001110; // vC= -370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b1111111001110111; // vC= -393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b1111111001101110; // vC= -402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b1111111010011011; // vC= -357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b1111111011100000; // vC= -288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b1111111010001010; // vC= -374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b1111111010101000; // vC= -344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010011; // iC=-1581 
vC = 14'b1111111010010000; // vC= -368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001010; // iC=-1590 
vC = 14'b1111111010010101; // vC= -363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b1111111010111101; // vC= -323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001110; // iC=-1586 
vC = 14'b1111111001111110; // vC= -386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b1111111000101110; // vC= -466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b1111111000110011; // vC= -461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b1111111000011100; // vC= -484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b1111111000101101; // vC= -467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b1111111010010101; // vC= -363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011101; // iC=-1699 
vC = 14'b1111111001001000; // vC= -440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b1111111010001110; // vC= -370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100100; // iC=-1628 
vC = 14'b1111111000011110; // vC= -482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000101; // iC=-1595 
vC = 14'b1111111001011111; // vC= -417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b1111111001101001; // vC= -407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b1111111000001011; // vC= -501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b1111111001100100; // vC= -412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100101; // iC=-1691 
vC = 14'b1111110111010100; // vC= -556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b1111111000010111; // vC= -489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111100; // iC=-1668 
vC = 14'b1111111000101111; // vC= -465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110110; // iC=-1674 
vC = 14'b1111111000111100; // vC= -452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b1111111001010111; // vC= -425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010001; // iC=-1647 
vC = 14'b1111110111010100; // vC= -556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101100; // iC=-1556 
vC = 14'b1111110110101110; // vC= -594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b1111110111110110; // vC= -522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b1111110111000001; // vC= -575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b1111110110101100; // vC= -596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101001; // iC=-1623 
vC = 14'b1111111000011100; // vC= -484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010111; // iC=-1641 
vC = 14'b1111111000000000; // vC= -512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b1111111000001001; // vC= -503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b1111110111111001; // vC= -519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b1111111000001100; // vC= -500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b1111110101110000; // vC= -656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b1111110111000100; // vC= -572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b1111110101101010; // vC= -662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100100; // iC=-1564 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b1111110110000011; // vC= -637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101101; // iC=-1491 
vC = 14'b1111110110101011; // vC= -597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b1111110110010110; // vC= -618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b1111110110110000; // vC= -592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011011; // iC=-1573 
vC = 14'b1111110110011010; // vC= -614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010100; // iC=-1580 
vC = 14'b1111110110100000; // vC= -608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b1111110111001000; // vC= -568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b1111110100100101; // vC= -731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000100; // iC=-1468 
vC = 14'b1111110100110110; // vC= -714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b1111110110000000; // vC= -640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b1111110101101110; // vC= -658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100011; // iC=-1501 
vC = 14'b1111110100100100; // vC= -732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011101; // iC=-1443 
vC = 14'b1111110110010100; // vC= -620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001101; // iC=-1459 
vC = 14'b1111110100001011; // vC= -757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110010; // iC=-1486 
vC = 14'b1111110100100111; // vC= -729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101100; // iC=-1428 
vC = 14'b1111110100011011; // vC= -741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b1111110011110010; // vC= -782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010011; // iC=-1517 
vC = 14'b1111110101010100; // vC= -684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b1111110100000001; // vC= -767 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000100; // iC=-1468 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110110; // iC=-1418 
vC = 14'b1111110101100101; // vC= -667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001011; // iC=-1397 
vC = 14'b1111110100101100; // vC= -724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111001; // iC=-1415 
vC = 14'b1111110011110001; // vC= -783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100101; // iC=-1435 
vC = 14'b1111110011110001; // vC= -783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011101; // iC=-1379 
vC = 14'b1111110011001000; // vC= -824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000111; // iC=-1401 
vC = 14'b1111110011011100; // vC= -804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100011; // iC=-1501 
vC = 14'b1111110100111110; // vC= -706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011000; // iC=-1512 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001101; // iC=-1395 
vC = 14'b1111110101001011; // vC= -693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100101; // iC=-1371 
vC = 14'b1111110011100011; // vC= -797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010011; // iC=-1453 
vC = 14'b1111110100000000; // vC= -768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111111; // iC=-1473 
vC = 14'b1111110010100110; // vC= -858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b1111110011010111; // vC= -809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100110; // iC=-1434 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110000; // iC=-1488 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111111; // iC=-1345 
vC = 14'b1111110010101110; // vC= -850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b1111110100011101; // vC= -739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100110; // iC=-1370 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011000; // iC=-1320 
vC = 14'b1111110011010010; // vC= -814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100011; // iC=-1373 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b1111110010110101; // vC= -843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100000; // iC=-1376 
vC = 14'b1111110010110000; // vC= -848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100101; // iC=-1307 
vC = 14'b1111110001101000; // vC= -920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101010; // iC=-1430 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101001; // iC=-1431 
vC = 14'b1111110011001011; // vC= -821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b1111110010010000; // vC= -880 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011001; // iC=-1447 
vC = 14'b1111110010010000; // vC= -880 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000001; // iC=-1407 
vC = 14'b1111110011001001; // vC= -823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110111; // iC=-1353 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111010; // iC=-1286 
vC = 14'b1111110001110110; // vC= -906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111110010000000; // vC= -896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110001; // iC=-1359 
vC = 14'b1111110010100001; // vC= -863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011001; // iC=-1383 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101000; // iC=-1368 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000000; // iC=-1344 
vC = 14'b1111110001000010; // vC= -958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001111; // iC=-1265 
vC = 14'b1111110010110111; // vC= -841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011010; // iC=-1318 
vC = 14'b1111110001110010; // vC= -910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001000; // iC=-1272 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010011; // iC=-1325 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001111; // iC=-1329 
vC = 14'b1111110000110110; // vC= -970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010111; // iC=-1257 
vC = 14'b1111110000101110; // vC= -978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100000; // iC=-1248 
vC = 14'b1111110010100101; // vC= -859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101001; // iC=-1303 
vC = 14'b1111110001100011; // vC= -925 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111110; // iC=-1218 
vC = 14'b1111110010010111; // vC= -873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100100; // iC=-1244 
vC = 14'b1111110000110001; // vC= -975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101010; // iC=-1366 
vC = 14'b1111110001010101; // vC= -939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110100; // iC=-1292 
vC = 14'b1111110001110111; // vC= -905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001111; // iC=-1265 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111010; // iC=-1286 
vC = 14'b1111101111110100; // vC=-1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011101; // iC=-1315 
vC = 14'b1111110001101100; // vC= -916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100100; // iC=-1308 
vC = 14'b1111110001001111; // vC= -945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001101; // iC=-1331 
vC = 14'b1111101111100011; // vC=-1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000101; // iC=-1275 
vC = 14'b1111110000000111; // vC=-1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101101; // iC=-1235 
vC = 14'b1111110001001111; // vC= -945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010110; // iC=-1258 
vC = 14'b1111101111111001; // vC=-1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111010; // iC=-1222 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001111; // iC=-1265 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000001; // iC=-1215 
vC = 14'b1111101111110110; // vC=-1034 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b1111101111011001; // vC=-1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001110; // iC=-1202 
vC = 14'b1111110000110001; // vC= -975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101111; // iC=-1169 
vC = 14'b1111101111111100; // vC=-1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111110; // iC=-1282 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010011; // iC=-1261 
vC = 14'b1111101111010001; // vC=-1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110100; // iC=-1228 
vC = 14'b1111110000101111; // vC= -977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000110; // iC=-1210 
vC = 14'b1111101111001001; // vC=-1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011010; // iC=-1190 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100110; // iC=-1242 
vC = 14'b1111101110010100; // vC=-1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101010; // iC=-1174 
vC = 14'b1111110000010000; // vC=-1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000011; // iC=-1149 
vC = 14'b1111101110001110; // vC=-1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101111; // iC=-1169 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010001; // iC=-1199 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111001; // iC=-1159 
vC = 14'b1111101111100111; // vC=-1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000101; // iC=-1147 
vC = 14'b1111101111001101; // vC=-1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101001; // iC=-1175 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010101; // iC=-1195 
vC = 14'b1111101110111100; // vC=-1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010101; // iC=-1195 
vC = 14'b1111101111100100; // vC=-1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111101; // iC=-1219 
vC = 14'b1111101110010000; // vC=-1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001001; // iC=-1143 
vC = 14'b1111101111100010; // vC=-1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001101; // iC=-1075 
vC = 14'b1111101110001110; // vC=-1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110111; // iC=-1161 
vC = 14'b1111101111001110; // vC=-1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101011; // iC=-1045 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010010; // iC=-1134 
vC = 14'b1111101110000000; // vC=-1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010101; // iC=-1067 
vC = 14'b1111101110100111; // vC=-1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010011; // iC=-1069 
vC = 14'b1111101101111011; // vC=-1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010100; // iC=-1068 
vC = 14'b1111101110011001; // vC=-1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000001; // iC=-1023 
vC = 14'b1111101101110101; // vC=-1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001101; // iC=-1075 
vC = 14'b1111101110111100; // vC=-1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111101; // iC=-1091 
vC = 14'b1111101101101101; // vC=-1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101000; // iC=-1112 
vC = 14'b1111101101110111; // vC=-1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101101; // iC=-1043 
vC = 14'b1111101111000110; // vC=-1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011100; // iC=-1060 
vC = 14'b1111101101110011; // vC=-1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100110; // iC=-1050 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000101; // iC=-1083 
vC = 14'b1111101110011010; // vC=-1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111010; // iC=-1030 
vC = 14'b1111101100110010; // vC=-1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100011; // iC= -989 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011110; // iC=-1058 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011011; // iC= -997 
vC = 14'b1111101101010011; // vC=-1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110100; // iC=-1100 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111101; // iC= -963 
vC = 14'b1111101101100110; // vC=-1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000011; // iC=-1085 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101111; // iC=-1041 
vC = 14'b1111101110010001; // vC=-1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101100; // iC=-1044 
vC = 14'b1111101101100110; // vC=-1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100101; // iC=-1051 
vC = 14'b1111101101110111; // vC=-1161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011011; // iC= -933 
vC = 14'b1111101101111100; // vC=-1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111010; // iC= -966 
vC = 14'b1111101101010001; // vC=-1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001011; // iC=-1077 
vC = 14'b1111101110001100; // vC=-1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110000; // iC=-1040 
vC = 14'b1111101100110100; // vC=-1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010000; // iC= -944 
vC = 14'b1111101100100000; // vC=-1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000010; // iC= -958 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111110; // iC=-1026 
vC = 14'b1111101100010011; // vC=-1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001010; // iC=-1014 
vC = 14'b1111101100111010; // vC=-1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011001; // iC= -999 
vC = 14'b1111101011011111; // vC=-1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b1111101100101011; // vC=-1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000000; // iC=-1024 
vC = 14'b1111101101110110; // vC=-1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101111; // iC= -977 
vC = 14'b1111101101000001; // vC=-1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010011; // iC=-1005 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001001; // iC=-1015 
vC = 14'b1111101101100111; // vC=-1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010101; // iC= -939 
vC = 14'b1111101011100110; // vC=-1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011010; // iC= -998 
vC = 14'b1111101100011101; // vC=-1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011111; // iC= -993 
vC = 14'b1111101101000110; // vC=-1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000110; // iC= -890 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100010; // iC= -862 
vC = 14'b1111101100111110; // vC=-1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001110; // iC= -946 
vC = 14'b1111101011000001; // vC=-1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101111; // iC= -849 
vC = 14'b1111101101001010; // vC=-1206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111110; // iC= -962 
vC = 14'b1111101100100000; // vC=-1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011010; // iC= -934 
vC = 14'b1111101100011011; // vC=-1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011000; // iC= -872 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000100; // iC= -828 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011110; // iC= -802 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110111; // iC= -905 
vC = 14'b1111101010111101; // vC=-1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101001; // iC= -791 
vC = 14'b1111101100100101; // vC=-1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110101; // iC= -843 
vC = 14'b1111101100111100; // vC=-1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100000; // iC= -800 
vC = 14'b1111101011110001; // vC=-1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110111; // iC= -841 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111010; // iC= -774 
vC = 14'b1111101010111100; // vC=-1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110101; // iC= -907 
vC = 14'b1111101010110101; // vC=-1355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001011; // iC= -885 
vC = 14'b1111101100101111; // vC=-1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101101; // iC= -851 
vC = 14'b1111101011111010; // vC=-1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110101; // iC= -843 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110101; // iC= -843 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010110; // iC= -810 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110111; // iC= -777 
vC = 14'b1111101011011110; // vC=-1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000001; // iC= -767 
vC = 14'b1111101100010111; // vC=-1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010101; // iC= -747 
vC = 14'b1111101011101001; // vC=-1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010100; // iC= -748 
vC = 14'b1111101100001000; // vC=-1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111010; // iC= -838 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111001; // iC= -839 
vC = 14'b1111101011101101; // vC=-1299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101001; // iC= -855 
vC = 14'b1111101011001110; // vC=-1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010001; // iC= -751 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100100; // iC= -796 
vC = 14'b1111101010100001; // vC=-1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000011; // iC= -701 
vC = 14'b1111101100000100; // vC=-1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000011; // iC= -829 
vC = 14'b1111101010001110; // vC=-1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000100; // iC= -764 
vC = 14'b1111101011111000; // vC=-1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100011; // iC= -733 
vC = 14'b1111101011110110; // vC=-1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100101; // iC= -731 
vC = 14'b1111101011010011; // vC=-1325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100011; // iC= -797 
vC = 14'b1111101001100100; // vC=-1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001011; // iC= -757 
vC = 14'b1111101010101111; // vC=-1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011100; // iC= -676 
vC = 14'b1111101011001101; // vC=-1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111001; // iC= -647 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011100; // iC= -676 
vC = 14'b1111101001110010; // vC=-1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111110; // iC= -706 
vC = 14'b1111101011010001; // vC=-1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111000; // iC= -648 
vC = 14'b1111101001100101; // vC=-1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000101; // iC= -699 
vC = 14'b1111101001111101; // vC=-1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110100; // iC= -652 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101111; // iC= -657 
vC = 14'b1111101010100010; // vC=-1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001011; // iC= -757 
vC = 14'b1111101011001010; // vC=-1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010101; // iC= -683 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100010; // iC= -606 
vC = 14'b1111101001110101; // vC=-1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110101; // iC= -715 
vC = 14'b1111101001101000; // vC=-1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101110; // iC= -594 
vC = 14'b1111101011011001; // vC=-1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111101001011000; // vC=-1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101001; // iC= -663 
vC = 14'b1111101010111010; // vC=-1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111101; // iC= -579 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011000; // iC= -616 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000100; // iC= -700 
vC = 14'b1111101001110001; // vC=-1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110011; // iC= -653 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001110; // iC= -626 
vC = 14'b1111101000100111; // vC=-1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010100; // iC= -556 
vC = 14'b1111101010001110; // vC=-1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100101; // iC= -667 
vC = 14'b1111101010011011; // vC=-1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111110; // iC= -578 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b1111101010011010; // vC=-1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110001; // iC= -655 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110110; // iC= -650 
vC = 14'b1111101001110100; // vC=-1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111010; // iC= -518 
vC = 14'b1111101010110111; // vC=-1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001110; // iC= -626 
vC = 14'b1111101000111111; // vC=-1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000100; // iC= -636 
vC = 14'b1111101010110100; // vC=-1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011011; // iC= -485 
vC = 14'b1111101001001110; // vC=-1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100001; // iC= -479 
vC = 14'b1111101000011111; // vC=-1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100011; // iC= -477 
vC = 14'b1111101000100000; // vC=-1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111000; // iC= -520 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011111; // iC= -481 
vC = 14'b1111101001111101; // vC=-1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000110; // iC= -506 
vC = 14'b1111101000100001; // vC=-1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101000; // iC= -472 
vC = 14'b1111101010000011; // vC=-1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100001; // iC= -543 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001001; // iC= -567 
vC = 14'b1111101000111110; // vC=-1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011001; // iC= -423 
vC = 14'b1111101001100110; // vC=-1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001000; // iC= -440 
vC = 14'b1111101001011010; // vC=-1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101110; // iC= -530 
vC = 14'b1111101001110010; // vC=-1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101001; // iC= -535 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100100; // iC= -540 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110110; // iC= -458 
vC = 14'b1111101000011110; // vC=-1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101000; // iC= -536 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000111; // iC= -377 
vC = 14'b1111101000101111; // vC=-1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110111; // iC= -457 
vC = 14'b1111101000100101; // vC=-1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110011; // iC= -525 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001011; // iC= -437 
vC = 14'b1111101000100110; // vC=-1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100101; // iC= -475 
vC = 14'b1111101000110100; // vC=-1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010011; // iC= -429 
vC = 14'b1111101000001111; // vC=-1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010001; // iC= -431 
vC = 14'b1111101000111100; // vC=-1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000011; // iC= -381 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010100; // iC= -364 
vC = 14'b1111101000001000; // vC=-1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011001; // iC= -423 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000110; // iC= -378 
vC = 14'b1111101000100000; // vC=-1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100001; // iC= -351 
vC = 14'b1111101000110110; // vC=-1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001001; // iC= -311 
vC = 14'b1111100111101010; // vC=-1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011010; // iC= -294 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010110; // iC= -298 
vC = 14'b1111100111110101; // vC=-1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100000; // iC= -288 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111011; // iC= -261 
vC = 14'b1111101000000100; // vC=-1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111000; // iC= -200 
vC = 14'b1111101001011111; // vC=-1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000101; // iC= -187 
vC = 14'b1111101001110110; // vC=-1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001001; // iC= -311 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101000; // iC= -152 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010010; // iC= -174 
vC = 14'b1111100111100100; // vC=-1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100110; // iC= -154 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001101; // iC= -179 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111101; // iC= -131 
vC = 14'b1111101000001000; // vC=-1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010110; // iC= -106 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010011; // iC= -173 
vC = 14'b1111101001100110; // vC=-1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111011; // iC= -197 
vC = 14'b1111100111101011; // vC=-1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000101; // iC= -123 
vC = 14'b1111101001011000; // vC=-1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110011; // iC= -141 
vC = 14'b1111101001101001; // vC=-1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100010; // iC=  -30 
vC = 14'b1111101001001000; // vC=-1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000110; // iC=    6 
vC = 14'b1111101000100110; // vC=-1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000010; // iC=    2 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100001; // iC=  -95 
vC = 14'b1111101000000001; // vC=-1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100110; // iC=  -26 
vC = 14'b1111100111101001; // vC=-1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001000; // iC=  -56 
vC = 14'b1111101000011001; // vC=-1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011101; // iC=   29 
vC = 14'b1111101001101010; // vC=-1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110101; // iC=   53 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011111; // iC=   95 
vC = 14'b1111100111100111; // vC=-1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010001; // iC=   81 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011011; // iC=   27 
vC = 14'b1111100111011001; // vC=-1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000010; // iC=  194 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000011; // iC=  131 
vC = 14'b1111100111101111; // vC=-1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100100; // iC=  100 
vC = 14'b1111101001000011; // vC=-1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011011; // iC=  219 
vC = 14'b1111100111111001; // vC=-1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100011; // iC=  163 
vC = 14'b1111101001000000; // vC=-1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001100; // iC=  204 
vC = 14'b1111101000100011; // vC=-1501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101000; // iC=  296 
vC = 14'b1111101000010110; // vC=-1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101000; // iC=  232 
vC = 14'b1111101001110010; // vC=-1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000100; // iC=  260 
vC = 14'b1111100111110011; // vC=-1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101000; // iC=  360 
vC = 14'b1111101000100010; // vC=-1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010100; // iC=  276 
vC = 14'b1111101000111011; // vC=-1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110111; // iC=  311 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000011; // iC=  451 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110111; // iC=  439 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000101; // iC=  389 
vC = 14'b1111101000010111; // vC=-1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010010; // iC=  530 
vC = 14'b1111101010001010; // vC=-1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100000; // iC=  480 
vC = 14'b1111101000011101; // vC=-1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010110; // iC=  470 
vC = 14'b1111100111111000; // vC=-1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000000; // iC=  576 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110011; // iC=  627 
vC = 14'b1111101000100011; // vC=-1501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000011; // iC=  515 
vC = 14'b1111101000000111; // vC=-1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101100; // iC=  620 
vC = 14'b1111101001101010; // vC=-1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101101; // iC=  685 
vC = 14'b1111101000001101; // vC=-1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111011; // iC=  635 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000000; // iC=  640 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010001; // iC=  721 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001010; // iC=  778 
vC = 14'b1111101001111110; // vC=-1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110101; // iC=  693 
vC = 14'b1111101000000100; // vC=-1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110000; // iC=  688 
vC = 14'b1111101000111111; // vC=-1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011110; // iC=  862 
vC = 14'b1111101001110110; // vC=-1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010101; // iC=  789 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001011; // iC=  907 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000111; // iC=  839 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110100; // iC=  948 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111011; // iC=  827 
vC = 14'b1111101000111001; // vC=-1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010001; // iC=  849 
vC = 14'b1111101001110001; // vC=-1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011000; // iC=  984 
vC = 14'b1111101000100110; // vC=-1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001101; // iC=  909 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011000; // iC= 1048 
vC = 14'b1111101010101110; // vC=-1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011111; // iC= 1055 
vC = 14'b1111101010101111; // vC=-1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000011; // iC= 1091 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011010; // iC=  986 
vC = 14'b1111101011000010; // vC=-1342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000001; // iC= 1025 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001001; // iC= 1161 
vC = 14'b1111101001010001; // vC=-1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111110; // iC= 1086 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110000; // iC= 1072 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001100; // iC= 1164 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010101; // iC= 1173 
vC = 14'b1111101001100110; // vC=-1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100000; // iC= 1184 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011100; // iC= 1244 
vC = 14'b1111101010111010; // vC=-1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110110; // iC= 1270 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111110; // iC= 1214 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001101; // iC= 1293 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111110; // iC= 1278 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100000; // iC= 1312 
vC = 14'b1111101011101100; // vC=-1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100011; // iC= 1379 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101001; // iC= 1385 
vC = 14'b1111101010110001; // vC=-1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010110; // iC= 1302 
vC = 14'b1111101011110100; // vC=-1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001000; // iC= 1416 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000000; // iC= 1344 
vC = 14'b1111101010111101; // vC=-1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111010; // iC= 1466 
vC = 14'b1111101011001000; // vC=-1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000011; // iC= 1475 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100100; // iC= 1508 
vC = 14'b1111101010010110; // vC=-1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110111; // iC= 1399 
vC = 14'b1111101100010001; // vC=-1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011101; // iC= 1437 
vC = 14'b1111101011010000; // vC=-1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000011; // iC= 1475 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101000; // iC= 1448 
vC = 14'b1111101011001010; // vC=-1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100001; // iC= 1441 
vC = 14'b1111101011011001; // vC=-1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001010; // iC= 1546 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001110; // iC= 1550 
vC = 14'b1111101100011110; // vC=-1250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010111; // iC= 1623 
vC = 14'b1111101011010111; // vC=-1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100000; // iC= 1504 
vC = 14'b1111101011101000; // vC=-1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110101; // iC= 1589 
vC = 14'b1111101100110011; // vC=-1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000101; // iC= 1669 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000111; // iC= 1671 
vC = 14'b1111101100111100; // vC=-1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111100; // iC= 1596 
vC = 14'b1111101100100110; // vC=-1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011011; // iC= 1563 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100001; // iC= 1633 
vC = 14'b1111101100011011; // vC=-1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011111; // iC= 1631 
vC = 14'b1111101011110010; // vC=-1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001111; // iC= 1679 
vC = 14'b1111101011111001; // vC=-1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011000; // iC= 1624 
vC = 14'b1111101101100011; // vC=-1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000101; // iC= 1669 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100001; // iC= 1633 
vC = 14'b1111101100100110; // vC=-1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b1111101100011011; // vC=-1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111110; // iC= 1662 
vC = 14'b1111101110000001; // vC=-1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110001; // iC= 1777 
vC = 14'b1111101100111000; // vC=-1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b1111101101000000; // vC=-1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b1111101101100000; // vC=-1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101111; // iC= 1711 
vC = 14'b1111101110000110; // vC=-1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b1111101110010001; // vC=-1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b1111101101111010; // vC=-1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101001; // iC= 1833 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b1111101111100100; // vC=-1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111111; // iC= 1791 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b1111101110010100; // vC=-1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111001; // iC= 1785 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100011; // iC= 1827 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100100; // iC= 1764 
vC = 14'b1111101111001100; // vC=-1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011000; // iC= 1880 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111101111111000; // vC=-1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b1111101111110100; // vC=-1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111101111100100; // vC=-1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b1111110000010101; // vC=-1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110100; // iC= 1780 
vC = 14'b1111101111101000; // vC=-1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111101111011101; // vC=-1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101011; // iC= 1835 
vC = 14'b1111110000101001; // vC= -983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111101111011010; // vC=-1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111101110111001; // vC=-1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111101110111100; // vC=-1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111110000010001; // vC=-1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111101111111011; // vC=-1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b1111110001000111; // vC= -953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111110001010010; // vC= -942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b1111110000110010; // vC= -974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111110001111100; // vC= -900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110001; // iC= 1841 
vC = 14'b1111110001000010; // vC= -958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110000; // iC= 1840 
vC = 14'b1111110000011111; // vC= -993 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110001001000; // vC= -952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000010; // iC= 1858 
vC = 14'b1111110010110011; // vC= -845 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b1111110000101101; // vC= -979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001010; // iC= 1994 
vC = 14'b1111110010100101; // vC= -859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111110001111110; // vC= -898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110011001000; // vC= -824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111110011001011; // vC= -821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111110011011001; // vC= -807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000101; // iC= 1861 
vC = 14'b1111110001101110; // vC= -914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b1111110010111000; // vC= -840 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111110001111100; // vC= -900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b1111110100011101; // vC= -739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b1111110011100110; // vC= -794 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111110010011101; // vC= -867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b1111110101000000; // vC= -704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100001; // iC= 2017 
vC = 14'b1111110010111110; // vC= -834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111110011011111; // vC= -801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b1111110100100111; // vC= -729 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111110011001111; // vC= -817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111110100000010; // vC= -766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111110100101111; // vC= -721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111110101101111; // vC= -657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111110100101000; // vC= -728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b1111110101111100; // vC= -644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111110100001011; // vC= -757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b1111110110001100; // vC= -628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b1111110100100100; // vC= -732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b1111110110100010; // vC= -606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000000; // iC= 1984 
vC = 14'b1111110110101000; // vC= -600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b1111110101001000; // vC= -696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b1111110100111110; // vC= -706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111110110111011; // vC= -581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111110101000001; // vC= -703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111110101001001; // vC= -695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b1111110101001111; // vC= -689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111110101111101; // vC= -643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111110110001000; // vC= -632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111110110100100; // vC= -604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111110101110010; // vC= -654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111110110110110; // vC= -586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111100; // iC= 2044 
vC = 14'b1111110110001011; // vC= -629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111110111100110; // vC= -538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110110110110; // vC= -586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000100; // iC= 2052 
vC = 14'b1111110111100001; // vC= -543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111110111011111; // vC= -545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100011; // iC= 2019 
vC = 14'b1111111000100011; // vC= -477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111110110100100; // vC= -604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001010; // iC= 2058 
vC = 14'b1111111000111010; // vC= -454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010001; // iC= 2065 
vC = 14'b1111111000000011; // vC= -509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101110; // iC= 2030 
vC = 14'b1111110111100001; // vC= -543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111000010101; // vC= -491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b1111111000000000; // vC= -512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110100; // iC= 1972 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b1111111001001001; // vC= -439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111111001011100; // vC= -420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101110; // iC= 2030 
vC = 14'b1111111000001001; // vC= -503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111111000101100; // vC= -468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b1111111010000010; // vC= -382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b1111111000010110; // vC= -490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000100; // iC= 1924 
vC = 14'b1111111001111011; // vC= -389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111111001101000; // vC= -408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b1111111010010011; // vC= -365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111111001110000; // vC= -400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111111000011010; // vC= -486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011000; // iC= 2072 
vC = 14'b1111111001001101; // vC= -435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111111000110100; // vC= -460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111111010100100; // vC= -348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b1111111010010100; // vC= -364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011100; // iC= 2076 
vC = 14'b1111111010001011; // vC= -373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111111001111000; // vC= -392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111011100100; // vC= -284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b1111111001010001; // vC= -431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111111; // iC= 2047 
vC = 14'b1111111010101011; // vC= -341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111111011001011; // vC= -309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b1111111100000010; // vC= -254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111111011100101; // vC= -283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001011; // iC= 2059 
vC = 14'b1111111011000011; // vC= -317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111111011010101; // vC= -299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000111; // iC= 1991 
vC = 14'b1111111010000101; // vC= -379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011010; // iC= 2074 
vC = 14'b1111111100010110; // vC= -234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111011010101; // vC= -299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111111100101010; // vC= -214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111111011000001; // vC= -319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011111; // iC= 2079 
vC = 14'b1111111010100010; // vC= -350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000111; // iC= 2055 
vC = 14'b1111111011010011; // vC= -301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000010; // iC= 2050 
vC = 14'b1111111100100011; // vC= -221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111011000111; // vC= -313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101011; // iC= 2027 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010100; // iC= 2068 
vC = 14'b1111111011101001; // vC= -279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111111011111010; // vC= -262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b1111111100111101; // vC= -195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010110; // iC= 2070 
vC = 14'b1111111110000011; // vC= -125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111111101111010; // vC= -134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111111100010001; // vC= -239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b1111111100011101; // vC= -227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b1111111100001001; // vC= -247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111111101011011; // vC= -165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b1111111110100000; // vC=  -96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111111101011100; // vC= -164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101011; // iC= 2027 
vC = 14'b1111111111001001; // vC=  -55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000011; // iC= 2051 
vC = 14'b1111111101101111; // vC= -145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111111110101111; // vC=  -81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111100; // iC= 2044 
vC = 14'b1111111101100110; // vC= -154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111000; // iC= 2040 
vC = 14'b1111111110100101; // vC=  -91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111111111011101; // vC=  -35 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111111101100110; // vC= -154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111101111110; // vC= -130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b0000000000000001; // vC=    1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b1111111110110000; // vC=  -80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b0000000000001111; // vC=   15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b1111111110110100; // vC=  -76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b1111111111011111; // vC=  -33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111111110001111; // vC= -113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001001; // iC= 2057 
vC = 14'b1111111110011001; // vC= -103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111111111101000; // vC=  -24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111111110110100; // vC=  -76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111111110101111; // vC=  -81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b0000000000010110; // vC=   22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b0000000000110001; // vC=   49 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111111111010011; // vC=  -45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b0000000001101100; // vC=  108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b0000000001011010; // vC=   90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b0000000000101110; // vC=   46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b0000000010000101; // vC=  133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011001; // iC= 1881 
vC = 14'b0000000000100110; // vC=   38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b0000000001010011; // vC=   83 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b0000000001010000; // vC=   80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b0000000001011001; // vC=   89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011110; // iC= 1886 
vC = 14'b0000000001110010; // vC=  114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b0000000000111100; // vC=   60 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b0000000010101111; // vC=  175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b0000000011001100; // vC=  204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b0000000011011100; // vC=  220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b0000000010110000; // vC=  176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000100; // iC= 1860 
vC = 14'b0000000011110010; // vC=  242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000000011000111; // vC=  199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110111; // iC= 1975 
vC = 14'b0000000011001010; // vC=  202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b0000000010101101; // vC=  173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000011001111; // vC=  207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b0000000100010001; // vC=  273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b0000000010111100; // vC=  188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b0000000010110110; // vC=  182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b0000000011110001; // vC=  241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001101; // iC= 1869 
vC = 14'b0000000100101100; // vC=  300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b0000000011001000; // vC=  200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000101; // iC= 1861 
vC = 14'b0000000011101111; // vC=  239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b0000000101100100; // vC=  356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b0000000101100001; // vC=  353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000111; // iC= 1863 
vC = 14'b0000000101010010; // vC=  338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b0000000101100000; // vC=  352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b0000000101101011; // vC=  363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101001; // iC= 1833 
vC = 14'b0000000100111000; // vC=  312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b0000000100100101; // vC=  293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101001; // iC= 1833 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b0000000110010111; // vC=  407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b0000000101101101; // vC=  365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b0000000110100001; // vC=  417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b0000000110101100; // vC=  428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b0000000100111111; // vC=  319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b0000000100100110; // vC=  294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111001; // iC= 1913 
vC = 14'b0000000100111111; // vC=  319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b0000000100110010; // vC=  306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b0000000100111101; // vC=  317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b0000000101011110; // vC=  350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b0000000111000100; // vC=  452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b0000000111001100; // vC=  460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100011; // iC= 1827 
vC = 14'b0000000110110111; // vC=  439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b0000000101101011; // vC=  363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011110; // iC= 1886 
vC = 14'b0000000101101101; // vC=  365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100000; // iC= 1824 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111100; // iC= 1788 
vC = 14'b0000000111001100; // vC=  460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010100; // iC= 1876 
vC = 14'b0000000111110101; // vC=  501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b0000000101111000; // vC=  376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111011; // iC= 1851 
vC = 14'b0000000110100001; // vC=  417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001100; // iC= 1804 
vC = 14'b0000000111111001; // vC=  505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011100; // iC= 1820 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b0000000110100001; // vC=  417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b0000000111100001; // vC=  481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110010; // iC= 1778 
vC = 14'b0000000111010110; // vC=  470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010000; // iC= 1808 
vC = 14'b0000001000011000; // vC=  536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b0000001000110111; // vC=  567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b0000000111001101; // vC=  461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000000111110011; // vC=  499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b0000001001010101; // vC=  597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100010; // iC= 1826 
vC = 14'b0000001000000000; // vC=  512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000110; // iC= 1798 
vC = 14'b0000001000101001; // vC=  553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b0000001000000110; // vC=  518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b0000000111100111; // vC=  487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111000; // iC= 1784 
vC = 14'b0000001001011010; // vC=  602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011100; // iC= 1884 
vC = 14'b0000001000010100; // vC=  532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b0000001010000001; // vC=  641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010010; // iC= 1874 
vC = 14'b0000001001001000; // vC=  584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010001; // iC= 1873 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b0000001000001101; // vC=  525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b0000001010000000; // vC=  640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001000; // iC= 1864 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b0000001001100011; // vC=  611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b0000001000101110; // vC=  558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b0000001011000000; // vC=  704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b0000001001010000; // vC=  592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001001; // iC= 1737 
vC = 14'b0000001010100111; // vC=  679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100011; // iC= 1699 
vC = 14'b0000001001011101; // vC=  605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b0000001001000110; // vC=  582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101001; // iC= 1705 
vC = 14'b0000001001011100; // vC=  604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010110; // iC= 1686 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000100; // iC= 1668 
vC = 14'b0000001011101000; // vC=  744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000111; // iC= 1799 
vC = 14'b0000001010101011; // vC=  683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000001010010001; // vC=  657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b0000001011111001; // vC=  761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111000; // iC= 1720 
vC = 14'b0000001010100100; // vC=  676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b0000001010101110; // vC=  686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100110; // iC= 1702 
vC = 14'b0000001010110011; // vC=  691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b0000001010110101; // vC=  693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b0000001010101100; // vC=  684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b0000001100110001; // vC=  817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000110; // iC= 1670 
vC = 14'b0000001011001010; // vC=  714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b0000001010101000; // vC=  680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111010; // iC= 1658 
vC = 14'b0000001010110110; // vC=  694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011000; // iC= 1752 
vC = 14'b0000001101001011; // vC=  843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010100; // iC= 1620 
vC = 14'b0000001100001111; // vC=  783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010010; // iC= 1618 
vC = 14'b0000001101001010; // vC=  842 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001000; // iC= 1672 
vC = 14'b0000001011111001; // vC=  761 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011000; // iC= 1624 
vC = 14'b0000001011110100; // vC=  756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110001; // iC= 1649 
vC = 14'b0000001100110001; // vC=  817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110110; // iC= 1654 
vC = 14'b0000001101010001; // vC=  849 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110000; // iC= 1648 
vC = 14'b0000001011111111; // vC=  767 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b0000001100010111; // vC=  791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b0000001101010111; // vC=  855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110100; // iC= 1588 
vC = 14'b0000001011111100; // vC=  764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101001; // iC= 1705 
vC = 14'b0000001101010101; // vC=  853 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000001; // iC= 1729 
vC = 14'b0000001101011010; // vC=  858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b0000001100010000; // vC=  784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110110; // iC= 1590 
vC = 14'b0000001100100011; // vC=  803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001110; // iC= 1614 
vC = 14'b0000001101110001; // vC=  881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000001100110000; // vC=  816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100100; // iC= 1572 
vC = 14'b0000001110100100; // vC=  932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011010; // iC= 1562 
vC = 14'b0000001110010001; // vC=  913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b0000001101110010; // vC=  882 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100000; // iC= 1632 
vC = 14'b0000001110110101; // vC=  949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111100; // iC= 1596 
vC = 14'b0000001110010001; // vC=  913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111101; // iC= 1597 
vC = 14'b0000001110000101; // vC=  901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001111; // iC= 1615 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101011; // iC= 1579 
vC = 14'b0000001111010100; // vC=  980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110011; // iC= 1523 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100110; // iC= 1574 
vC = 14'b0000001110010101; // vC=  917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001000; // iC= 1544 
vC = 14'b0000001110001011; // vC=  907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101001; // iC= 1641 
vC = 14'b0000001111100101; // vC=  997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010111; // iC= 1623 
vC = 14'b0000001110001111; // vC=  911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001110010000; // vC=  912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011001; // iC= 1561 
vC = 14'b0000001110011011; // vC=  923 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111101; // iC= 1597 
vC = 14'b0000001111010000; // vC=  976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000010; // iC= 1538 
vC = 14'b0000001111101011; // vC= 1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011100; // iC= 1564 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101010; // iC= 1642 
vC = 14'b0000001110011001; // vC=  921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000000; // iC= 1600 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b0000001110101011; // vC=  939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b0000001110001111; // vC=  911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010010; // iC= 1490 
vC = 14'b0000001111011111; // vC=  991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010000; // iC= 1552 
vC = 14'b0000001110011100; // vC=  924 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011100; // iC= 1500 
vC = 14'b0000010000101011; // vC= 1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111101; // iC= 1597 
vC = 14'b0000001111010110; // vC=  982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100010; // iC= 1506 
vC = 14'b0000010000011100; // vC= 1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110000; // iC= 1456 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111101; // iC= 1597 
vC = 14'b0000001110101101; // vC=  941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001111; // iC= 1487 
vC = 14'b0000010000000011; // vC= 1027 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101110; // iC= 1582 
vC = 14'b0000001111110010; // vC= 1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100000; // iC= 1504 
vC = 14'b0000010000000010; // vC= 1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001111; // iC= 1423 
vC = 14'b0000001111100011; // vC=  995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111110; // iC= 1534 
vC = 14'b0000001111100011; // vC=  995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001010; // iC= 1482 
vC = 14'b0000010001000010; // vC= 1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b0000010000000111; // vC= 1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100111; // iC= 1447 
vC = 14'b0000010000000101; // vC= 1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000011; // iC= 1475 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000010; // iC= 1538 
vC = 14'b0000010001000010; // vC= 1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100100; // iC= 1444 
vC = 14'b0000010001001110; // vC= 1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011000; // iC= 1432 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b0000010010000100; // vC= 1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100001; // iC= 1377 
vC = 14'b0000010001011100; // vC= 1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111011; // iC= 1531 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111100; // iC= 1404 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100000; // iC= 1376 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110010; // iC= 1394 
vC = 14'b0000010001111000; // vC= 1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000110; // iC= 1414 
vC = 14'b0000010000000100; // vC= 1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010001; // iC= 1489 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101011; // iC= 1451 
vC = 14'b0000010010011110; // vC= 1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111000; // iC= 1464 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100001; // iC= 1377 
vC = 14'b0000010010000001; // vC= 1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100111; // iC= 1447 
vC = 14'b0000010001100001; // vC= 1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110110; // iC= 1334 
vC = 14'b0000010001111011; // vC= 1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111100; // iC= 1404 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011100; // iC= 1436 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001110; // iC= 1358 
vC = 14'b0000010010111101; // vC= 1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100110; // iC= 1318 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110011; // iC= 1331 
vC = 14'b0000010010011001; // vC= 1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100111; // iC= 1447 
vC = 14'b0000010010001011; // vC= 1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010000; // iC= 1424 
vC = 14'b0000010001101000; // vC= 1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110100; // iC= 1332 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001111; // iC= 1295 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001011; // iC= 1355 
vC = 14'b0000010001111000; // vC= 1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010110; // iC= 1430 
vC = 14'b0000010010001101; // vC= 1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101011; // iC= 1387 
vC = 14'b0000010001010110; // vC= 1110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100111; // iC= 1319 
vC = 14'b0000010011001101; // vC= 1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011001; // iC= 1369 
vC = 14'b0000010011110011; // vC= 1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011001; // iC= 1305 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001001; // iC= 1353 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110000; // iC= 1328 
vC = 14'b0000010010001111; // vC= 1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111110; // iC= 1342 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110100; // iC= 1396 
vC = 14'b0000010011001110; // vC= 1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000100; // iC= 1348 
vC = 14'b0000010010011110; // vC= 1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001101; // iC= 1357 
vC = 14'b0000010010100000; // vC= 1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100001; // iC= 1313 
vC = 14'b0000010010101111; // vC= 1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100001; // iC= 1377 
vC = 14'b0000010100011010; // vC= 1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100000; // iC= 1376 
vC = 14'b0000010100000001; // vC= 1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101100; // iC= 1260 
vC = 14'b0000010011111010; // vC= 1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011101; // iC= 1309 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110101; // iC= 1205 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111110; // iC= 1214 
vC = 14'b0000010100100101; // vC= 1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001001; // iC= 1353 
vC = 14'b0000010011111000; // vC= 1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101000; // iC= 1320 
vC = 14'b0000010100000011; // vC= 1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000001; // iC= 1217 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000111; // iC= 1287 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110111; // iC= 1335 
vC = 14'b0000010011111100; // vC= 1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101101; // iC= 1197 
vC = 14'b0000010100100101; // vC= 1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000010100001000; // vC= 1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010010; // iC= 1170 
vC = 14'b0000010011011010; // vC= 1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011101; // iC= 1309 
vC = 14'b0000010101010001; // vC= 1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010000; // iC= 1296 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010011; // iC= 1235 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101111; // iC= 1199 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001011; // iC= 1163 
vC = 14'b0000010011110111; // vC= 1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001100; // iC= 1164 
vC = 14'b0000010011111000; // vC= 1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000001; // iC= 1153 
vC = 14'b0000010101010011; // vC= 1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011010; // iC= 1178 
vC = 14'b0000010011111010; // vC= 1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001100; // iC= 1164 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101110; // iC= 1262 
vC = 14'b0000010011100010; // vC= 1250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101111; // iC= 1135 
vC = 14'b0000010100001110; // vC= 1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011000; // iC= 1176 
vC = 14'b0000010100101011; // vC= 1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010111; // iC= 1111 
vC = 14'b0000010101001001; // vC= 1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000101; // iC= 1221 
vC = 14'b0000010100101010; // vC= 1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000100; // iC= 1156 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000000; // iC= 1152 
vC = 14'b0000010100001000; // vC= 1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100101; // iC= 1189 
vC = 14'b0000010101010011; // vC= 1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111111; // iC= 1215 
vC = 14'b0000010011111110; // vC= 1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111011; // iC= 1147 
vC = 14'b0000010100110100; // vC= 1332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011010; // iC= 1114 
vC = 14'b0000010110000101; // vC= 1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101100; // iC= 1068 
vC = 14'b0000010101001111; // vC= 1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000010110011001; // vC= 1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010111; // iC= 1047 
vC = 14'b0000010101101011; // vC= 1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001111; // iC= 1103 
vC = 14'b0000010101010100; // vC= 1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100101; // iC= 1125 
vC = 14'b0000010110101000; // vC= 1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010101; // iC= 1045 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000100; // iC= 1028 
vC = 14'b0000010100011100; // vC= 1308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000010101100111; // vC= 1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111100; // iC= 1148 
vC = 14'b0000010110010011; // vC= 1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110010; // iC= 1074 
vC = 14'b0000010100110010; // vC= 1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001111; // iC= 1039 
vC = 14'b0000010101111110; // vC= 1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011011; // iC= 1115 
vC = 14'b0000010100110111; // vC= 1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011100; // iC= 1116 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011101; // iC=  989 
vC = 14'b0000010101110001; // vC= 1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110100; // iC= 1140 
vC = 14'b0000010100101100; // vC= 1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000010; // iC= 1090 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010001; // iC= 1041 
vC = 14'b0000010111000011; // vC= 1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100001; // iC= 1121 
vC = 14'b0000010101000011; // vC= 1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100110; // iC=  998 
vC = 14'b0000010101101101; // vC= 1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111110; // iC= 1022 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001110; // iC=  974 
vC = 14'b0000010101111001; // vC= 1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000110; // iC= 1030 
vC = 14'b0000010111010010; // vC= 1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111000; // iC=  952 
vC = 14'b0000010101000111; // vC= 1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001110; // iC=  974 
vC = 14'b0000010101101001; // vC= 1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010111; // iC=  983 
vC = 14'b0000010110011011; // vC= 1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001111; // iC=  975 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011111; // iC=  991 
vC = 14'b0000010101110001; // vC= 1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110110; // iC= 1014 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001010; // iC=  906 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101101; // iC= 1005 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000010; // iC= 1026 
vC = 14'b0000010110100000; // vC= 1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100100; // iC=  996 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011001; // iC=  921 
vC = 14'b0000010110111110; // vC= 1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110000; // iC= 1008 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110101; // iC= 1013 
vC = 14'b0000010111100001; // vC= 1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111111; // iC=  895 
vC = 14'b0000010111110011; // vC= 1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010100; // iC=  980 
vC = 14'b0000010110001011; // vC= 1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111001; // iC=  889 
vC = 14'b0000010111011011; // vC= 1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100110; // iC=  998 
vC = 14'b0000010111010101; // vC= 1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001110; // iC=  846 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111000; // iC=  952 
vC = 14'b0000010111000000; // vC= 1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111110; // iC=  894 
vC = 14'b0000010111111001; // vC= 1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000101; // iC=  837 
vC = 14'b0000010110000100; // vC= 1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110100; // iC=  820 
vC = 14'b0000010111111101; // vC= 1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110000; // iC=  816 
vC = 14'b0000010110101000; // vC= 1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101100; // iC=  812 
vC = 14'b0000010110010001; // vC= 1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010110; // iC=  854 
vC = 14'b0000010111001000; // vC= 1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101010; // iC=  810 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111001; // iC=  825 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010100; // iC=  788 
vC = 14'b0000011000001101; // vC= 1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000001; // iC=  897 
vC = 14'b0000010110011001; // vC= 1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100101; // iC=  933 
vC = 14'b0000010110110100; // vC= 1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001000; // iC=  840 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000001; // iC=  833 
vC = 14'b0000010111001010; // vC= 1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001001; // iC=  841 
vC = 14'b0000010110011100; // vC= 1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001001; // iC=  905 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101001; // iC=  809 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110001; // iC=  881 
vC = 14'b0000011001000110; // vC= 1606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001011; // iC=  779 
vC = 14'b0000010111010000; // vC= 1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101100; // iC=  812 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111011; // iC=  763 
vC = 14'b0000011001001001; // vC= 1609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010001; // iC=  721 
vC = 14'b0000010111000011; // vC= 1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110001; // iC=  753 
vC = 14'b0000010111100101; // vC= 1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111101; // iC=  829 
vC = 14'b0000011000110101; // vC= 1589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000000; // iC=  768 
vC = 14'b0000010110111000; // vC= 1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000001; // iC=  769 
vC = 14'b0000011000110001; // vC= 1585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111111; // iC=  703 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001101; // iC=  717 
vC = 14'b0000011000001101; // vC= 1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000000; // iC=  704 
vC = 14'b0000011001011101; // vC= 1629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000010; // iC=  706 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001010; // iC=  778 
vC = 14'b0000011000110100; // vC= 1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101011; // iC=  747 
vC = 14'b0000011000101000; // vC= 1576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001010; // iC=  778 
vC = 14'b0000011001001110; // vC= 1614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010010; // iC=  722 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010110; // iC=  790 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010111; // iC=  791 
vC = 14'b0000011001101001; // vC= 1641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111110; // iC=  766 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011001; // iC=  729 
vC = 14'b0000011000010010; // vC= 1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011100; // iC=  732 
vC = 14'b0000011001101100; // vC= 1644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100111; // iC=  615 
vC = 14'b0000011001010010; // vC= 1618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101001; // iC=  745 
vC = 14'b0000011000010111; // vC= 1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010111; // iC=  727 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011100; // iC=  668 
vC = 14'b0000011001011000; // vC= 1624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111001; // iC=  633 
vC = 14'b0000010111100011; // vC= 1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111010; // iC=  634 
vC = 14'b0000011001011011; // vC= 1627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101001; // iC=  681 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011011; // iC=  603 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000101; // iC=  645 
vC = 14'b0000011000010111; // vC= 1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000010; // iC=  578 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001110; // iC=  654 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110100; // iC=  564 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100110; // iC=  614 
vC = 14'b0000010111110111; // vC= 1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100101; // iC=  549 
vC = 14'b0000011000000110; // vC= 1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011000; // iC=  536 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000100; // iC=  644 
vC = 14'b0000011000010010; // vC= 1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000011; // iC=  579 
vC = 14'b0000011001111001; // vC= 1657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010000; // iC=  528 
vC = 14'b0000011001010101; // vC= 1621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100110; // iC=  614 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100001; // iC=  609 
vC = 14'b0000011001111110; // vC= 1662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000010; // iC=  578 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101101; // iC=  557 
vC = 14'b0000011010001111; // vC= 1679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101000; // iC=  616 
vC = 14'b0000011000001000; // vC= 1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111001; // iC=  505 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101001; // iC=  489 
vC = 14'b0000011001000011; // vC= 1603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011110; // iC=  478 
vC = 14'b0000011001110011; // vC= 1651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100011; // iC=  547 
vC = 14'b0000011001100100; // vC= 1636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001000; // iC=  456 
vC = 14'b0000011000001001; // vC= 1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111000; // iC=  568 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011001; // iC=  473 
vC = 14'b0000011000111101; // vC= 1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110000; // iC=  560 
vC = 14'b0000011000101101; // vC= 1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010100; // iC=  532 
vC = 14'b0000011000011101; // vC= 1565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001000; // iC=  456 
vC = 14'b0000011010011111; // vC= 1695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010110; // iC=  470 
vC = 14'b0000011001010101; // vC= 1621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011001; // iC=  537 
vC = 14'b0000011010011101; // vC= 1693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010110; // iC=  534 
vC = 14'b0000011010011000; // vC= 1688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010001; // iC=  401 
vC = 14'b0000011010010110; // vC= 1686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000010; // iC=  386 
vC = 14'b0000011010000001; // vC= 1665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110110; // iC=  502 
vC = 14'b0000011000111000; // vC= 1592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100001; // iC=  353 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111110; // iC=  446 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011011; // iC=  475 
vC = 14'b0000011001101110; // vC= 1646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110000; // iC=  432 
vC = 14'b0000011010011011; // vC= 1691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101001; // iC=  425 
vC = 14'b0000011010010010; // vC= 1682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111010; // iC=  378 
vC = 14'b0000011010000011; // vC= 1667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010011; // iC=  275 
vC = 14'b0000011010000001; // vC= 1665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101000; // iC=  360 
vC = 14'b0000011001011011; // vC= 1627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011010; // iC=  282 
vC = 14'b0000011001101010; // vC= 1642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111111; // iC=  383 
vC = 14'b0000011001011000; // vC= 1624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010000; // iC=  336 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110000; // iC=  304 
vC = 14'b0000011010110001; // vC= 1713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010000; // iC=  272 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100110; // iC=  230 
vC = 14'b0000011001011101; // vC= 1629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000111; // iC=  263 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011010; // iC=  282 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010110; // iC=  214 
vC = 14'b0000011001010110; // vC= 1622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011001; // iC=  217 
vC = 14'b0000011010001000; // vC= 1672 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101000; // iC=  232 
vC = 14'b0000011001111101; // vC= 1661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100001; // iC=  225 
vC = 14'b0000011001110011; // vC= 1651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100101; // iC=  165 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010100; // iC=  148 
vC = 14'b0000011010001011; // vC= 1675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111010; // iC=  122 
vC = 14'b0000011000110110; // vC= 1590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000011; // iC=   67 
vC = 14'b0000011010001111; // vC= 1679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100101; // iC=  101 
vC = 14'b0000011001111110; // vC= 1662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001101; // iC=   77 
vC = 14'b0000011010100100; // vC= 1700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110100; // iC=  -12 
vC = 14'b0000011001011100; // vC= 1628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111101000; // iC=  -24 
vC = 14'b0000011001000101; // vC= 1605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011101; // iC=  -35 
vC = 14'b0000011001100010; // vC= 1634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001111; // iC=  -49 
vC = 14'b0000011001111111; // vC= 1663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111101; // iC=   -3 
vC = 14'b0000011001010101; // vC= 1621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001010; // iC=  -54 
vC = 14'b0000011000110101; // vC= 1589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100010; // iC=  -30 
vC = 14'b0000011001000010; // vC= 1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100010; // iC= -158 
vC = 14'b0000011000110110; // vC= 1590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110001; // iC=  -79 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111001; // iC= -135 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010110; // iC= -234 
vC = 14'b0000011010000000; // vC= 1664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110100; // iC= -204 
vC = 14'b0000011001011110; // vC= 1630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000111; // iC= -249 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001101; // iC= -243 
vC = 14'b0000011010001001; // vC= 1673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011010; // iC= -294 
vC = 14'b0000011001100001; // vC= 1633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111000; // iC= -264 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001101; // iC= -307 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101101; // iC= -339 
vC = 14'b0000011010010010; // vC= 1682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110000; // iC= -400 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011101; // iC= -291 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000111; // iC= -313 
vC = 14'b0000011000000100; // vC= 1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011010; // iC= -422 
vC = 14'b0000011001010001; // vC= 1617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011000; // iC= -360 
vC = 14'b0000011000011001; // vC= 1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000011; // iC= -509 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101100; // iC= -468 
vC = 14'b0000011000110001; // vC= 1585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111011; // iC= -517 
vC = 14'b0000011000101111; // vC= 1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101001; // iC= -471 
vC = 14'b0000011001100111; // vC= 1639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100111; // iC= -473 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000101; // iC= -635 
vC = 14'b0000011000010111; // vC= 1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001000; // iC= -632 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111010; // iC= -582 
vC = 14'b0000010111111000; // vC= 1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111000; // iC= -584 
vC = 14'b0000011001000001; // vC= 1601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111111; // iC= -577 
vC = 14'b0000011001111100; // vC= 1660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111011; // iC= -645 
vC = 14'b0000011001111010; // vC= 1658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000011; // iC= -765 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100111; // iC= -665 
vC = 14'b0000010111101001; // vC= 1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111011; // iC= -773 
vC = 14'b0000011001010111; // vC= 1623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011101; // iC= -803 
vC = 14'b0000011001010001; // vC= 1617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111011; // iC= -837 
vC = 14'b0000010111111111; // vC= 1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001100; // iC= -884 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110100; // iC= -908 
vC = 14'b0000011001011011; // vC= 1627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110011; // iC= -845 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101000; // iC= -792 
vC = 14'b0000010111011100; // vC= 1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011010; // iC= -934 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001111; // iC= -881 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011010; // iC= -870 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000110; // iC= -954 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111111; // iC=-1025 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101010; // iC=-1046 
vC = 14'b0000010110100101; // vC= 1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001100; // iC=-1012 
vC = 14'b0000011000111000; // vC= 1592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111110; // iC=-1026 
vC = 14'b0000010111010111; // vC= 1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010110; // iC=-1066 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000110; // iC=-1018 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101110; // iC=-1042 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111110; // iC=-1154 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100100; // iC=-1052 
vC = 14'b0000010111111101; // vC= 1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100000; // iC=-1056 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110101; // iC=-1163 
vC = 14'b0000010101111001; // vC= 1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011101; // iC=-1187 
vC = 14'b0000010111100110; // vC= 1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010110; // iC=-1130 
vC = 14'b0000010110100101; // vC= 1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b0000010110001011; // vC= 1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011110; // iC=-1250 
vC = 14'b0000010110011111; // vC= 1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010111; // iC=-1257 
vC = 14'b0000010110001010; // vC= 1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b0000010110101010; // vC= 1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101011; // iC=-1301 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100001; // iC=-1247 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100011; // iC=-1309 
vC = 14'b0000010101011110; // vC= 1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001010; // iC=-1334 
vC = 14'b0000010101010101; // vC= 1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000100; // iC=-1340 
vC = 14'b0000010110101000; // vC= 1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100011; // iC=-1373 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001101; // iC=-1395 
vC = 14'b0000010110110011; // vC= 1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001001; // iC=-1399 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b0000010111000101; // vC= 1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011110; // iC=-1314 
vC = 14'b0000010101101001; // vC= 1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001000; // iC=-1336 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b0000010100100000; // vC= 1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111001; // iC=-1479 
vC = 14'b0000010101101010; // vC= 1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110001; // iC=-1359 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b0000010110011001; // vC= 1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b0000010110011000; // vC= 1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110010; // iC=-1486 
vC = 14'b0000010100010000; // vC= 1296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010011; // iC=-1517 
vC = 14'b0000010101010101; // vC= 1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b0000010101001101; // vC= 1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011111; // iC=-1505 
vC = 14'b0000010101101100; // vC= 1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101111; // iC=-1489 
vC = 14'b0000010101000111; // vC= 1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b0000010100011011; // vC= 1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111110; // iC=-1538 
vC = 14'b0000010101001001; // vC= 1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010100; // iC=-1580 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b0000010101100011; // vC= 1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001110; // iC=-1586 
vC = 14'b0000010011101001; // vC= 1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101100; // iC=-1556 
vC = 14'b0000010100110000; // vC= 1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b0000010010110001; // vC= 1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b0000010100101001; // vC= 1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101111; // iC=-1617 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b0000010010011111; // vC= 1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b0000010011111100; // vC= 1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110111; // iC=-1545 
vC = 14'b0000010010011110; // vC= 1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100100; // iC=-1692 
vC = 14'b0000010010110111; // vC= 1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b0000010010011010; // vC= 1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b0000010100001101; // vC= 1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b0000010010110110; // vC= 1206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000010010100111; // vC= 1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b0000010010100111; // vC= 1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000010010011101; // vC= 1181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000101; // iC=-1595 
vC = 14'b0000010001100101; // vC= 1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000010001101100; // vC= 1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010000; // iC=-1648 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b0000010001101000; // vC= 1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b0000010001101000; // vC= 1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000010010010111; // vC= 1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b0000010001001000; // vC= 1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b0000010010101100; // vC= 1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000111; // iC=-1657 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101110; // iC=-1618 
vC = 14'b0000010010100101; // vC= 1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000010000011101; // vC= 1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000010010010011; // vC= 1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000010000000100; // vC= 1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000100; // iC=-1724 
vC = 14'b0000010000101010; // vC= 1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011010; // iC=-1702 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000001111111000; // vC= 1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000001111111010; // vC= 1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b0000001111101110; // vC= 1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b0000010000010100; // vC= 1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b0000001111110100; // vC= 1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000010000000001; // vC= 1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000001111111010; // vC= 1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000001111110101; // vC= 1013 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000010000101010; // vC= 1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001110100111; // vC=  935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b0000001111111101; // vC= 1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011010; // iC=-1702 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000001110110101; // vC=  949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000001111010011; // vC=  979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101001; // iC=-1815 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000001111111010; // vC= 1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011010; // iC=-1830 
vC = 14'b0000001111100000; // vC=  992 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101101; // iC=-1683 
vC = 14'b0000001101111010; // vC=  890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000001111001101; // vC=  973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b0000001111100100; // vC=  996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001111010110; // vC=  982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000001101001001; // vC=  841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000001110111011; // vC=  955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b0000001100101110; // vC=  814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b0000001101111110; // vC=  894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b0000001110000100; // vC=  900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000001100011001; // vC=  793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011101; // iC=-1699 
vC = 14'b0000001101100010; // vC=  866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b0000001101001100; // vC=  844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000000; // iC=-1792 
vC = 14'b0000001110010101; // vC=  917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000001100111011; // vC=  827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000001101011010; // vC=  858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001010; // iC=-1846 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000001011110111; // vC=  759 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000001100100101; // vC=  805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000001100110101; // vC=  821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110011; // iC=-1869 
vC = 14'b0000001011001001; // vC=  713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000001101000011; // vC=  835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000001101001000; // vC=  840 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b0000001100000001; // vC=  769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b0000001010101010; // vC=  682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000001100101111; // vC=  815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000001011110011; // vC=  755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000001100011001; // vC=  793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000001100101111; // vC=  815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111110; // iC=-1858 
vC = 14'b0000001010001001; // vC=  649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000001011011000; // vC=  728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b0000001100010101; // vC=  789 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000001010010000; // vC=  656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000001011100011; // vC=  739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000001010110001; // vC=  689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101100; // iC=-1876 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000001011110110; // vC=  758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000001010010001; // vC=  657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101011; // iC=-1877 
vC = 14'b0000001001100100; // vC=  612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000001011010011; // vC=  723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100111; // iC=-1881 
vC = 14'b0000001001010001; // vC=  593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000001000111101; // vC=  573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101100; // iC=-1876 
vC = 14'b0000001001011101; // vC=  605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000001001011101; // vC=  605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b0000001001100110; // vC=  614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100001; // iC=-1887 
vC = 14'b0000001000111111; // vC=  575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111001; // iC=-1863 
vC = 14'b0000001001111101; // vC=  637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000001000001111; // vC=  527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000001000100010; // vC=  546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000001001101001; // vC=  617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000001000000100; // vC=  516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000001001111010; // vC=  634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000001000011111; // vC=  543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000001000000010; // vC=  514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110000; // iC=-1872 
vC = 14'b0000001000010101; // vC=  533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000001000100000; // vC=  544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010110; // iC=-1898 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011110; // iC=-1890 
vC = 14'b0000001000111001; // vC=  569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000000111111100; // vC=  508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001111; // iC=-1841 
vC = 14'b0000000110111101; // vC=  445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000001000100111; // vC=  551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000000110110101; // vC=  437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110010; // iC=-1806 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000000101110010; // vC=  370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111110; // iC=-1858 
vC = 14'b0000000110110000; // vC=  432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000000111011111; // vC=  479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000000110100011; // vC=  419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000000111010010; // vC=  466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000000; // iC=-1792 
vC = 14'b0000000111000011; // vC=  451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100001; // iC=-1887 
vC = 14'b0000000101111100; // vC=  380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101001; // iC=-1879 
vC = 14'b0000000101000100; // vC=  324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000000101011110; // vC=  350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100000; // iC=-1888 
vC = 14'b0000000110100000; // vC=  416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000000101001000; // vC=  328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000000100110011; // vC=  307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101011; // iC=-1877 
vC = 14'b0000000101111101; // vC=  381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011001; // iC=-1895 
vC = 14'b0000000110101011; // vC=  427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100000; // iC=-1888 
vC = 14'b0000000100010111; // vC=  279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000111; // iC=-1849 
vC = 14'b0000000100011010; // vC=  282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011010; // iC=-1894 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000000101111001; // vC=  377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000000011101011; // vC=  235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000000100110000; // vC=  304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000000100111110; // vC=  318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000000101100001; // vC=  353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100001; // iC=-1887 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110010; // iC=-1806 
vC = 14'b0000000101000100; // vC=  324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000000100111101; // vC=  317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000000100110011; // vC=  307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000000011100001; // vC=  225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000000011101001; // vC=  233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000000100101001; // vC=  297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000000011010001; // vC=  209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000000010100100; // vC=  164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000000010111100; // vC=  188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000000001100111; // vC=  103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000000001111000; // vC=  120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000111; // iC=-1849 
vC = 14'b0000000011011101; // vC=  221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000000001100000; // vC=   96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000000001000010; // vC=   66 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000000000110111; // vC=   55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000000000011100; // vC=   28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000000001110011; // vC=  115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000000000100000; // vC=   32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000000001000100; // vC=   68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000000000101000; // vC=   40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000000010001000; // vC=  136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000000001101110; // vC=  110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b0000000000100000; // vC=   32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000000001111001; // vC=  121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000000000110100; // vC=   52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000000000011101; // vC=   29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000000000001011; // vC=   11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000000000101110; // vC=   46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000000001010000; // vC=   80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101001; // iC=-1815 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111111; // iC=-1857 
vC = 14'b1111111111011000; // vC=  -40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b1111111110110011; // vC=  -77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000000001000101; // vC=   69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b1111111111011011; // vC=  -37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000000000011001; // vC=   25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b1111111111000001; // vC=  -63 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b1111111111011001; // vC=  -39 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b1111111111000101; // vC=  -59 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b1111111111101101; // vC=  -19 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b1111111111110110; // vC=  -10 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b1111111111010010; // vC=  -46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b1111111110111001; // vC=  -71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b1111111101111100; // vC= -132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b1111111111001101; // vC=  -51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b1111111101111010; // vC= -134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000000; // iC=-1792 
vC = 14'b1111111111001100; // vC=  -52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011011; // iC=-1829 
vC = 14'b1111111101100000; // vC= -160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011101; // iC=-1827 
vC = 14'b1111111101011010; // vC= -166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b1111111101110001; // vC= -143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b1111111110111101; // vC=  -67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b1111111101011101; // vC= -163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101000; // iC=-1688 
vC = 14'b1111111100101000; // vC= -216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b1111111101000110; // vC= -186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b1111111100100010; // vC= -222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b1111111100111100; // vC= -196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b1111111101100100; // vC= -156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111101; // iC=-1667 
vC = 14'b1111111100111011; // vC= -197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b1111111100001011; // vC= -245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100000; // iC=-1760 
vC = 14'b1111111100110111; // vC= -201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b1111111101010101; // vC= -171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b1111111110000001; // vC= -127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b1111111101011010; // vC= -166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111011; // iC=-1797 
vC = 14'b1111111101111011; // vC= -133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b1111111100101111; // vC= -209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b1111111011101001; // vC= -279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b1111111101001110; // vC= -178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b1111111100101111; // vC= -209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b1111111011011100; // vC= -292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001000; // iC=-1656 
vC = 14'b1111111010111001; // vC= -327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b1111111011100110; // vC= -282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b1111111100101001; // vC= -215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b1111111011010101; // vC= -299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b1111111011101100; // vC= -276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b1111111010010110; // vC= -362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b1111111010110100; // vC= -332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101111; // iC=-1617 
vC = 14'b1111111100000010; // vC= -254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111100; // iC=-1668 
vC = 14'b1111111010111000; // vC= -328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b1111111011110001; // vC= -271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b1111111001111010; // vC= -390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110001; // iC=-1679 
vC = 14'b1111111011100110; // vC= -282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b1111111010110100; // vC= -332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101111; // iC=-1617 
vC = 14'b1111111010011101; // vC= -355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b1111111001101000; // vC= -408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b1111111011001000; // vC= -312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111101; // iC=-1667 
vC = 14'b1111111001011101; // vC= -419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011001; // iC=-1639 
vC = 14'b1111111001100000; // vC= -416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b1111111011000000; // vC= -320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b1111111001010001; // vC= -431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b1111111000110111; // vC= -457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010111; // iC=-1641 
vC = 14'b1111111001000011; // vC= -445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b1111111010100100; // vC= -348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101101; // iC=-1619 
vC = 14'b1111111010000111; // vC= -377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001100; // iC=-1588 
vC = 14'b1111111010110000; // vC= -336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001101; // iC=-1587 
vC = 14'b1111111001101011; // vC= -405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011010; // iC=-1702 
vC = 14'b1111111010101101; // vC= -339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b1111111000110000; // vC= -464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111111; // iC=-1665 
vC = 14'b1111111001101110; // vC= -402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b1111111000110010; // vC= -462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b1111111001001000; // vC= -440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b1111111000010001; // vC= -495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b1111110111111111; // vC= -513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110001; // iC=-1615 
vC = 14'b1111110111110110; // vC= -522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110100; // iC=-1612 
vC = 14'b1111111000101110; // vC= -466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b1111111001110110; // vC= -394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b1111111000111001; // vC= -455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101000; // iC=-1624 
vC = 14'b1111111001001000; // vC= -440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b1111111000011001; // vC= -487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b1111110111101110; // vC= -530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b1111111000100000; // vC= -480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b1111111001000110; // vC= -442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110111; // iC=-1673 
vC = 14'b1111110111101111; // vC= -529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b1111111000011010; // vC= -486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b1111110111010001; // vC= -559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b1111110111111100; // vC= -516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111101; // iC=-1603 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b1111110111100110; // vC= -538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b1111110110101110; // vC= -594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011100; // iC=-1572 
vC = 14'b1111111000000100; // vC= -508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110000; // iC=-1552 
vC = 14'b1111110110010000; // vC= -624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b1111110110010100; // vC= -620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b1111110101111011; // vC= -645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b1111110110011011; // vC= -613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b1111110101101001; // vC= -663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b1111110111011101; // vC= -547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111100; // iC=-1604 
vC = 14'b1111110101110010; // vC= -654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b1111110101011010; // vC= -678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b1111110111000111; // vC= -569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010100; // iC=-1580 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110101; // iC=-1483 
vC = 14'b1111110110000010; // vC= -638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001010; // iC=-1462 
vC = 14'b1111110110111100; // vC= -580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b1111110101011001; // vC= -679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b1111110101101010; // vC= -662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010010; // iC=-1582 
vC = 14'b1111110100101001; // vC= -727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000000; // iC=-1472 
vC = 14'b1111110101110100; // vC= -652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b1111110101110001; // vC= -655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b1111110110000101; // vC= -635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001100; // iC=-1524 
vC = 14'b1111110101100101; // vC= -667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001111; // iC=-1521 
vC = 14'b1111110110001100; // vC= -628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b1111110101011001; // vC= -679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101011; // iC=-1493 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111101; // iC=-1539 
vC = 14'b1111110100100100; // vC= -732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b1111110100011111; // vC= -737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b1111110100010000; // vC= -752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010110; // iC=-1450 
vC = 14'b1111110101100110; // vC= -666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b1111110101111101; // vC= -643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b1111110011111011; // vC= -773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111010; // iC=-1478 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b1111110101101110; // vC= -658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111101; // iC=-1539 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100101; // iC=-1435 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011110; // iC=-1378 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000110; // iC=-1402 
vC = 14'b1111110011000111; // vC= -825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101000; // iC=-1368 
vC = 14'b1111110011101100; // vC= -788 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111100; // iC=-1476 
vC = 14'b1111110101000000; // vC= -704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010111; // iC=-1513 
vC = 14'b1111110010100110; // vC= -858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111010; // iC=-1414 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101011; // iC=-1493 
vC = 14'b1111110010110010; // vC= -846 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001010; // iC=-1398 
vC = 14'b1111110100010001; // vC= -751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111010; // iC=-1350 
vC = 14'b1111110011011100; // vC= -804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010010; // iC=-1390 
vC = 14'b1111110011011001; // vC= -807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000011; // iC=-1405 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b1111110100001000; // vC= -760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110010; // iC=-1486 
vC = 14'b1111110011110011; // vC= -781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b1111110010110111; // vC= -841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001100; // iC=-1332 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100001; // iC=-1375 
vC = 14'b1111110010011000; // vC= -872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001000; // iC=-1336 
vC = 14'b1111110010100101; // vC= -859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001101; // iC=-1331 
vC = 14'b1111110011000110; // vC= -826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000000; // iC=-1344 
vC = 14'b1111110010011111; // vC= -865 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100001; // iC=-1311 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011111; // iC=-1377 
vC = 14'b1111110011001111; // vC= -817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011100; // iC=-1444 
vC = 14'b1111110001001001; // vC= -951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111110; // iC=-1346 
vC = 14'b1111110010110001; // vC= -847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010101; // iC=-1323 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010100; // iC=-1388 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001100; // iC=-1332 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111101; // iC=-1411 
vC = 14'b1111110001000101; // vC= -955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101010; // iC=-1366 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011101; // iC=-1379 
vC = 14'b1111110001011111; // vC= -929 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101000; // iC=-1368 
vC = 14'b1111110010011001; // vC= -871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010101; // iC=-1259 
vC = 14'b1111110001110011; // vC= -909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101101; // iC=-1363 
vC = 14'b1111110001001110; // vC= -946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011111; // iC=-1313 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b1111110000110010; // vC= -974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101100; // iC=-1364 
vC = 14'b1111110001010111; // vC= -937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110110; // iC=-1354 
vC = 14'b1111110001010101; // vC= -939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111100; // iC=-1284 
vC = 14'b1111110001000010; // vC= -958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100011; // iC=-1309 
vC = 14'b1111110000010111; // vC=-1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110101; // iC=-1291 
vC = 14'b1111110001110111; // vC= -905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110010; // iC=-1294 
vC = 14'b1111110001101111; // vC= -913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101010; // iC=-1238 
vC = 14'b1111110000100001; // vC= -991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111001; // iC=-1223 
vC = 14'b1111110000111101; // vC= -963 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001010; // iC=-1270 
vC = 14'b1111110001111001; // vC= -903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001111; // iC=-1265 
vC = 14'b1111110000100011; // vC= -989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111110001001011; // vC= -949 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010000; // iC=-1200 
vC = 14'b1111101111100000; // vC=-1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001001; // iC=-1207 
vC = 14'b1111110001100010; // vC= -926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100000; // iC=-1184 
vC = 14'b1111110000000110; // vC=-1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011110; // iC=-1186 
vC = 14'b1111101111010011; // vC=-1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b1111101111110011; // vC=-1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010110; // iC=-1258 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111110; // iC=-1154 
vC = 14'b1111110000000011; // vC=-1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100111; // iC=-1241 
vC = 14'b1111101110111101; // vC=-1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101001; // iC=-1175 
vC = 14'b1111101111101011; // vC=-1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b1111101111001111; // vC=-1073 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100110; // iC=-1178 
vC = 14'b1111101111100110; // vC=-1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001100; // iC=-1140 
vC = 14'b1111101111111000; // vC=-1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001001; // iC=-1271 
vC = 14'b1111110000001101; // vC=-1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000100; // iC=-1148 
vC = 14'b1111101110111010; // vC=-1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011010; // iC=-1126 
vC = 14'b1111101110011011; // vC=-1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010000; // iC=-1200 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001100; // iC=-1140 
vC = 14'b1111101111010110; // vC=-1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011000; // iC=-1192 
vC = 14'b1111101111010100; // vC=-1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101001; // iC=-1175 
vC = 14'b1111101111100111; // vC=-1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101001; // iC=-1175 
vC = 14'b1111101110111000; // vC=-1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100111; // iC=-1113 
vC = 14'b1111110000001100; // vC=-1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100100; // iC=-1180 
vC = 14'b1111101110110111; // vC=-1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000100; // iC=-1148 
vC = 14'b1111101101110011; // vC=-1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111011; // iC=-1221 
vC = 14'b1111101101101111; // vC=-1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011100; // iC=-1188 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110100; // iC=-1100 
vC = 14'b1111101111000101; // vC=-1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001101; // iC=-1203 
vC = 14'b1111101110111000; // vC=-1096 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101111; // iC=-1105 
vC = 14'b1111101111001001; // vC=-1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100100; // iC=-1180 
vC = 14'b1111101111001101; // vC=-1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001010; // iC=-1206 
vC = 14'b1111101101010101; // vC=-1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001001; // iC=-1143 
vC = 14'b1111101111101100; // vC=-1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000110; // iC=-1082 
vC = 14'b1111101111100111; // vC=-1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011010; // iC=-1062 
vC = 14'b1111101101010101; // vC=-1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011100; // iC=-1060 
vC = 14'b1111101110010111; // vC=-1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001010; // iC=-1078 
vC = 14'b1111101101110000; // vC=-1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001100; // iC=-1140 
vC = 14'b1111101101100100; // vC=-1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011110; // iC=-1122 
vC = 14'b1111101110100111; // vC=-1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011001; // iC=-1127 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011000; // iC=-1064 
vC = 14'b1111101101111100; // vC=-1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000011; // iC=-1149 
vC = 14'b1111101100111111; // vC=-1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110010; // iC=-1102 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000100; // iC=-1148 
vC = 14'b1111101110001011; // vC=-1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100100; // iC=-1052 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000001; // iC=-1023 
vC = 14'b1111101110011110; // vC=-1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111001; // iC=-1095 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100010; // iC=-1054 
vC = 14'b1111101101100010; // vC=-1182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101011; // iC=-1045 
vC = 14'b1111101110100010; // vC=-1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011001; // iC= -999 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110111; // iC=-1097 
vC = 14'b1111101101000001; // vC=-1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011011; // iC= -997 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101010; // iC=-1046 
vC = 14'b1111101101001101; // vC=-1203 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110100; // iC=-1036 
vC = 14'b1111101100110101; // vC=-1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100110; // iC= -986 
vC = 14'b1111101101010011; // vC=-1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100001; // iC= -991 
vC = 14'b1111101011111010; // vC=-1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100001; // iC= -927 
vC = 14'b1111101100100011; // vC=-1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100000; // iC= -928 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111101101000000; // vC=-1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011101; // iC= -931 
vC = 14'b1111101101011011; // vC=-1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010001; // iC= -943 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101111; // iC= -913 
vC = 14'b1111101100001010; // vC=-1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100000; // iC= -928 
vC = 14'b1111101101000011; // vC=-1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000011; // iC= -957 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111101; // iC= -899 
vC = 14'b1111101011101110; // vC=-1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010100; // iC= -940 
vC = 14'b1111101011011111; // vC=-1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010111; // iC= -873 
vC = 14'b1111101101101011; // vC=-1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110111; // iC= -969 
vC = 14'b1111101101101010; // vC=-1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011010; // iC= -870 
vC = 14'b1111101100001101; // vC=-1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110110; // iC= -906 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011110; // iC= -866 
vC = 14'b1111101100001101; // vC=-1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000100; // iC= -956 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000100; // iC= -956 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011010; // iC= -998 
vC = 14'b1111101011100010; // vC=-1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110011; // iC= -845 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111001; // iC= -967 
vC = 14'b1111101010110001; // vC=-1359 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110011; // iC= -973 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000101; // iC= -891 
vC = 14'b1111101011011100; // vC=-1316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110000; // iC= -912 
vC = 14'b1111101011111101; // vC=-1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000111; // iC= -889 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011111; // iC= -801 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011101; // iC= -867 
vC = 14'b1111101011100010; // vC=-1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011001; // iC= -807 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100110; // iC= -858 
vC = 14'b1111101100010011; // vC=-1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101100; // iC= -916 
vC = 14'b1111101010011010; // vC=-1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010001; // iC= -815 
vC = 14'b1111101100010000; // vC=-1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000100; // iC= -892 
vC = 14'b1111101010100001; // vC=-1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111011; // iC= -901 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011010; // iC= -806 
vC = 14'b1111101100010111; // vC=-1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010000; // iC= -880 
vC = 14'b1111101011000011; // vC=-1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011111; // iC= -865 
vC = 14'b1111101011110110; // vC=-1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101101; // iC= -787 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101001; // iC= -791 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100100; // iC= -796 
vC = 14'b1111101010010111; // vC=-1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110100; // iC= -844 
vC = 14'b1111101011010101; // vC=-1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101101; // iC= -723 
vC = 14'b1111101010001101; // vC=-1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111010; // iC= -774 
vC = 14'b1111101010110011; // vC=-1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011101; // iC= -867 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000000; // iC= -768 
vC = 14'b1111101010011101; // vC=-1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001101; // iC= -819 
vC = 14'b1111101010001010; // vC=-1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110001; // iC= -847 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000001; // iC= -703 
vC = 14'b1111101011101100; // vC=-1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100110; // iC= -730 
vC = 14'b1111101010010001; // vC=-1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011010; // iC= -742 
vC = 14'b1111101010110000; // vC=-1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101111; // iC= -785 
vC = 14'b1111101010110011; // vC=-1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101100; // iC= -788 
vC = 14'b1111101010010000; // vC=-1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101011; // iC= -789 
vC = 14'b1111101011010001; // vC=-1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011000; // iC= -680 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110001; // iC= -783 
vC = 14'b1111101011000011; // vC=-1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110001; // iC= -719 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000001; // iC= -703 
vC = 14'b1111101011011110; // vC=-1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000111; // iC= -697 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000110; // iC= -762 
vC = 14'b1111101001111111; // vC=-1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000011; // iC= -637 
vC = 14'b1111101011000100; // vC=-1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001101; // iC= -691 
vC = 14'b1111101010010110; // vC=-1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110010; // iC= -718 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010000; // iC= -624 
vC = 14'b1111101010001101; // vC=-1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000110; // iC= -698 
vC = 14'b1111101010001111; // vC=-1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010101; // iC= -683 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111001; // iC= -711 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111000; // iC= -712 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100001; // iC= -671 
vC = 14'b1111101010111101; // vC=-1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101001; // iC= -727 
vC = 14'b1111101010010100; // vC=-1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001001; // iC= -695 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010010; // iC= -558 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b1111101011000001; // vC=-1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101010; // iC= -662 
vC = 14'b1111101010100010; // vC=-1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100010; // iC= -670 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001111; // iC= -625 
vC = 14'b1111101001110011; // vC=-1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111101; // iC= -579 
vC = 14'b1111101010111101; // vC=-1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101110; // iC= -530 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111010; // iC= -646 
vC = 14'b1111101001101001; // vC=-1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011001; // iC= -615 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110101; // iC= -523 
vC = 14'b1111101010001110; // vC=-1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010100; // iC= -620 
vC = 14'b1111101010001000; // vC=-1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010000; // iC= -496 
vC = 14'b1111101010011010; // vC=-1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000010; // iC= -574 
vC = 14'b1111101000110000; // vC=-1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011001; // iC= -487 
vC = 14'b1111101010010110; // vC=-1386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100110; // iC= -602 
vC = 14'b1111101000111100; // vC=-1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011100; // iC= -612 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001101; // iC= -627 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011101; // iC= -547 
vC = 14'b1111101000010010; // vC=-1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110100; // iC= -460 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101000; // iC= -536 
vC = 14'b1111101000001110; // vC=-1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101100; // iC= -468 
vC = 14'b1111101001111100; // vC=-1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000001; // iC= -575 
vC = 14'b1111101000011010; // vC=-1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110101; // iC= -587 
vC = 14'b1111101000000001; // vC=-1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010011; // iC= -493 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111110; // iC= -450 
vC = 14'b1111101001010100; // vC=-1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000111; // iC= -569 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001101; // iC= -563 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001001; // iC= -439 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010100; // iC= -556 
vC = 14'b1111101000011100; // vC=-1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100111; // iC= -409 
vC = 14'b1111101001011000; // vC=-1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110010; // iC= -398 
vC = 14'b1111100111110000; // vC=-1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000111010; // iC= -454 
vC = 14'b1111101000110011; // vC=-1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011100; // iC= -484 
vC = 14'b1111101001101010; // vC=-1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010110; // iC= -490 
vC = 14'b1111100111111001; // vC=-1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101011; // iC= -469 
vC = 14'b1111101010001001; // vC=-1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000111; // iC= -377 
vC = 14'b1111101000000110; // vC=-1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110100; // iC= -396 
vC = 14'b1111101000011000; // vC=-1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111101; // iC= -387 
vC = 14'b1111100111110101; // vC=-1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110010; // iC= -398 
vC = 14'b1111101000000000; // vC=-1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011000001; // iC= -319 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110000; // iC= -400 
vC = 14'b1111101000110000; // vC=-1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010001; // iC= -431 
vC = 14'b1111101001101010; // vC=-1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001010; // iC= -310 
vC = 14'b1111100111101110; // vC=-1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101101; // iC= -339 
vC = 14'b1111100111101100; // vC=-1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010111; // iC= -361 
vC = 14'b1111101000110100; // vC=-1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100111; // iC= -409 
vC = 14'b1111101000111011; // vC=-1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001110100; // iC= -396 
vC = 14'b1111100111101000; // vC=-1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101101; // iC= -339 
vC = 14'b1111101001001101; // vC=-1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010011; // iC= -237 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100101; // iC= -347 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000010; // iC= -190 
vC = 14'b1111101000111100; // vC=-1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110110; // iC= -266 
vC = 14'b1111101000000010; // vC=-1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001001; // iC= -311 
vC = 14'b1111100111100001; // vC=-1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110101; // iC= -203 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110110; // iC= -266 
vC = 14'b1111101000010000; // vC=-1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111010; // iC= -198 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001000; // iC= -184 
vC = 14'b1111101000010001; // vC=-1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101000; // iC= -216 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101001; // iC= -151 
vC = 14'b1111100111101111; // vC=-1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010100; // iC= -172 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001011; // iC=  -53 
vC = 14'b1111100111111011; // vC=-1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000101; // iC= -123 
vC = 14'b1111101001001001; // vC=-1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001101; // iC= -115 
vC = 14'b1111101000100100; // vC=-1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110010; // iC=  -14 
vC = 14'b1111101000000110; // vC=-1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011010; // iC=  -38 
vC = 14'b1111100111101001; // vC=-1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110110001; // iC=  -79 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010100; // iC=   20 
vC = 14'b1111100111100111; // vC=-1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000100; // iC=  -60 
vC = 14'b1111101000101011; // vC=-1493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111100100; // iC=  -28 
vC = 14'b1111101000000111; // vC=-1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110100; // iC=  -12 
vC = 14'b1111101001101000; // vC=-1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100100; // iC=  100 
vC = 14'b1111101000000000; // vC=-1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100110; // iC=  102 
vC = 14'b1111101001000011; // vC=-1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010000; // iC=   80 
vC = 14'b1111100111111110; // vC=-1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001001; // iC=  201 
vC = 14'b1111101000011010; // vC=-1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011001; // iC=  217 
vC = 14'b1111101001110011; // vC=-1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100001; // iC=   97 
vC = 14'b1111101000100101; // vC=-1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111010; // iC=  122 
vC = 14'b1111101000011001; // vC=-1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100111; // iC=  167 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010111; // iC=  279 
vC = 14'b1111101000011111; // vC=-1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111111; // iC=  255 
vC = 14'b1111101001101010; // vC=-1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010010; // iC=  274 
vC = 14'b1111101000100011; // vC=-1501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110110; // iC=  310 
vC = 14'b1111101000110001; // vC=-1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110111; // iC=  247 
vC = 14'b1111101000010000; // vC=-1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011010; // iC=  346 
vC = 14'b1111101000010100; // vC=-1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010100; // iC=  340 
vC = 14'b1111101000001100; // vC=-1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100001; // iC=  417 
vC = 14'b1111100111101001; // vC=-1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100111; // iC=  423 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011000; // iC=  472 
vC = 14'b1111100111101000; // vC=-1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111111; // iC=  447 
vC = 14'b1111101001010100; // vC=-1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110111; // iC=  439 
vC = 14'b1111101000000111; // vC=-1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000100; // iC=  580 
vC = 14'b1111101001001001; // vC=-1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001000; // iC=  456 
vC = 14'b1111101000000001; // vC=-1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101011; // iC=  491 
vC = 14'b1111101001000000; // vC=-1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000111; // iC=  583 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011001; // iC=  601 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110001; // iC=  561 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011001; // iC=  665 
vC = 14'b1111101000000010; // vC=-1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100011; // iC=  739 
vC = 14'b1111101001001110; // vC=-1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111011; // iC=  699 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111101; // iC=  701 
vC = 14'b1111101000100001; // vC=-1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010011; // iC=  723 
vC = 14'b1111101000100101; // vC=-1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110101; // iC=  821 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010011; // iC=  787 
vC = 14'b1111101000001000; // vC=-1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111111; // iC=  831 
vC = 14'b1111101000010010; // vC=-1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010000; // iC=  912 
vC = 14'b1111101001111101; // vC=-1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001110; // iC=  910 
vC = 14'b1111101001011111; // vC=-1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011000; // iC=  856 
vC = 14'b1111101000010011; // vC=-1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101111; // iC=  943 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100100; // iC=  868 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011010; // iC=  986 
vC = 14'b1111101010001111; // vC=-1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011000; // iC=  984 
vC = 14'b1111101000101111; // vC=-1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111101; // iC= 1085 
vC = 14'b1111101010011000; // vC=-1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000101; // iC=  965 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011111; // iC= 1119 
vC = 14'b1111101001010001; // vC=-1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100111; // iC=  999 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001000; // iC= 1160 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001100; // iC= 1036 
vC = 14'b1111101001001101; // vC=-1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110011; // iC= 1203 
vC = 14'b1111101010001000; // vC=-1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110010; // iC= 1138 
vC = 14'b1111101010000010; // vC=-1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110101; // iC= 1141 
vC = 14'b1111101001011001; // vC=-1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011000; // iC= 1240 
vC = 14'b1111101010001110; // vC=-1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000111; // iC= 1159 
vC = 14'b1111101001001110; // vC=-1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011100; // iC= 1180 
vC = 14'b1111101011110010; // vC=-1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001010; // iC= 1226 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110010; // iC= 1202 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011000; // iC= 1240 
vC = 14'b1111101011101110; // vC=-1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111001; // iC= 1273 
vC = 14'b1111101010011011; // vC=-1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101001; // iC= 1257 
vC = 14'b1111101010110011; // vC=-1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010111; // iC= 1431 
vC = 14'b1111101011101000; // vC=-1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010001; // iC= 1425 
vC = 14'b1111101011010011; // vC=-1325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011101; // iC= 1309 
vC = 14'b1111101011111110; // vC=-1282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010011; // iC= 1363 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000110; // iC= 1478 
vC = 14'b1111101010011011; // vC=-1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101110; // iC= 1390 
vC = 14'b1111101010100101; // vC=-1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011010; // iC= 1434 
vC = 14'b1111101100011001; // vC=-1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111011; // iC= 1467 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001010; // iC= 1418 
vC = 14'b1111101011101011; // vC=-1301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100000; // iC= 1504 
vC = 14'b1111101100111100; // vC=-1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b1111101011110001; // vC=-1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110101; // iC= 1589 
vC = 14'b1111101100010000; // vC=-1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000000; // iC= 1600 
vC = 14'b1111101011001110; // vC=-1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111001; // iC= 1593 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100000; // iC= 1504 
vC = 14'b1111101101100000; // vC=-1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110001; // iC= 1649 
vC = 14'b1111101100010010; // vC=-1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001011; // iC= 1611 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010011; // iC= 1619 
vC = 14'b1111101101001100; // vC=-1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101001; // iC= 1641 
vC = 14'b1111101101001010; // vC=-1206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b1111101101011011; // vC=-1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b1111101110001100; // vC=-1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101011; // iC= 1643 
vC = 14'b1111101011110111; // vC=-1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110001; // iC= 1713 
vC = 14'b1111101100010100; // vC=-1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000001; // iC= 1665 
vC = 14'b1111101110001101; // vC=-1139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000110; // iC= 1798 
vC = 14'b1111101101111010; // vC=-1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b1111101100110111; // vC=-1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b1111101100010001; // vC=-1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001101; // iC= 1677 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b1111101101010111; // vC=-1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b1111101110110100; // vC=-1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b1111101110000001; // vC=-1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b1111101101110100; // vC=-1164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b1111101101101111; // vC=-1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111101110110000; // vC=-1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010100; // iC= 1876 
vC = 14'b1111101110000001; // vC=-1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010100; // iC= 1748 
vC = 14'b1111101111011100; // vC=-1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b1111101110000111; // vC=-1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100010; // iC= 1762 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b1111101111010010; // vC=-1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100010; // iC= 1826 
vC = 14'b1111101101111001; // vC=-1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b1111101111011000; // vC=-1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111011; // iC= 1851 
vC = 14'b1111101101111111; // vC=-1153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010101; // iC= 1813 
vC = 14'b1111101111001001; // vC=-1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111101111111100; // vC=-1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111110000100110; // vC= -986 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111101110110101; // vC=-1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b1111101110111001; // vC=-1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000111; // iC= 1863 
vC = 14'b1111101111101000; // vC=-1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b1111101111100000; // vC=-1056 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111101111100001; // vC=-1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b1111110001001100; // vC= -948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b1111110000011101; // vC= -995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b1111101111100011; // vC=-1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110001; // iC= 1841 
vC = 14'b1111101111100100; // vC=-1052 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001111; // iC= 1871 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110101; // iC= 1845 
vC = 14'b1111110000001111; // vC=-1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111110010001111; // vC= -881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b1111110001101000; // vC= -920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b1111110000100001; // vC= -991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111110000001100; // vC=-1012 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000100; // iC= 1924 
vC = 14'b1111110000010100; // vC=-1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111110010000001; // vC= -895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111110000110010; // vC= -974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111110001001101; // vC= -947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b1111110010010111; // vC= -873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001001; // iC= 1865 
vC = 14'b1111110001000101; // vC= -955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b1111110011011110; // vC= -802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b1111110001110101; // vC= -907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101111; // iC= 1903 
vC = 14'b1111110011101001; // vC= -791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011011; // iC= 2011 
vC = 14'b1111110010111100; // vC= -836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111110001100110; // vC= -922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b1111110010011100; // vC= -868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b1111110010010001; // vC= -879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111110010000101; // vC= -891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111110100000010; // vC= -766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111110011101111; // vC= -785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b1111110100001100; // vC= -756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111001; // iC= 2041 
vC = 14'b1111110100111000; // vC= -712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111110011100010; // vC= -798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111110100110001; // vC= -719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b1111110011111100; // vC= -772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111110011110000; // vC= -784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b1111110100001101; // vC= -755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b1111110101001010; // vC= -694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111110011110000; // vC= -784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111110011110011; // vC= -781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111110101011111; // vC= -673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b1111110011111110; // vC= -770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b1111110101110001; // vC= -655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b1111110101111010; // vC= -646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111110101100110; // vC= -666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b1111110110010101; // vC= -619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b1111110101100001; // vC= -671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110101010001; // vC= -687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b1111110110011010; // vC= -614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111110110101111; // vC= -593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111110101001100; // vC= -692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010011; // iC= 2067 
vC = 14'b1111110111010011; // vC= -557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000010; // iC= 2050 
vC = 14'b1111110110010011; // vC= -621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111110101111010; // vC= -646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111110110000111; // vC= -633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b1111110111110011; // vC= -525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001000; // iC= 2056 
vC = 14'b1111110101100001; // vC= -671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111110111101000; // vC= -536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111110110101011; // vC= -597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111101; // iC= 2045 
vC = 14'b1111110110000100; // vC= -636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111111000010000; // vC= -496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111111000010111; // vC= -489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b1111110110010011; // vC= -621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111110111010011; // vC= -557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111110111110001; // vC= -527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101111; // iC= 2031 
vC = 14'b1111111000111011; // vC= -453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b1111110111100100; // vC= -540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011101; // iC= 2077 
vC = 14'b1111110111001111; // vC= -561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111000100101; // vC= -475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111111000100110; // vC= -474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b1111110111011001; // vC= -551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010001; // iC= 2065 
vC = 14'b1111110111101111; // vC= -529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101111; // iC= 2031 
vC = 14'b1111111000100110; // vC= -474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000111; // iC= 2055 
vC = 14'b1111110111011101; // vC= -547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111111001110010; // vC= -398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111111000110011; // vC= -461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111111001101111; // vC= -401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111111000010011; // vC= -493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111111010010110; // vC= -362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b1111111000101111; // vC= -465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111111000111001; // vC= -455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b1111111000110001; // vC= -463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111111000011001; // vC= -487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111111001101100; // vC= -404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000010; // iC= 2050 
vC = 14'b1111111000101101; // vC= -467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001010; // iC= 2058 
vC = 14'b1111111000110100; // vC= -460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b1111111011000000; // vC= -320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100111; // iC= 2087 
vC = 14'b1111111001011000; // vC= -424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100111; // iC= 2087 
vC = 14'b1111111010011110; // vC= -354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011111; // iC= 2079 
vC = 14'b1111111011001110; // vC= -306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111111010100101; // vC= -347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101111; // iC= 2031 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010110; // iC= 2070 
vC = 14'b1111111010110001; // vC= -335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000100; // iC= 2052 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100111; // iC= 2087 
vC = 14'b1111111001101001; // vC= -407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001001; // iC= 2057 
vC = 14'b1111111010010110; // vC= -362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111111011111110; // vC= -258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010011; // iC= 2067 
vC = 14'b1111111010011011; // vC= -357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111111001111111; // vC= -385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111111011001101; // vC= -307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111111100010010; // vC= -238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111111010011100; // vC= -356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b1111111100001010; // vC= -246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111111100110011; // vC= -205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111111011111001; // vC= -263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111111011011011; // vC= -293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111111011011111; // vC= -289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b1111111100011011; // vC= -229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111011100000; // vC= -288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011001; // iC= 2073 
vC = 14'b1111111011001110; // vC= -306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111111101001010; // vC= -182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111111100100101; // vC= -219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011101; // iC= 2013 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011011; // iC= 2075 
vC = 14'b1111111101110100; // vC= -140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b1111111101011000; // vC= -168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111111100101100; // vC= -212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111111100011110; // vC= -226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011000; // iC= 2072 
vC = 14'b1111111101011101; // vC= -163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111111101110001; // vC= -143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011101; // iC= 2077 
vC = 14'b1111111110001011; // vC= -117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b1111111100111010; // vC= -198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111101001100; // vC= -180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000100; // iC= 2052 
vC = 14'b1111111110100101; // vC=  -91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b1111111101011110; // vC= -162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111111101001100; // vC= -180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b1111111101111001; // vC= -135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110111; // iC= 1975 
vC = 14'b1111111101110001; // vC= -143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111111101100100; // vC= -156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b1111111101111101; // vC= -131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b1111111111110001; // vC=  -15 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b0000000000010101; // vC=   21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111111111001111; // vC=  -49 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b1111111110011011; // vC= -101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001000; // iC= 2056 
vC = 14'b1111111110100101; // vC=  -91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111111110101111; // vC=  -81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b0000000000011101; // vC=   29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111111111011111; // vC=  -33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110111; // iC= 1975 
vC = 14'b0000000000101101; // vC=   45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111111111101100; // vC=  -20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b0000000000101000; // vC=   40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000101; // iC= 2053 
vC = 14'b0000000000000001; // vC=    1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b0000000000101111; // vC=   47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b0000000001011011; // vC=   91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b0000000000110011; // vC=   51 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b0000000000011111; // vC=   31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111100; // iC= 2044 
vC = 14'b0000000001101100; // vC=  108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b0000000000001011; // vC=   11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000001; // iC= 2049 
vC = 14'b0000000001111000; // vC=  120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b0000000001010110; // vC=   86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b0000000001000101; // vC=   69 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011011; // iC= 2011 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011001; // iC= 1881 
vC = 14'b0000000010001111; // vC=  143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b0000000001110100; // vC=  116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b0000000010101110; // vC=  174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b0000000001101010; // vC=  106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000111; // iC= 1991 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b0000000011010000; // vC=  208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b0000000010011000; // vC=  152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111010; // iC= 1978 
vC = 14'b0000000011111110; // vC=  254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b0000000100000100; // vC=  260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b0000000100000111; // vC=  263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b0000000010001010; // vC=  138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b0000000010010010; // vC=  146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b0000000100101000; // vC=  296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011001; // iC= 1881 
vC = 14'b0000000010111110; // vC=  190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b0000000011110100; // vC=  244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000000; // iC= 1984 
vC = 14'b0000000100100010; // vC=  290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b0000000011100110; // vC=  230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b0000000100100011; // vC=  291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b0000000011100000; // vC=  224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b0000000100110001; // vC=  305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001111; // iC= 1871 
vC = 14'b0000000101010101; // vC=  341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110010; // iC= 1906 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b0000000100011110; // vC=  286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b0000000101011100; // vC=  348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b0000000100011111; // vC=  287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b0000000101110010; // vC=  370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000000110001011; // vC=  395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110000; // iC= 1840 
vC = 14'b0000000101111010; // vC=  378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b0000000101010101; // vC=  341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b0000000110100101; // vC=  421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b0000000100011000; // vC=  280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b0000000101010010; // vC=  338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b0000000100110110; // vC=  310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000110100100; // vC=  420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b0000000111001011; // vC=  459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b0000000101010011; // vC=  339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000000101010001; // vC=  337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110001; // iC= 1841 
vC = 14'b0000000110011110; // vC=  414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000000111101000; // vC=  488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b0000000110101111; // vC=  431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b0000000110111101; // vC=  445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b0000000101111000; // vC=  376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b0000000110101110; // vC=  430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110110; // iC= 1846 
vC = 14'b0000000110111101; // vC=  445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b0000000110011001; // vC=  409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100000; // iC= 1824 
vC = 14'b0000000110010110; // vC=  406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000000; // iC= 1856 
vC = 14'b0000000110100110; // vC=  422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b0000000110010011; // vC=  403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000000110101111; // vC=  431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011111; // iC= 1887 
vC = 14'b0000001000000010; // vC=  514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b0000001000011011; // vC=  539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b0000001000101000; // vC=  552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b0000001000101001; // vC=  553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b0000001000101000; // vC=  552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b0000000110111000; // vC=  440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b0000001000100100; // vC=  548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000111; // iC= 1799 
vC = 14'b0000001001010001; // vC=  593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b0000001000101110; // vC=  558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010001; // iC= 1809 
vC = 14'b0000001001100100; // vC=  612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b0000000111011101; // vC=  477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000010; // iC= 1858 
vC = 14'b0000000111111101; // vC=  509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b0000001000100010; // vC=  546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b0000001000111010; // vC=  570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100110; // iC= 1766 
vC = 14'b0000001001011110; // vC=  606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b0000001000011011; // vC=  539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b0000001001111101; // vC=  637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110000; // iC= 1776 
vC = 14'b0000001000100101; // vC=  549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b0000001010001001; // vC=  649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b0000001000011111; // vC=  543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b0000001010011001; // vC=  665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000101; // iC= 1733 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001011; // iC= 1867 
vC = 14'b0000001010100101; // vC=  677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000111; // iC= 1863 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000001010000011; // vC=  643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b0000001000110101; // vC=  565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110101; // iC= 1845 
vC = 14'b0000001001110110; // vC=  630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000101; // iC= 1797 
vC = 14'b0000001010001110; // vC=  654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b0000001001101010; // vC=  618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000001001011100; // vC=  604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b0000001011101010; // vC=  746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b0000001010011111; // vC=  671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b0000001001011110; // vC=  606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100111; // iC= 1703 
vC = 14'b0000001010101111; // vC=  687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b0000001011000000; // vC=  704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b0000001011010010; // vC=  722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011000; // iC= 1688 
vC = 14'b0000001011010010; // vC=  722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100010; // iC= 1698 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b0000001010111110; // vC=  702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111100; // iC= 1788 
vC = 14'b0000001011100101; // vC=  741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111100; // iC= 1788 
vC = 14'b0000001100101111; // vC=  815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b0000001011000000; // vC=  704 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000001; // iC= 1665 
vC = 14'b0000001011010101; // vC=  725 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b0000001100011001; // vC=  793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b0000001011100101; // vC=  741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011010; // iC= 1626 
vC = 14'b0000001101000010; // vC=  834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011110; // iC= 1758 
vC = 14'b0000001100101000; // vC=  808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001000; // iC= 1736 
vC = 14'b0000001011010100; // vC=  724 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011001; // iC= 1689 
vC = 14'b0000001011011110; // vC=  734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001011; // iC= 1675 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010000; // iC= 1680 
vC = 14'b0000001011111000; // vC=  760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010100; // iC= 1748 
vC = 14'b0000001101100111; // vC=  871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010000; // iC= 1616 
vC = 14'b0000001100010111; // vC=  791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111010; // iC= 1658 
vC = 14'b0000001100101100; // vC=  812 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110110; // iC= 1590 
vC = 14'b0000001011110010; // vC=  754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b0000001101011110; // vC=  862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110110; // iC= 1654 
vC = 14'b0000001101100111; // vC=  871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011110; // iC= 1630 
vC = 14'b0000001101100111; // vC=  871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010010; // iC= 1682 
vC = 14'b0000001100110000; // vC=  816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011110; // iC= 1566 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b0000001110001001; // vC=  905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111001; // iC= 1657 
vC = 14'b0000001100111100; // vC=  828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010001; // iC= 1681 
vC = 14'b0000001110101001; // vC=  937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000110; // iC= 1670 
vC = 14'b0000001101101001; // vC=  873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b0000001101111110; // vC=  894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b0000001110111100; // vC=  956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110001; // iC= 1585 
vC = 14'b0000001110110100; // vC=  948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100000; // iC= 1632 
vC = 14'b0000001100111000; // vC=  824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b0000001101011001; // vC=  857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000100; // iC= 1540 
vC = 14'b0000001110011111; // vC=  927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000111; // iC= 1543 
vC = 14'b0000001111010101; // vC=  981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100100; // iC= 1572 
vC = 14'b0000001111000001; // vC=  961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010000; // iC= 1616 
vC = 14'b0000001111110001; // vC= 1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001000; // iC= 1608 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111001; // iC= 1529 
vC = 14'b0000001111000000; // vC=  960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b0000001110110000; // vC=  944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110101; // iC= 1589 
vC = 14'b0000001110001110; // vC=  910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001010; // iC= 1610 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b0000010000000110; // vC= 1030 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000001101111010; // vC=  890 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010010; // iC= 1618 
vC = 14'b0000001111101011; // vC= 1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100110; // iC= 1638 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000011; // iC= 1603 
vC = 14'b0000010000010000; // vC= 1040 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000101; // iC= 1605 
vC = 14'b0000001111111010; // vC= 1018 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000100; // iC= 1604 
vC = 14'b0000001111001001; // vC=  969 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010110; // iC= 1494 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011001; // iC= 1561 
vC = 14'b0000010000010110; // vC= 1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001111; // iC= 1615 
vC = 14'b0000001111101110; // vC= 1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111010; // iC= 1530 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011000; // iC= 1496 
vC = 14'b0000010000111111; // vC= 1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000110; // iC= 1542 
vC = 14'b0000010001000111; // vC= 1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101011; // iC= 1451 
vC = 14'b0000010000010110; // vC= 1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001111; // iC= 1551 
vC = 14'b0000010001010010; // vC= 1106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001100; // iC= 1484 
vC = 14'b0000001111010111; // vC=  983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010101; // iC= 1429 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000000; // iC= 1472 
vC = 14'b0000010000001111; // vC= 1039 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110111; // iC= 1463 
vC = 14'b0000010000001100; // vC= 1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001000; // iC= 1416 
vC = 14'b0000010001000111; // vC= 1095 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111010; // iC= 1530 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010100; // iC= 1428 
vC = 14'b0000010000011001; // vC= 1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001101; // iC= 1421 
vC = 14'b0000010001110010; // vC= 1138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001001; // iC= 1545 
vC = 14'b0000010000010101; // vC= 1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100011; // iC= 1507 
vC = 14'b0000010001110111; // vC= 1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100000; // iC= 1504 
vC = 14'b0000010000100011; // vC= 1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001000; // iC= 1480 
vC = 14'b0000010010001011; // vC= 1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000100; // iC= 1412 
vC = 14'b0000010000111100; // vC= 1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011111; // iC= 1375 
vC = 14'b0000010000101100; // vC= 1068 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011000; // iC= 1496 
vC = 14'b0000010001010100; // vC= 1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011111; // iC= 1503 
vC = 14'b0000010001100101; // vC= 1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100010; // iC= 1378 
vC = 14'b0000010001101011; // vC= 1131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001111; // iC= 1423 
vC = 14'b0000010001100001; // vC= 1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110101; // iC= 1461 
vC = 14'b0000010000101000; // vC= 1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000001; // iC= 1409 
vC = 14'b0000010010010011; // vC= 1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011010; // iC= 1434 
vC = 14'b0000010000110110; // vC= 1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111011; // iC= 1467 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100010; // iC= 1442 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101000; // iC= 1320 
vC = 14'b0000010010101100; // vC= 1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011100; // iC= 1436 
vC = 14'b0000010010110001; // vC= 1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001111; // iC= 1359 
vC = 14'b0000010011010101; // vC= 1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011000; // iC= 1432 
vC = 14'b0000010010101101; // vC= 1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b0000010001011110; // vC= 1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011100; // iC= 1372 
vC = 14'b0000010010100111; // vC= 1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001110; // iC= 1358 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010010; // iC= 1298 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010011; // iC= 1299 
vC = 14'b0000010010100010; // vC= 1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001101; // iC= 1357 
vC = 14'b0000010001111010; // vC= 1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000001; // iC= 1345 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010001; // iC= 1297 
vC = 14'b0000010011001111; // vC= 1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000001; // iC= 1281 
vC = 14'b0000010010101111; // vC= 1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111000; // iC= 1272 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101110; // iC= 1326 
vC = 14'b0000010011101110; // vC= 1262 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010110; // iC= 1302 
vC = 14'b0000010011101100; // vC= 1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111010; // iC= 1274 
vC = 14'b0000010010111111; // vC= 1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011110; // iC= 1246 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010100; // iC= 1300 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100100; // iC= 1316 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001111; // iC= 1295 
vC = 14'b0000010100010111; // vC= 1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100011; // iC= 1379 
vC = 14'b0000010011101100; // vC= 1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101100; // iC= 1260 
vC = 14'b0000010010100111; // vC= 1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101000; // iC= 1320 
vC = 14'b0000010011010111; // vC= 1239 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010101; // iC= 1237 
vC = 14'b0000010100111010; // vC= 1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001010; // iC= 1354 
vC = 14'b0000010100010111; // vC= 1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110100; // iC= 1268 
vC = 14'b0000010100110011; // vC= 1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010001; // iC= 1233 
vC = 14'b0000010011001001; // vC= 1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000111; // iC= 1223 
vC = 14'b0000010011110100; // vC= 1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101001; // iC= 1257 
vC = 14'b0000010100100011; // vC= 1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011000; // iC= 1304 
vC = 14'b0000010011110101; // vC= 1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011010; // iC= 1306 
vC = 14'b0000010100100011; // vC= 1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101111; // iC= 1263 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110111; // iC= 1207 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100110; // iC= 1254 
vC = 14'b0000010101000100; // vC= 1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111100; // iC= 1276 
vC = 14'b0000010101011100; // vC= 1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010110; // iC= 1302 
vC = 14'b0000010011001011; // vC= 1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000011; // iC= 1283 
vC = 14'b0000010011110000; // vC= 1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010001; // iC= 1169 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110010; // iC= 1202 
vC = 14'b0000010011110110; // vC= 1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100000; // iC= 1248 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110000; // iC= 1264 
vC = 14'b0000010101001100; // vC= 1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001001; // iC= 1225 
vC = 14'b0000010101011111; // vC= 1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011111; // iC= 1119 
vC = 14'b0000010101010000; // vC= 1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100011; // iC= 1123 
vC = 14'b0000010011100101; // vC= 1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101010; // iC= 1258 
vC = 14'b0000010011101010; // vC= 1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101001; // iC= 1129 
vC = 14'b0000010100001111; // vC= 1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011111; // iC= 1183 
vC = 14'b0000010100000110; // vC= 1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001110; // iC= 1230 
vC = 14'b0000010100011001; // vC= 1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110111; // iC= 1207 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111101; // iC= 1149 
vC = 14'b0000010101010110; // vC= 1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000100; // iC= 1156 
vC = 14'b0000010110001010; // vC= 1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010011; // iC= 1171 
vC = 14'b0000010101001011; // vC= 1355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100011; // iC= 1059 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110001; // iC= 1201 
vC = 14'b0000010101110111; // vC= 1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001001; // iC= 1161 
vC = 14'b0000010100100011; // vC= 1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000001; // iC= 1153 
vC = 14'b0000010101111111; // vC= 1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100001; // iC= 1057 
vC = 14'b0000010101010101; // vC= 1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011100; // iC= 1180 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001011; // iC= 1099 
vC = 14'b0000010101001000; // vC= 1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100100; // iC= 1124 
vC = 14'b0000010110001110; // vC= 1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111111; // iC= 1023 
vC = 14'b0000010101101101; // vC= 1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111010; // iC= 1146 
vC = 14'b0000010110001101; // vC= 1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000100; // iC= 1092 
vC = 14'b0000010110011010; // vC= 1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000100; // iC= 1092 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100101; // iC= 1061 
vC = 14'b0000010110000110; // vC= 1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101011; // iC= 1131 
vC = 14'b0000010101111010; // vC= 1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011000; // iC= 1112 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111101; // iC= 1021 
vC = 14'b0000010110010011; // vC= 1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111011; // iC= 1083 
vC = 14'b0000010101100001; // vC= 1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111101; // iC= 1085 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110000; // iC= 1008 
vC = 14'b0000010111100001; // vC= 1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100000; // iC=  992 
vC = 14'b0000010110001110; // vC= 1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000010; // iC= 1026 
vC = 14'b0000010110001111; // vC= 1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010100; // iC=  980 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010010; // iC=  978 
vC = 14'b0000010111000000; // vC= 1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101001; // iC= 1001 
vC = 14'b0000010101100111; // vC= 1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010110; // iC=  982 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101001; // iC= 1001 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010111; // iC=  983 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100110; // iC=  998 
vC = 14'b0000010110110100; // vC= 1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100000; // iC= 1056 
vC = 14'b0000010111011110; // vC= 1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001100; // iC=  972 
vC = 14'b0000010111111001; // vC= 1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b0000010110101010; // vC= 1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001101; // iC=  909 
vC = 14'b0000010111000100; // vC= 1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001000; // iC=  904 
vC = 14'b0000010110110011; // vC= 1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000001; // iC=  897 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000000; // iC=  960 
vC = 14'b0000010111001101; // vC= 1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110011; // iC= 1011 
vC = 14'b0000010110011000; // vC= 1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011110; // iC=  862 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011001; // iC=  985 
vC = 14'b0000010110011111; // vC= 1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010011; // iC=  979 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010101; // iC=  981 
vC = 14'b0000011000010111; // vC= 1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101011; // iC=  875 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000011; // iC=  963 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010001; // iC=  849 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101110; // iC=  878 
vC = 14'b0000010111011001; // vC= 1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010111; // iC=  919 
vC = 14'b0000010111010011; // vC= 1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110010; // iC=  946 
vC = 14'b0000010111101001; // vC= 1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001101; // iC=  845 
vC = 14'b0000011000101100; // vC= 1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101111; // iC=  815 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101101; // iC=  813 
vC = 14'b0000010110111010; // vC= 1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101001; // iC=  937 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011110; // iC=  862 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100111; // iC=  807 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111001; // iC=  889 
vC = 14'b0000011001000010; // vC= 1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101010; // iC=  874 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001001; // iC=  905 
vC = 14'b0000010111001010; // vC= 1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110101; // iC=  885 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000110; // iC=  838 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010100; // iC=  788 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110111; // iC=  887 
vC = 14'b0000010111001000; // vC= 1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000100; // iC=  772 
vC = 14'b0000011000001101; // vC= 1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100010; // iC=  866 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111111; // iC=  767 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000011; // iC=  835 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010110; // iC=  854 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100010; // iC=  866 
vC = 14'b0000010111001011; // vC= 1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110110; // iC=  758 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111001; // iC=  825 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000111; // iC=  775 
vC = 14'b0000011000010011; // vC= 1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101111; // iC=  815 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111001; // iC=  825 
vC = 14'b0000010111101100; // vC= 1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010101; // iC=  789 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b0000010111011001; // vC= 1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101000; // iC=  680 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011011; // iC=  731 
vC = 14'b0000011000110010; // vC= 1586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100100; // iC=  804 
vC = 14'b0000010111101010; // vC= 1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001011; // iC=  651 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100100; // iC=  676 
vC = 14'b0000011001110100; // vC= 1652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010100; // iC=  660 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010010; // iC=  786 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110110; // iC=  630 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001000; // iC=  712 
vC = 14'b0000010111101100; // vC= 1516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100010; // iC=  610 
vC = 14'b0000011001010101; // vC= 1621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011101; // iC=  669 
vC = 14'b0000010111100011; // vC= 1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101111; // iC=  751 
vC = 14'b0000011001000010; // vC= 1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001100; // iC=  652 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011100; // iC=  604 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111011; // iC=  699 
vC = 14'b0000011000110001; // vC= 1585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010110; // iC=  662 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001010; // iC=  714 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001100; // iC=  588 
vC = 14'b0000011000010011; // vC= 1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100011; // iC=  611 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111010; // iC=  634 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011011; // iC=  667 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000101; // iC=  581 
vC = 14'b0000011010000111; // vC= 1671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001110; // iC=  654 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100100; // iC=  548 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001010; // iC=  586 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011011; // iC=  539 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000101; // iC=  645 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000101; // iC=  517 
vC = 14'b0000011001000001; // vC= 1601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111111; // iC=  575 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011111; // iC=  543 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000111; // iC=  519 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110101; // iC=  565 
vC = 14'b0000011001101111; // vC= 1647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001100; // iC=  524 
vC = 14'b0000011001110101; // vC= 1653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101000; // iC=  488 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010100; // iC=  596 
vC = 14'b0000011001011110; // vC= 1630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110101; // iC=  565 
vC = 14'b0000011001011001; // vC= 1625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010011; // iC=  595 
vC = 14'b0000011000110110; // vC= 1590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101001; // iC=  553 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111111; // iC=  511 
vC = 14'b0000011010011110; // vC= 1694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101010; // iC=  490 
vC = 14'b0000011010010101; // vC= 1685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101000; // iC=  488 
vC = 14'b0000011001000101; // vC= 1605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011101; // iC=  541 
vC = 14'b0000011001011001; // vC= 1625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011101; // iC=  541 
vC = 14'b0000011010101011; // vC= 1707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101010; // iC=  426 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011110; // iC=  478 
vC = 14'b0000011010110101; // vC= 1717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111000; // iC=  504 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010110; // iC=  470 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010111; // iC=  407 
vC = 14'b0000011010101010; // vC= 1706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100111; // iC=  487 
vC = 14'b0000011001010010; // vC= 1618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011101; // iC=  349 
vC = 14'b0000011010110010; // vC= 1714 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100010; // iC=  418 
vC = 14'b0000011010101011; // vC= 1707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001010; // iC=  458 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000101; // iC=  325 
vC = 14'b0000011001100001; // vC= 1633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011010; // iC=  410 
vC = 14'b0000011010011100; // vC= 1692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011111; // iC=  287 
vC = 14'b0000011010100100; // vC= 1700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000111; // iC=  327 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111101; // iC=  253 
vC = 14'b0000011010101110; // vC= 1710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011111; // iC=  287 
vC = 14'b0000011010101110; // vC= 1710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000011; // iC=  259 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010111; // iC=  215 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110111; // iC=  311 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110100; // iC=  180 
vC = 14'b0000011001100011; // vC= 1635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011100110; // iC=  230 
vC = 14'b0000011010101010; // vC= 1706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010000111; // iC=  135 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011001; // iC=  153 
vC = 14'b0000011010000111; // vC= 1671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111001; // iC=  249 
vC = 14'b0000011010101101; // vC= 1709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101111; // iC=  111 
vC = 14'b0000011001100100; // vC= 1636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100110; // iC=  102 
vC = 14'b0000011010000101; // vC= 1669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001000; // iC=  200 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111110; // iC=   62 
vC = 14'b0000011010010011; // vC= 1683 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110001; // iC=   49 
vC = 14'b0000011001001010; // vC= 1610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010110000; // iC=  176 
vC = 14'b0000011010100111; // vC= 1703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001100; // iC=  140 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111101; // iC=   61 
vC = 14'b0000011001010111; // vC= 1623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011000; // iC=   24 
vC = 14'b0000011001101001; // vC= 1641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011010; // iC=   90 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001001; // iC=    9 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011111; // iC=   31 
vC = 14'b0000011001100110; // vC= 1638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000111; // iC=  -57 
vC = 14'b0000011010001111; // vC= 1679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001000; // iC=    8 
vC = 14'b0000011010100011; // vC= 1699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110010; // iC=  -14 
vC = 14'b0000011001111101; // vC= 1661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010100; // iC= -108 
vC = 14'b0000011001111010; // vC= 1658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001110; // iC=  -50 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101000; // iC= -216 
vC = 14'b0000011001111010; // vC= 1658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000101; // iC= -123 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011101; // iC= -227 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110000; // iC= -272 
vC = 14'b0000011001100011; // vC= 1635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011111; // iC= -289 
vC = 14'b0000011001100011; // vC= 1635 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110101; // iC= -267 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000101; // iC= -251 
vC = 14'b0000011010011010; // vC= 1690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001111; // iC= -369 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010100; // iC= -300 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000100; // iC= -380 
vC = 14'b0000011001111110; // vC= 1662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011101; // iC= -355 
vC = 14'b0000011010000110; // vC= 1670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011110; // iC= -418 
vC = 14'b0000011001011010; // vC= 1626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100000; // iC= -416 
vC = 14'b0000011010010100; // vC= 1684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100000; // iC= -416 
vC = 14'b0000011001101100; // vC= 1644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001110; // iC= -498 
vC = 14'b0000011000010010; // vC= 1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101110; // iC= -530 
vC = 14'b0000011001111011; // vC= 1659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100101; // iC= -411 
vC = 14'b0000011001011100; // vC= 1628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111111; // iC= -513 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001101; // iC= -499 
vC = 14'b0000011001110111; // vC= 1655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001111; // iC= -497 
vC = 14'b0000011000101011; // vC= 1579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010100; // iC= -684 
vC = 14'b0000011000111110; // vC= 1598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001110; // iC= -690 
vC = 14'b0000011000000001; // vC= 1537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100110; // iC= -602 
vC = 14'b0000010111111101; // vC= 1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111111; // iC= -641 
vC = 14'b0000010111110100; // vC= 1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010000; // iC= -688 
vC = 14'b0000010111100100; // vC= 1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101011; // iC= -661 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110111; // iC= -713 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001011; // iC= -693 
vC = 14'b0000011001010001; // vC= 1617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101100; // iC= -724 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111111; // iC= -769 
vC = 14'b0000011001101111; // vC= 1647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101110; // iC= -914 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010101; // iC= -939 
vC = 14'b0000010111001001; // vC= 1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001001; // iC= -951 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111100; // iC= -964 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110011; // iC= -909 
vC = 14'b0000010111000110; // vC= 1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010110; // iC=-1002 
vC = 14'b0000010111000000; // vC= 1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111100; // iC= -900 
vC = 14'b0000011001000101; // vC= 1605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011011; // iC= -997 
vC = 14'b0000010111111111; // vC= 1535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000100; // iC= -956 
vC = 14'b0000010111001011; // vC= 1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011011; // iC=-1061 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111011; // iC= -965 
vC = 14'b0000011000111000; // vC= 1592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101001; // iC=-1047 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011101; // iC=-1059 
vC = 14'b0000011000101010; // vC= 1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110000; // iC=-1168 
vC = 14'b0000010111101010; // vC= 1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000110; // iC=-1082 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101110; // iC=-1170 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010001; // iC=-1199 
vC = 14'b0000010110010001; // vC= 1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001001; // iC=-1143 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100001; // iC=-1119 
vC = 14'b0000010111110111; // vC= 1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000000; // iC=-1152 
vC = 14'b0000010110001111; // vC= 1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001011; // iC=-1269 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b0000010111001000; // vC= 1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110111; // iC=-1161 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011111; // iC=-1249 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100100; // iC=-1308 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000011; // iC=-1213 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110110; // iC=-1290 
vC = 14'b0000010110001111; // vC= 1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011100; // iC=-1252 
vC = 14'b0000010101110000; // vC= 1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011100; // iC=-1252 
vC = 14'b0000010101011011; // vC= 1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011110; // iC=-1314 
vC = 14'b0000010110100010; // vC= 1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000111; // iC=-1273 
vC = 14'b0000010110100101; // vC= 1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110010; // iC=-1422 
vC = 14'b0000010101111010; // vC= 1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101010; // iC=-1302 
vC = 14'b0000010110101001; // vC= 1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000111; // iC=-1337 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b0000010110001010; // vC= 1418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111110; // iC=-1474 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111001; // iC=-1415 
vC = 14'b0000010101011111; // vC= 1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b0000010101100100; // vC= 1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010000; // iC=-1392 
vC = 14'b0000010101001010; // vC= 1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000011; // iC=-1469 
vC = 14'b0000010100100111; // vC= 1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011100; // iC=-1444 
vC = 14'b0000010110001100; // vC= 1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b0000010101100000; // vC= 1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b0000010101100101; // vC= 1381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b0000010101110000; // vC= 1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b0000010100000100; // vC= 1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b0000010101101111; // vC= 1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b0000010100110001; // vC= 1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001101; // iC=-1587 
vC = 14'b0000010100111001; // vC= 1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b0000010100110011; // vC= 1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b0000010100010000; // vC= 1296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001010; // iC=-1654 
vC = 14'b0000010011000111; // vC= 1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111110; // iC=-1538 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b0000010011000011; // vC= 1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000010011011100; // vC= 1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b0000010101001010; // vC= 1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000001; // iC=-1599 
vC = 14'b0000010010110000; // vC= 1200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100100; // iC=-1628 
vC = 14'b0000010010100011; // vC= 1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b0000010010101000; // vC= 1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b0000010011000011; // vC= 1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000010010011001; // vC= 1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b0000010010101000; // vC= 1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000010010101000; // vC= 1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010000; // iC=-1648 
vC = 14'b0000010100000010; // vC= 1282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b0000010001111011; // vC= 1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011000; // iC=-1640 
vC = 14'b0000010001010111; // vC= 1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011111; // iC=-1633 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b0000010010100000; // vC= 1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000010011010010; // vC= 1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010110; // iC=-1642 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b0000010010110010; // vC= 1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000010000101111; // vC= 1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b0000010010010011; // vC= 1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111101; // iC=-1667 
vC = 14'b0000010010000010; // vC= 1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100100; // iC=-1628 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000010000000101; // vC= 1029 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000010000110101; // vC= 1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101000; // iC=-1688 
vC = 14'b0000010000110111; // vC= 1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000001111111111; // vC= 1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000010000101010; // vC= 1066 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100111; // iC=-1689 
vC = 14'b0000010001001100; // vC= 1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000001111111110; // vC= 1022 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111101; // iC=-1667 
vC = 14'b0000001111000101; // vC=  965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000010; // iC=-1662 
vC = 14'b0000001111110110; // vC= 1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101101; // iC=-1683 
vC = 14'b0000010000110111; // vC= 1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000010000111111; // vC= 1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b0000001110011001; // vC=  921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000001110110100; // vC=  948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b0000001111010110; // vC=  982 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000001110111011; // vC=  955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000001110101000; // vC=  936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b0000001111011011; // vC=  987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b0000001101101110; // vC=  878 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b0000001111010010; // vC=  978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b0000001110000010; // vC=  898 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000001101011000; // vC=  856 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001111100010; // vC=  994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000001110011011; // vC=  923 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000001110010011; // vC=  915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000001110010110; // vC=  918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000001110010001; // vC=  913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000001100110101; // vC=  821 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000001110101011; // vC=  939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b0000001110110110; // vC=  950 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000001101000111; // vC=  839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000100; // iC=-1724 
vC = 14'b0000001100100101; // vC=  805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001110011011; // vC=  923 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000001101001100; // vC=  844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b0000001110000100; // vC=  900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b0000001110000000; // vC=  896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010011; // iC=-1709 
vC = 14'b0000001100001110; // vC=  782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000001100100011; // vC=  803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110010; // iC=-1806 
vC = 14'b0000001101011100; // vC=  860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000001101100101; // vC=  869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100100; // iC=-1820 
vC = 14'b0000001100000010; // vC=  770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b0000001100100110; // vC=  806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000001100111000; // vC=  824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000001011010011; // vC=  723 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b0000001010101101; // vC=  685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000001011101011; // vC=  747 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011100; // iC=-1828 
vC = 14'b0000001011010111; // vC=  727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000001011110100; // vC=  756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101111; // iC=-1873 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111011; // iC=-1861 
vC = 14'b0000001010111010; // vC=  698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000001010100100; // vC=  676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110001; // iC=-1871 
vC = 14'b0000001011111011; // vC=  763 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001111; // iC=-1841 
vC = 14'b0000001011001101; // vC=  717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101010; // iC=-1750 
vC = 14'b0000001001101001; // vC=  617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100111; // iC=-1881 
vC = 14'b0000001011001111; // vC=  719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011111; // iC=-1889 
vC = 14'b0000001001111110; // vC=  638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000001011100110; // vC=  742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110010; // iC=-1870 
vC = 14'b0000001001101011; // vC=  619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001001101001; // vC=  617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111111; // iC=-1857 
vC = 14'b0000001010001010; // vC=  650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000001010011001; // vC=  665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000001001011111; // vC=  607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000001010110101; // vC=  693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000111; // iC=-1849 
vC = 14'b0000001001000001; // vC=  577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001011; // iC=-1845 
vC = 14'b0000001001111110; // vC=  638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b0000001001110011; // vC=  627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000001000001001; // vC=  521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001011; // iC=-1845 
vC = 14'b0000001001100101; // vC=  613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000001000111110; // vC=  574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000001001011010; // vC=  602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000000111110101; // vC=  501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000000111111101; // vC=  509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000001000011011; // vC=  539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011010; // iC=-1894 
vC = 14'b0000001000101011; // vC=  555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011110; // iC=-1890 
vC = 14'b0000001000010101; // vC=  533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010110; // iC=-1898 
vC = 14'b0000001000100001; // vC=  545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000111110100; // vC=  500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000000111001011; // vC=  459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000000111100000; // vC=  480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010101; // iC=-1899 
vC = 14'b0000000111000010; // vC=  450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001000000000; // vC=  512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000000111001001; // vC=  457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000001000010111; // vC=  535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110010; // iC=-1870 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000000110111001; // vC=  441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000000110100111; // vC=  423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000111; // iC=-1849 
vC = 14'b0000000101110110; // vC=  374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000000110011110; // vC=  414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010100; // iC=-1900 
vC = 14'b0000000111110100; // vC=  500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000000111000000; // vC=  448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000000101111111; // vC=  383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010001; // iC=-1903 
vC = 14'b0000000110110111; // vC=  439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000000110111110; // vC=  446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b0000000110001010; // vC=  394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000000100111001; // vC=  313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000110011110; // vC=  414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000000110011000; // vC=  408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b0000000110011010; // vC=  410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000000110110110; // vC=  438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111010; // iC=-1862 
vC = 14'b0000000101011100; // vC=  348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110101; // iC=-1867 
vC = 14'b0000000100001101; // vC=  269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000000101111000; // vC=  376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b0000000101001111; // vC=  335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000000100110011; // vC=  307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000000101100100; // vC=  356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000000100101000; // vC=  296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000010; // iC=-1854 
vC = 14'b0000000101101010; // vC=  362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010101; // iC=-1899 
vC = 14'b0000000101110110; // vC=  374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000000100110001; // vC=  305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000000101011011; // vC=  347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111000; // iC=-1864 
vC = 14'b0000000100000000; // vC=  256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111101; // iC=-1859 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000000100011100; // vC=  284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000000011000000; // vC=  192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011101; // iC=-1827 
vC = 14'b0000000101001011; // vC=  331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000011001010; // vC=  202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000000010011110; // vC=  158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000000100011011; // vC=  283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111011; // iC=-1797 
vC = 14'b0000000100010100; // vC=  276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101011; // iC=-1877 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b0000000010000110; // vC=  134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000011000000; // vC=  192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101000; // iC=-1880 
vC = 14'b0000000100000010; // vC=  258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100010; // iC=-1886 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b0000000011111100; // vC=  252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101001; // iC=-1879 
vC = 14'b0000000011011010; // vC=  218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000000001011101; // vC=   93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b0000000001100000; // vC=   96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111011; // iC=-1861 
vC = 14'b0000000010111000; // vC=  184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000000; // iC=-1792 
vC = 14'b0000000001101101; // vC=  109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000000001101111; // vC=  111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b0000000010110100; // vC=  180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b0000000010001101; // vC=  141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000000001101011; // vC=  107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b0000000001111001; // vC=  121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000000010001110; // vC=  142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110101; // iC=-1867 
vC = 14'b0000000001100010; // vC=   98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000000000100101; // vC=   37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000000001011101; // vC=   93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000000000100001; // vC=   33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011000; // iC=-1832 
vC = 14'b0000000000011001; // vC=   25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b0000000001000111; // vC=   71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011110; // iC=-1762 
vC = 14'b1111111111011111; // vC=  -33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b1111111110101111; // vC=  -81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001110; // iC=-1778 
vC = 14'b1111111111000011; // vC=  -61 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b1111111110111010; // vC=  -70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001110; // iC=-1842 
vC = 14'b1111111111001010; // vC=  -54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b1111111111111000; // vC=   -8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100011; // iC=-1821 
vC = 14'b1111111110000000; // vC= -128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b1111111111011011; // vC=  -37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b1111111110001011; // vC= -117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b1111111110000110; // vC= -122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b1111111111100000; // vC=  -32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b1111111101100000; // vC= -160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b1111111101100010; // vC= -158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b1111111110000000; // vC= -128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110000; // iC=-1680 
vC = 14'b1111111110100001; // vC=  -95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010110; // iC=-1706 
vC = 14'b1111111110101000; // vC=  -88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b1111111101101100; // vC= -148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b1111111111010000; // vC=  -48 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111000; // iC=-1800 
vC = 14'b1111111110000100; // vC= -124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b1111111110001000; // vC= -120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110110; // iC=-1674 
vC = 14'b1111111100111000; // vC= -200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b1111111101000011; // vC= -189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b1111111101111011; // vC= -133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b1111111101111100; // vC= -132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b1111111101010001; // vC= -175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b1111111100110000; // vC= -208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001010; // iC=-1654 
vC = 14'b1111111011111100; // vC= -260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b1111111110000010; // vC= -126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b1111111100000100; // vC= -252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100101; // iC=-1691 
vC = 14'b1111111101101101; // vC= -147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b1111111100001101; // vC= -243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b1111111100101000; // vC= -216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b1111111101001110; // vC= -178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b1111111011101010; // vC= -278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b1111111101001110; // vC= -178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b1111111100011110; // vC= -226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b1111111011011010; // vC= -294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b1111111010101010; // vC= -342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b1111111011010001; // vC= -303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b1111111011010000; // vC= -304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b1111111010011010; // vC= -358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110001; // iC=-1679 
vC = 14'b1111111100000100; // vC= -252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b1111111011010000; // vC= -304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b1111111011001101; // vC= -307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b1111111011011111; // vC= -289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b1111111011001011; // vC= -309 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111111; // iC=-1665 
vC = 14'b1111111100001100; // vC= -244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b1111111011010111; // vC= -297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b1111111001100100; // vC= -412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000001; // iC=-1663 
vC = 14'b1111111011110111; // vC= -265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b1111111010101101; // vC= -339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b1111111001101101; // vC= -403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b1111111010111011; // vC= -325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011011; // iC=-1637 
vC = 14'b1111111001100100; // vC= -412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010000; // iC=-1648 
vC = 14'b1111111010100101; // vC= -347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101001; // iC=-1623 
vC = 14'b1111111010011101; // vC= -355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b1111111000111010; // vC= -454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010000; // iC=-1584 
vC = 14'b1111111000111011; // vC= -453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b1111111000111010; // vC= -454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b1111111001111001; // vC= -391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b1111111000110011; // vC= -461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011001; // iC=-1639 
vC = 14'b1111111001010111; // vC= -425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b1111111010001100; // vC= -372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b1111111000001110; // vC= -498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b1111111010011010; // vC= -358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000010; // iC=-1598 
vC = 14'b1111111000011010; // vC= -486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b1111110111110111; // vC= -521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b1111111001110000; // vC= -400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100011; // iC=-1693 
vC = 14'b1111111000111110; // vC= -450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000011; // iC=-1661 
vC = 14'b1111111001110111; // vC= -393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000010; // iC=-1662 
vC = 14'b1111111000001011; // vC= -501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b1111110111101100; // vC= -532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b1111111001101111; // vC= -401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001110; // iC=-1650 
vC = 14'b1111110111100000; // vC= -544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b1111111001010001; // vC= -431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b1111111000001000; // vC= -504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111101; // iC=-1667 
vC = 14'b1111111000110101; // vC= -459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b1111110111110000; // vC= -528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b1111110111100111; // vC= -537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b1111110111011001; // vC= -551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010110; // iC=-1578 
vC = 14'b1111110111000011; // vC= -573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b1111110111101111; // vC= -529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111100; // iC=-1668 
vC = 14'b1111110110110111; // vC= -585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b1111110111001000; // vC= -568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101111; // iC=-1617 
vC = 14'b1111110110000010; // vC= -638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010101; // iC=-1515 
vC = 14'b1111110110011110; // vC= -610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001110; // iC=-1586 
vC = 14'b1111110111100111; // vC= -537 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000010; // iC=-1534 
vC = 14'b1111110110010101; // vC= -619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b1111110110000111; // vC= -633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b1111110101111001; // vC= -647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b1111110110100101; // vC= -603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101100; // iC=-1556 
vC = 14'b1111110110111111; // vC= -577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b1111110110001010; // vC= -630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100011; // iC=-1501 
vC = 14'b1111110101011010; // vC= -678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001110; // iC=-1586 
vC = 14'b1111110110010100; // vC= -620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100001; // iC=-1503 
vC = 14'b1111110101110110; // vC= -650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101011; // iC=-1557 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001100; // iC=-1588 
vC = 14'b1111110101100010; // vC= -670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111101; // iC=-1539 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b1111110101101100; // vC= -660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001110; // iC=-1458 
vC = 14'b1111110110101011; // vC= -597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b1111110110100010; // vC= -606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010010; // iC=-1582 
vC = 14'b1111110101100000; // vC= -672 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011001; // iC=-1447 
vC = 14'b1111110110101100; // vC= -596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010001; // iC=-1519 
vC = 14'b1111110101111001; // vC= -647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b1111110110100100; // vC= -604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011100; // iC=-1444 
vC = 14'b1111110100011000; // vC= -744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100110; // iC=-1434 
vC = 14'b1111110100011110; // vC= -738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110110; // iC=-1546 
vC = 14'b1111110100001100; // vC= -756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001101; // iC=-1523 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b1111110110000100; // vC= -636 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111000; // iC=-1416 
vC = 14'b1111110100101011; // vC= -725 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000011; // iC=-1469 
vC = 14'b1111110011011101; // vC= -803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b1111110100011100; // vC= -740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b1111110101010011; // vC= -685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011100; // iC=-1444 
vC = 14'b1111110100111110; // vC= -706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111011; // iC=-1413 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110000; // iC=-1488 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001010; // iC=-1526 
vC = 14'b1111110101000110; // vC= -698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b1111110100011111; // vC= -737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011000; // iC=-1448 
vC = 14'b1111110010111010; // vC= -838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100000; // iC=-1440 
vC = 14'b1111110100001000; // vC= -760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011110; // iC=-1378 
vC = 14'b1111110100001000; // vC= -760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110000; // iC=-1424 
vC = 14'b1111110100011001; // vC= -743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b1111110011111100; // vC= -772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101110; // iC=-1426 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111101; // iC=-1347 
vC = 14'b1111110011110011; // vC= -781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101000; // iC=-1432 
vC = 14'b1111110011100011; // vC= -797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b1111110001111011; // vC= -901 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101110; // iC=-1490 
vC = 14'b1111110010111000; // vC= -840 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011011; // iC=-1445 
vC = 14'b1111110010110111; // vC= -841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101001; // iC=-1431 
vC = 14'b1111110010011001; // vC= -871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010000; // iC=-1392 
vC = 14'b1111110011010001; // vC= -815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b1111110011011110; // vC= -802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010011; // iC=-1453 
vC = 14'b1111110010100001; // vC= -863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101001; // iC=-1367 
vC = 14'b1111110011100011; // vC= -797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110110; // iC=-1418 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100010; // iC=-1310 
vC = 14'b1111110010001010; // vC= -886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011001; // iC=-1383 
vC = 14'b1111110001101100; // vC= -916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110011; // iC=-1293 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111010; // iC=-1414 
vC = 14'b1111110010100000; // vC= -864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b1111110010011111; // vC= -865 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111001; // iC=-1351 
vC = 14'b1111110010010001; // vC= -879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001000; // iC=-1400 
vC = 14'b1111110010111100; // vC= -836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110000; // iC=-1296 
vC = 14'b1111110001111010; // vC= -902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001111; // iC=-1329 
vC = 14'b1111110010110010; // vC= -846 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111101; // iC=-1283 
vC = 14'b1111110001101101; // vC= -915 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110111; // iC=-1289 
vC = 14'b1111110010011101; // vC= -867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111110001000110; // vC= -954 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011001; // iC=-1319 
vC = 14'b1111110001000111; // vC= -953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010010; // iC=-1326 
vC = 14'b1111110010011100; // vC= -868 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011100; // iC=-1316 
vC = 14'b1111110001100110; // vC= -922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110101; // iC=-1291 
vC = 14'b1111110000100100; // vC= -988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101111; // iC=-1297 
vC = 14'b1111110000001010; // vC=-1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110100; // iC=-1292 
vC = 14'b1111110001110000; // vC= -912 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101111; // iC=-1361 
vC = 14'b1111110001100110; // vC= -922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100001; // iC=-1311 
vC = 14'b1111110000011110; // vC= -994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101010; // iC=-1302 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101010; // iC=-1238 
vC = 14'b1111110000011000; // vC=-1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011100; // iC=-1316 
vC = 14'b1111101111100011; // vC=-1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000010; // iC=-1278 
vC = 14'b1111110001110011; // vC= -909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100000; // iC=-1248 
vC = 14'b1111110000111110; // vC= -962 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001001; // iC=-1335 
vC = 14'b1111110000010100; // vC=-1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100111; // iC=-1241 
vC = 14'b1111110000111011; // vC= -965 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010101; // iC=-1259 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000101; // iC=-1211 
vC = 14'b1111101111010001; // vC=-1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011000; // iC=-1192 
vC = 14'b1111101111001001; // vC=-1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110101; // iC=-1227 
vC = 14'b1111110000010110; // vC=-1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111010; // iC=-1286 
vC = 14'b1111110000100011; // vC= -989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010011; // iC=-1325 
vC = 14'b1111101111100011; // vC=-1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111011; // iC=-1221 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011010; // iC=-1190 
vC = 14'b1111101110101001; // vC=-1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001011; // iC=-1205 
vC = 14'b1111110000010101; // vC=-1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b1111110000011110; // vC= -994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101110; // iC=-1298 
vC = 14'b1111101111011100; // vC=-1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010100; // iC=-1260 
vC = 14'b1111101110110111; // vC=-1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001011; // iC=-1269 
vC = 14'b1111110000011011; // vC= -997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001101; // iC=-1139 
vC = 14'b1111101110100100; // vC=-1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000011; // iC=-1149 
vC = 14'b1111101110101111; // vC=-1105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000010; // iC=-1150 
vC = 14'b1111110000100000; // vC= -992 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110000; // iC=-1232 
vC = 14'b1111110000011110; // vC= -994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100010; // iC=-1182 
vC = 14'b1111101110010111; // vC=-1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100111; // iC=-1177 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111001; // iC=-1223 
vC = 14'b1111101111101010; // vC=-1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100111; // iC=-1177 
vC = 14'b1111101111110011; // vC=-1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101110; // iC=-1234 
vC = 14'b1111101111001010; // vC=-1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101011; // iC=-1173 
vC = 14'b1111101110010010; // vC=-1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111000; // iC=-1096 
vC = 14'b1111101111010010; // vC=-1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010000; // iC=-1136 
vC = 14'b1111101111110101; // vC=-1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111001; // iC=-1095 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011001; // iC=-1127 
vC = 14'b1111101111000000; // vC=-1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001101; // iC=-1075 
vC = 14'b1111101111001010; // vC=-1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011101; // iC=-1059 
vC = 14'b1111101101110001; // vC=-1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110111; // iC=-1097 
vC = 14'b1111101101010011; // vC=-1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011111; // iC=-1121 
vC = 14'b1111101101011100; // vC=-1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111111; // iC=-1153 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110001; // iC=-1167 
vC = 14'b1111101101001000; // vC=-1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011110; // iC=-1186 
vC = 14'b1111101110010010; // vC=-1134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010110; // iC=-1130 
vC = 14'b1111101110101011; // vC=-1109 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011111; // iC=-1121 
vC = 14'b1111101101000100; // vC=-1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111101; // iC=-1091 
vC = 14'b1111101101110010; // vC=-1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101110; // iC=-1170 
vC = 14'b1111101101010110; // vC=-1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110100110; // iC=-1114 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111001; // iC=-1159 
vC = 14'b1111101100111111; // vC=-1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100100; // iC=-1052 
vC = 14'b1111101101101001; // vC=-1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111111; // iC=-1089 
vC = 14'b1111101110100100; // vC=-1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100000; // iC= -992 
vC = 14'b1111101110100101; // vC=-1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010101; // iC=-1003 
vC = 14'b1111101110000001; // vC=-1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110110; // iC=-1034 
vC = 14'b1111101101010111; // vC=-1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111000; // iC=-1096 
vC = 14'b1111101110011011; // vC=-1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011000; // iC=-1128 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001110; // iC=-1074 
vC = 14'b1111101100100001; // vC=-1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111010; // iC=-1094 
vC = 14'b1111101101110011; // vC=-1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101111; // iC=-1105 
vC = 14'b1111101101101000; // vC=-1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110001; // iC=-1039 
vC = 14'b1111101011111110; // vC=-1282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010010; // iC=-1006 
vC = 14'b1111101101101010; // vC=-1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100100; // iC= -988 
vC = 14'b1111101110000110; // vC=-1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110011; // iC= -973 
vC = 14'b1111101110010000; // vC=-1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001110; // iC= -946 
vC = 14'b1111101100110101; // vC=-1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001001; // iC= -951 
vC = 14'b1111101011111010; // vC=-1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111101101001001; // vC=-1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111101100111011; // vC=-1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111010; // iC= -966 
vC = 14'b1111101100010001; // vC=-1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110011; // iC= -973 
vC = 14'b1111101101110011; // vC=-1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101001; // iC=-1047 
vC = 14'b1111101100011000; // vC=-1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100011; // iC= -989 
vC = 14'b1111101100001001; // vC=-1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b1111101100001111; // vC=-1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001110; // iC=-1010 
vC = 14'b1111101101010111; // vC=-1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110111; // iC= -905 
vC = 14'b1111101011111100; // vC=-1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101010; // iC= -982 
vC = 14'b1111101100001110; // vC=-1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000111; // iC=-1017 
vC = 14'b1111101101100101; // vC=-1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110111; // iC= -905 
vC = 14'b1111101101010100; // vC=-1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000100; // iC= -892 
vC = 14'b1111101100110101; // vC=-1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100001; // iC= -927 
vC = 14'b1111101100011001; // vC=-1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110001; // iC= -911 
vC = 14'b1111101100010011; // vC=-1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111001; // iC= -967 
vC = 14'b1111101011010111; // vC=-1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001100; // iC= -948 
vC = 14'b1111101100110011; // vC=-1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011100; // iC= -868 
vC = 14'b1111101100010011; // vC=-1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001010; // iC= -886 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000000; // iC= -896 
vC = 14'b1111101010110101; // vC=-1355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010111; // iC= -937 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010100; // iC= -876 
vC = 14'b1111101100010101; // vC=-1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000111; // iC= -953 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111100; // iC= -836 
vC = 14'b1111101011111000; // vC=-1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000001; // iC= -895 
vC = 14'b1111101100010100; // vC=-1260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010110; // iC= -938 
vC = 14'b1111101100101110; // vC=-1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110010; // iC= -910 
vC = 14'b1111101011011001; // vC=-1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010001; // iC= -815 
vC = 14'b1111101100101110; // vC=-1234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000111; // iC= -825 
vC = 14'b1111101010001000; // vC=-1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110110; // iC= -906 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011000; // iC= -808 
vC = 14'b1111101100000011; // vC=-1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000110; // iC= -826 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001001; // iC= -823 
vC = 14'b1111101011111011; // vC=-1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110000; // iC= -848 
vC = 14'b1111101011001000; // vC=-1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101001; // iC= -791 
vC = 14'b1111101100000101; // vC=-1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110000; // iC= -784 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100101; // iC= -859 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101110; // iC= -786 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010111; // iC= -809 
vC = 14'b1111101010000011; // vC=-1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010011; // iC= -813 
vC = 14'b1111101100000010; // vC=-1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100011; // iC= -861 
vC = 14'b1111101001111110; // vC=-1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110100; // iC= -780 
vC = 14'b1111101010100010; // vC=-1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101110; // iC= -850 
vC = 14'b1111101011101000; // vC=-1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101111; // iC= -721 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000100; // iC= -828 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110110; // iC= -778 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001001; // iC= -695 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111000; // iC= -712 
vC = 14'b1111101010101100; // vC=-1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011011; // iC= -805 
vC = 14'b1111101001100111; // vC=-1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110110; // iC= -714 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001011; // iC= -693 
vC = 14'b1111101011011110; // vC=-1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001011; // iC= -693 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100100; // iC= -796 
vC = 14'b1111101010000110; // vC=-1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100000; // iC= -672 
vC = 14'b1111101010001001; // vC=-1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000000; // iC= -640 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111000; // iC= -776 
vC = 14'b1111101010100001; // vC=-1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001001; // iC= -631 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100000; // iC= -736 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001110; // iC= -690 
vC = 14'b1111101010001111; // vC=-1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011100; // iC= -740 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001101; // iC= -691 
vC = 14'b1111101010000110; // vC=-1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100100; // iC= -604 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111100; // iC= -644 
vC = 14'b1111101010100010; // vC=-1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101011; // iC= -597 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110101; // iC= -651 
vC = 14'b1111101010010111; // vC=-1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011001; // iC= -679 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111101; // iC= -579 
vC = 14'b1111101001000000; // vC=-1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010000; // iC= -688 
vC = 14'b1111101010011010; // vC=-1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001101; // iC= -627 
vC = 14'b1111101010000111; // vC=-1401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110111; // iC= -585 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000110; // iC= -634 
vC = 14'b1111101010101010; // vC=-1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010001; // iC= -559 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100111; // iC= -665 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101011; // iC= -661 
vC = 14'b1111101010010100; // vC=-1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000000; // iC= -512 
vC = 14'b1111101000100000; // vC=-1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001011; // iC= -501 
vC = 14'b1111101000010011; // vC=-1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110011; // iC= -525 
vC = 14'b1111101001100111; // vC=-1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001110; // iC= -562 
vC = 14'b1111101010010001; // vC=-1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001100; // iC= -500 
vC = 14'b1111101001001000; // vC=-1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111111; // iC= -577 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011000; // iC= -552 
vC = 14'b1111101010100100; // vC=-1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b1111101000010111; // vC=-1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111101000100111; // vC=-1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110110; // iC= -458 
vC = 14'b1111101000001100; // vC=-1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011100; // iC= -548 
vC = 14'b1111101000100010; // vC=-1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110011; // iC= -589 
vC = 14'b1111101010011100; // vC=-1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100100; // iC= -540 
vC = 14'b1111101000011110; // vC=-1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001011; // iC= -565 
vC = 14'b1111101000110011; // vC=-1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111001101; // iC= -563 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010100; // iC= -492 
vC = 14'b1111101000100001; // vC=-1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101010; // iC= -470 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110000; // iC= -464 
vC = 14'b1111101001100110; // vC=-1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000011; // iC= -509 
vC = 14'b1111100111111010; // vC=-1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011110; // iC= -546 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100101; // iC= -539 
vC = 14'b1111101001101001; // vC=-1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100111; // iC= -409 
vC = 14'b1111101000100111; // vC=-1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010001; // iC= -367 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110101; // iC= -459 
vC = 14'b1111100111101110; // vC=-1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101001; // iC= -471 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100010; // iC= -478 
vC = 14'b1111101000100101; // vC=-1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100001; // iC= -351 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010010; // iC= -430 
vC = 14'b1111101000010000; // vC=-1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011001; // iC= -423 
vC = 14'b1111101000011001; // vC=-1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100001; // iC= -351 
vC = 14'b1111101000011000; // vC=-1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011101100; // iC= -276 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000011; // iC= -253 
vC = 14'b1111101000100010; // vC=-1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010101; // iC= -299 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001010; // iC= -374 
vC = 14'b1111101000111100; // vC=-1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011011101; // iC= -291 
vC = 14'b1111101000101100; // vC=-1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111110; // iC= -322 
vC = 14'b1111101000000010; // vC=-1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010110; // iC= -298 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100100; // iC= -284 
vC = 14'b1111101001010100; // vC=-1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100011; // iC= -285 
vC = 14'b1111101001101101; // vC=-1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101000; // iC= -216 
vC = 14'b1111100111110001; // vC=-1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100110100; // iC= -204 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101011; // iC= -213 
vC = 14'b1111100111111100; // vC=-1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011100; // iC= -164 
vC = 14'b1111101000000000; // vC=-1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010100; // iC= -172 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011111; // iC=  -97 
vC = 14'b1111101000100100; // vC=-1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111100; // iC= -196 
vC = 14'b1111100111110110; // vC=-1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000100; // iC= -124 
vC = 14'b1111100111010011; // vC=-1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011100; // iC= -164 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001110; // iC= -114 
vC = 14'b1111101001001111; // vC=-1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011010; // iC= -102 
vC = 14'b1111101000011101; // vC=-1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111110011; // iC=  -13 
vC = 14'b1111101000110011; // vC=-1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110101101; // iC=  -83 
vC = 14'b1111101001001001; // vC=-1463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011100; // iC=   28 
vC = 14'b1111101001000011; // vC=-1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111001; // iC=   -7 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000101; // iC=   69 
vC = 14'b1111101001110000; // vC=-1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100101; // iC=  101 
vC = 14'b1111100111100000; // vC=-1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101000; // iC=  104 
vC = 14'b1111101001010000; // vC=-1456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010100111; // iC=  167 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101001; // iC=  105 
vC = 14'b1111101000001001; // vC=-1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001010; // iC=  202 
vC = 14'b1111101000100100; // vC=-1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111110; // iC=  126 
vC = 14'b1111101000010010; // vC=-1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000010; // iC=  194 
vC = 14'b1111101000111111; // vC=-1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000111; // iC=  199 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000111; // iC=  263 
vC = 14'b1111100111101000; // vC=-1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001011; // iC=  203 
vC = 14'b1111100111011011; // vC=-1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010010; // iC=  338 
vC = 14'b1111100111110000; // vC=-1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111101; // iC=  317 
vC = 14'b1111100111110100; // vC=-1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010101; // iC=  277 
vC = 14'b1111101000110000; // vC=-1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110111; // iC=  375 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111111; // iC=  447 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111101; // iC=  381 
vC = 14'b1111101000110101; // vC=-1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011001; // iC=  473 
vC = 14'b1111100111101101; // vC=-1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011101; // iC=  413 
vC = 14'b1111101001110000; // vC=-1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011111; // iC=  479 
vC = 14'b1111101000111001; // vC=-1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101001; // iC=  425 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101000; // iC=  552 
vC = 14'b1111101001000001; // vC=-1471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110001; // iC=  497 
vC = 14'b1111101000001101; // vC=-1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001011; // iC=  523 
vC = 14'b1111100111111001; // vC=-1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100000; // iC=  672 
vC = 14'b1111101000001101; // vC=-1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111010; // iC=  634 
vC = 14'b1111101000000111; // vC=-1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011011; // iC=  603 
vC = 14'b1111100111110010; // vC=-1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000110; // iC=  710 
vC = 14'b1111101001101010; // vC=-1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011111; // iC=  735 
vC = 14'b1111101000001101; // vC=-1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001110; // iC=  654 
vC = 14'b1111101010010101; // vC=-1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000101; // iC=  773 
vC = 14'b1111101001011000; // vC=-1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001011; // iC=  779 
vC = 14'b1111101001111000; // vC=-1416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001110; // iC=  718 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000000; // iC=  832 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110100; // iC=  756 
vC = 14'b1111101000001000; // vC=-1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000100; // iC=  900 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110110; // iC=  886 
vC = 14'b1111101010100001; // vC=-1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101101; // iC=  941 
vC = 14'b1111101001101010; // vC=-1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111110; // iC=  894 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010100; // iC=  916 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001111; // iC= 1039 
vC = 14'b1111101000111100; // vC=-1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100100; // iC=  932 
vC = 14'b1111101001100100; // vC=-1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011011; // iC= 1051 
vC = 14'b1111101001111011; // vC=-1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001100; // iC= 1036 
vC = 14'b1111101010101100; // vC=-1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111011; // iC= 1083 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b1111101010101001; // vC=-1367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110001; // iC= 1009 
vC = 14'b1111101000110001; // vC=-1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010101; // iC= 1173 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001000; // iC= 1160 
vC = 14'b1111101011001011; // vC=-1333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010110; // iC= 1174 
vC = 14'b1111101001101000; // vC=-1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100101; // iC= 1189 
vC = 14'b1111101001110010; // vC=-1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110001; // iC= 1201 
vC = 14'b1111101010000100; // vC=-1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110111; // iC= 1271 
vC = 14'b1111101001110101; // vC=-1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001111; // iC= 1167 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110010; // iC= 1202 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110011; // iC= 1203 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110100; // iC= 1268 
vC = 14'b1111101001100001; // vC=-1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000000; // iC= 1280 
vC = 14'b1111101011111000; // vC=-1288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010111; // iC= 1303 
vC = 14'b1111101001101101; // vC=-1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111001; // iC= 1273 
vC = 14'b1111101011001010; // vC=-1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001001; // iC= 1417 
vC = 14'b1111101001101110; // vC=-1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100000; // iC= 1312 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100000; // iC= 1312 
vC = 14'b1111101011010101; // vC=-1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101111; // iC= 1391 
vC = 14'b1111101010000101; // vC=-1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001001; // iC= 1481 
vC = 14'b1111101100000110; // vC=-1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010101; // iC= 1493 
vC = 14'b1111101010101110; // vC=-1362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111100; // iC= 1532 
vC = 14'b1111101010110100; // vC=-1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010111; // iC= 1495 
vC = 14'b1111101011000101; // vC=-1339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001011; // iC= 1419 
vC = 14'b1111101011100110; // vC=-1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010101; // iC= 1429 
vC = 14'b1111101100101011; // vC=-1237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110100; // iC= 1460 
vC = 14'b1111101011101001; // vC=-1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000101; // iC= 1477 
vC = 14'b1111101010101010; // vC=-1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000110; // iC= 1542 
vC = 14'b1111101010110110; // vC=-1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010011; // iC= 1619 
vC = 14'b1111101011100110; // vC=-1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010101; // iC= 1621 
vC = 14'b1111101100111001; // vC=-1223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011000; // iC= 1560 
vC = 14'b1111101011011000; // vC=-1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010100; // iC= 1556 
vC = 14'b1111101100000011; // vC=-1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010111; // iC= 1623 
vC = 14'b1111101100111110; // vC=-1218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101011; // iC= 1643 
vC = 14'b1111101011101000; // vC=-1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000000; // iC= 1600 
vC = 14'b1111101101010100; // vC=-1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100000; // iC= 1568 
vC = 14'b1111101101111001; // vC=-1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110100; // iC= 1716 
vC = 14'b1111101011110011; // vC=-1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000100; // iC= 1732 
vC = 14'b1111101100010011; // vC=-1261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b1111101101111001; // vC=-1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011001; // iC= 1625 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011000; // iC= 1752 
vC = 14'b1111101110010111; // vC=-1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100110; // iC= 1702 
vC = 14'b1111101101111000; // vC=-1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100011; // iC= 1699 
vC = 14'b1111101101000011; // vC=-1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001100; // iC= 1676 
vC = 14'b1111101100101010; // vC=-1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001111; // iC= 1679 
vC = 14'b1111101101010010; // vC=-1198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101010; // iC= 1834 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b1111101110010001; // vC=-1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001010; // iC= 1738 
vC = 14'b1111101100110110; // vC=-1226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100101; // iC= 1765 
vC = 14'b1111101110110101; // vC=-1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110010; // iC= 1778 
vC = 14'b1111101110110101; // vC=-1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010111; // iC= 1751 
vC = 14'b1111101111000011; // vC=-1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000000; // iC= 1792 
vC = 14'b1111101110000011; // vC=-1149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100110; // iC= 1766 
vC = 14'b1111101110011010; // vC=-1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b1111101111000011; // vC=-1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101110; // iC= 1838 
vC = 14'b1111101110100010; // vC=-1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b1111101111011011; // vC=-1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b1111101110000000; // vC=-1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b1111101101110011; // vC=-1165 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010111; // iC= 1815 
vC = 14'b1111101110011010; // vC=-1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000000; // iC= 1792 
vC = 14'b1111101110110111; // vC=-1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111101111101111; // vC=-1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101110; // iC= 1838 
vC = 14'b1111101110010001; // vC=-1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111110000000001; // vC=-1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b1111101111111110; // vC=-1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100110; // iC= 1830 
vC = 14'b1111110000000000; // vC=-1024 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111101111111110; // vC=-1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b1111101111110101; // vC=-1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b1111110000010101; // vC=-1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b1111110001001101; // vC= -947 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b1111110000000111; // vC=-1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b1111110001010100; // vC= -940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111110001011100; // vC= -932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110001000000; // vC= -960 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b1111110000010000; // vC=-1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b1111101111111100; // vC=-1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001011; // iC= 1867 
vC = 14'b1111110001000011; // vC= -957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b1111110010001001; // vC= -887 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110000111110; // vC= -962 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111110001010111; // vC= -937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111110001110100; // vC= -908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b1111110011000110; // vC= -826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b1111110001001111; // vC= -945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b1111110011001100; // vC= -820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111110001111101; // vC= -899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111110010100010; // vC= -862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111110011001001; // vC= -823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111110010000100; // vC= -892 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111110011110111; // vC= -777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111110100110100; // vC= -716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b1111110010011001; // vC= -871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111110100111001; // vC= -711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111110011110110; // vC= -778 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111110100110100; // vC= -716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b1111110100100000; // vC= -736 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101010; // iC= 1898 
vC = 14'b1111110011001001; // vC= -823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b1111110100000010; // vC= -766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110100100010; // vC= -734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111110011100100; // vC= -796 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111110011110101; // vC= -779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b1111110101110110; // vC= -650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010100; // iC= 2004 
vC = 14'b1111110101001000; // vC= -696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111110110001001; // vC= -631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111110101011001; // vC= -679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b1111110110001101; // vC= -627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111110101111100; // vC= -644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010110; // iC= 2070 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110100011001; // vC= -743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111110100011010; // vC= -742 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b1111110101011100; // vC= -676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111110110001010; // vC= -630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111110101110110; // vC= -650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001001; // iC= 2057 
vC = 14'b1111110110010110; // vC= -618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110111; // iC= 1975 
vC = 14'b1111110111011001; // vC= -551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111110110111010; // vC= -582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111110110100110; // vC= -602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001001; // iC= 2057 
vC = 14'b1111110110100101; // vC= -603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010011; // iC= 2067 
vC = 14'b1111110111001111; // vC= -561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111110110010010; // vC= -622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111110111101100; // vC= -532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111110101110101; // vC= -651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001001; // iC= 2057 
vC = 14'b1111110110001000; // vC= -632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111110111011111; // vC= -545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011010; // iC= 2074 
vC = 14'b1111110110001001; // vC= -631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111110111001110; // vC= -562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111110110111001; // vC= -583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001110; // iC= 2062 
vC = 14'b1111111000000111; // vC= -505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010101; // iC= 1941 
vC = 14'b1111110111001100; // vC= -564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110111; // iC= 2039 
vC = 14'b1111111000100011; // vC= -477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000111; // iC= 1991 
vC = 14'b1111110110111010; // vC= -582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010001; // iC= 2065 
vC = 14'b1111111001001100; // vC= -436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b1111111001010010; // vC= -430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111000010101; // vC= -491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b1111110111100011; // vC= -541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111000; // iC= 1976 
vC = 14'b1111111000111001; // vC= -455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111111001001011; // vC= -437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001101; // iC= 2061 
vC = 14'b1111111001001001; // vC= -439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111111000100011; // vC= -477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001110; // iC= 2062 
vC = 14'b1111111001010011; // vC= -429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000000; // iC= 1984 
vC = 14'b1111111000001001; // vC= -503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111111000110010; // vC= -462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111111000101111; // vC= -465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011110; // iC= 2078 
vC = 14'b1111111001111010; // vC= -390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111111001101010; // vC= -406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111111001011111; // vC= -417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111010011000; // vC= -360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100110; // iC= 2086 
vC = 14'b1111111001110101; // vC= -395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010101; // iC= 2069 
vC = 14'b1111111001000010; // vC= -446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b1111111001110001; // vC= -399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001101; // iC= 2061 
vC = 14'b1111111001111110; // vC= -386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000000; // iC= 2048 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100111; // iC= 2023 
vC = 14'b1111111011101010; // vC= -278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011101; // iC= 2077 
vC = 14'b1111111001111000; // vC= -392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111111010010001; // vC= -367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111111010100011; // vC= -349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b1111111100010000; // vC= -240 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010100; // iC= 2068 
vC = 14'b1111111010010101; // vC= -363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b1111111100101010; // vC= -214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101101; // iC= 2029 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b1111111010011111; // vC= -353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111111100000010; // vC= -254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110010; // iC= 2034 
vC = 14'b1111111010110111; // vC= -329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b1111111011110111; // vC= -265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111111100001101; // vC= -243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b1111111101001011; // vC= -181 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011110; // iC= 2078 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010010; // iC= 2066 
vC = 14'b1111111101100000; // vC= -160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000111; // iC= 2055 
vC = 14'b1111111100111101; // vC= -195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111111101100110; // vC= -154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111111101100101; // vC= -155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000001; // iC= 2049 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111011111100; // vC= -260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b1111111101111101; // vC= -131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b1111111101100110; // vC= -154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111111100111110; // vC= -194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b1111111101111110; // vC= -130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100101; // iC= 2021 
vC = 14'b1111111100101101; // vC= -211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111111100110111; // vC= -201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b1111111100101100; // vC= -212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010010; // iC= 2066 
vC = 14'b1111111100110110; // vC= -202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111111101111011; // vC= -133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111111110011101; // vC=  -99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111001; // iC= 2041 
vC = 14'b1111111100111111; // vC= -193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011001; // iC= 2073 
vC = 14'b1111111101110110; // vC= -138 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b1111111111010111; // vC=  -41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b1111111110101110; // vC=  -82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111111110110011; // vC=  -77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111111110000010; // vC= -126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111100; // iC= 2044 
vC = 14'b1111111110001011; // vC= -117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b0000000000000110; // vC=    6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111111101000; // vC=  -24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001101; // iC= 2061 
vC = 14'b0000000000000101; // vC=    5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b0000000000010101; // vC=   21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b1111111110100110; // vC=  -90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b0000000000000100; // vC=    4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b0000000000010011; // vC=   19 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111111111100011; // vC=  -29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b0000000000101100; // vC=   44 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111111110100110; // vC=  -90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111111111101111; // vC=  -17 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110011; // iC= 2035 
vC = 14'b1111111111010101; // vC=  -43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b0000000001011000; // vC=   88 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000111; // iC= 2055 
vC = 14'b1111111111111000; // vC=   -8 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b0000000000101011; // vC=   43 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b0000000001001111; // vC=   79 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111111111010111; // vC=  -41 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111111111110101; // vC=  -11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100101; // iC= 2021 
vC = 14'b0000000000000110; // vC=    6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b0000000001010010; // vC=   82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b0000000001010110; // vC=   86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b0000000001001101; // vC=   77 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b0000000000011001; // vC=   25 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000000000100110; // vC=   38 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b0000000010000000; // vC=  128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b0000000010101101; // vC=  173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b0000000001111101; // vC=  125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b0000000010010101; // vC=  149 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b0000000010100110; // vC=  166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b0000000010101100; // vC=  172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b0000000010100011; // vC=  163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b0000000010100110; // vC=  166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b0000000001100111; // vC=  103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b0000000011110110; // vC=  246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b0000000001100001; // vC=   97 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b0000000010000010; // vC=  130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b0000000011100100; // vC=  228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b0000000100000101; // vC=  261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011011; // iC= 2011 
vC = 14'b0000000100001100; // vC=  268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b0000000011011000; // vC=  216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000100011101; // vC=  285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b0000000100001000; // vC=  264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b0000000100010101; // vC=  277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b0000000010110111; // vC=  183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b0000000100000111; // vC=  263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000011; // iC= 1987 
vC = 14'b0000000100111100; // vC=  316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b0000000100000011; // vC=  259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010001; // iC= 1873 
vC = 14'b0000000101010101; // vC=  341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110101; // iC= 1845 
vC = 14'b0000000100100111; // vC=  295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b0000000011111010; // vC=  250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111001; // iC= 1849 
vC = 14'b0000000101010010; // vC=  338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b0000000101011100; // vC=  348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110010; // iC= 1970 
vC = 14'b0000000100010000; // vC=  272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101100; // iC= 1964 
vC = 14'b0000000100100101; // vC=  293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101100; // iC= 1964 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b0000000101010011; // vC=  339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b0000000100101101; // vC=  301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001110; // iC= 1870 
vC = 14'b0000000101100100; // vC=  356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b0000000101111001; // vC=  377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b0000000110100111; // vC=  423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b0000000101000000; // vC=  320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b0000000100011101; // vC=  285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b0000000100110011; // vC=  307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101010; // iC= 1898 
vC = 14'b0000000110110011; // vC=  435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b0000000100111010; // vC=  314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b0000000110111010; // vC=  442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b0000000101001011; // vC=  331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001100; // iC= 1804 
vC = 14'b0000000110000000; // vC=  384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101010; // iC= 1898 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111011; // iC= 1851 
vC = 14'b0000000101111011; // vC=  379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b0000000111011001; // vC=  473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b0000000110011100; // vC=  412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000011; // iC= 1795 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011111; // iC= 1823 
vC = 14'b0000000111111100; // vC=  508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b0000000110100000; // vC=  416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b0000000111101101; // vC=  493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b0000000111000101; // vC=  453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b0000000111100101; // vC=  485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b0000001000101001; // vC=  553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001000; // iC= 1864 
vC = 14'b0000000111100011; // vC=  483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b0000000110111011; // vC=  443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b0000001000110111; // vC=  567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110101; // iC= 1909 
vC = 14'b0000000110110111; // vC=  439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110010; // iC= 1906 
vC = 14'b0000001000111100; // vC=  572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100011; // iC= 1763 
vC = 14'b0000000111011011; // vC=  475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b0000000110111001; // vC=  441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b0000001001001100; // vC=  588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b0000000111010110; // vC=  470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001100; // iC= 1804 
vC = 14'b0000000111011110; // vC=  478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b0000000111111010; // vC=  506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010101; // iC= 1749 
vC = 14'b0000001000100001; // vC=  545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010110; // iC= 1814 
vC = 14'b0000000111011010; // vC=  474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b0000001000011111; // vC=  543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b0000001000011110; // vC=  542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b0000001000011010; // vC=  538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110001; // iC= 1777 
vC = 14'b0000001010001100; // vC=  652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111111; // iC= 1727 
vC = 14'b0000001001110101; // vC=  629 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000100; // iC= 1796 
vC = 14'b0000001001000010; // vC=  578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111110; // iC= 1726 
vC = 14'b0000001000011111; // vC=  543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110101; // iC= 1845 
vC = 14'b0000001010101000; // vC=  680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011000; // iC= 1816 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b0000001001101010; // vC=  618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110000; // iC= 1840 
vC = 14'b0000001001110011; // vC=  627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000011; // iC= 1859 
vC = 14'b0000001001100010; // vC=  610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110111; // iC= 1847 
vC = 14'b0000001001001110; // vC=  590 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111000; // iC= 1720 
vC = 14'b0000001010011111; // vC=  671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100010; // iC= 1762 
vC = 14'b0000001001101111; // vC=  623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100010; // iC= 1698 
vC = 14'b0000001010011000; // vC=  664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b0000001001010010; // vC=  594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b0000001010001010; // vC=  650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010111; // iC= 1751 
vC = 14'b0000001011000010; // vC=  706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b0000001011010010; // vC=  722 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001110; // iC= 1742 
vC = 14'b0000001010110111; // vC=  695 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000100; // iC= 1668 
vC = 14'b0000001010100010; // vC=  674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110110; // iC= 1782 
vC = 14'b0000001100000101; // vC=  773 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110011; // iC= 1715 
vC = 14'b0000001100001100; // vC=  780 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b0000001010111001; // vC=  697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100110; // iC= 1702 
vC = 14'b0000001011110000; // vC=  752 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111100; // iC= 1724 
vC = 14'b0000001011010111; // vC=  727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000000; // iC= 1664 
vC = 14'b0000001100000100; // vC=  772 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000001011110010; // vC=  754 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000101; // iC= 1669 
vC = 14'b0000001011101111; // vC=  751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110110; // iC= 1654 
vC = 14'b0000001011011100; // vC=  732 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001110; // iC= 1742 
vC = 14'b0000001100011100; // vC=  796 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101000; // iC= 1768 
vC = 14'b0000001010100101; // vC=  677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111000; // iC= 1656 
vC = 14'b0000001100011001; // vC=  793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010011; // iC= 1683 
vC = 14'b0000001011001100; // vC=  716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b0000001011000111; // vC=  711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010010; // iC= 1746 
vC = 14'b0000001011001101; // vC=  717 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001010; // iC= 1610 
vC = 14'b0000001011111101; // vC=  765 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b0000001011001011; // vC=  715 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110100; // iC= 1716 
vC = 14'b0000001011100001; // vC=  737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000001100010000; // vC=  784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001100; // iC= 1612 
vC = 14'b0000001101101101; // vC=  877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110000; // iC= 1648 
vC = 14'b0000001101101101; // vC=  877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000001100110110; // vC=  822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b0000001110000111; // vC=  903 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111110; // iC= 1598 
vC = 14'b0000001110001011; // vC=  907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011110; // iC= 1630 
vC = 14'b0000001101111111; // vC=  895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100101; // iC= 1573 
vC = 14'b0000001100010001; // vC=  785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010011; // iC= 1619 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101011; // iC= 1579 
vC = 14'b0000001101111110; // vC=  894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101010; // iC= 1578 
vC = 14'b0000001110010001; // vC=  913 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111010; // iC= 1594 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111110; // iC= 1662 
vC = 14'b0000001100101001; // vC=  809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111010; // iC= 1658 
vC = 14'b0000001110010111; // vC=  919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010100; // iC= 1684 
vC = 14'b0000001101000000; // vC=  832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100000; // iC= 1696 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111101; // iC= 1533 
vC = 14'b0000001101000101; // vC=  837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110111; // iC= 1655 
vC = 14'b0000001101010000; // vC=  848 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111100; // iC= 1596 
vC = 14'b0000001111000100; // vC=  964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001000; // iC= 1608 
vC = 14'b0000001101000101; // vC=  837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001100; // iC= 1548 
vC = 14'b0000001111010010; // vC=  978 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100111; // iC= 1575 
vC = 14'b0000001101100101; // vC=  869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100111; // iC= 1639 
vC = 14'b0000001110101110; // vC=  942 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011011; // iC= 1627 
vC = 14'b0000001101101001; // vC=  873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010110; // iC= 1622 
vC = 14'b0000001101011011; // vC=  859 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000001; // iC= 1601 
vC = 14'b0000001111100010; // vC=  994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110000; // iC= 1520 
vC = 14'b0000001110101010; // vC=  938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110110; // iC= 1526 
vC = 14'b0000001110000011; // vC=  899 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101000; // iC= 1512 
vC = 14'b0000001110011010; // vC=  922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101000; // iC= 1640 
vC = 14'b0000001111101000; // vC= 1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111111; // iC= 1599 
vC = 14'b0000001101111000; // vC=  888 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011110; // iC= 1566 
vC = 14'b0000001111101100; // vC= 1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001100; // iC= 1612 
vC = 14'b0000001111111101; // vC= 1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010000; // iC= 1552 
vC = 14'b0000001111011110; // vC=  990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111000; // iC= 1464 
vC = 14'b0000001110110010; // vC=  946 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b0000001110111101; // vC=  957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111111; // iC= 1471 
vC = 14'b0000010000000010; // vC= 1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110110; // iC= 1590 
vC = 14'b0000010000110101; // vC= 1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000101; // iC= 1477 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110001; // iC= 1457 
vC = 14'b0000010000011010; // vC= 1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111001; // iC= 1593 
vC = 14'b0000001110100011; // vC=  931 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101111; // iC= 1519 
vC = 14'b0000010000110111; // vC= 1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000000; // iC= 1472 
vC = 14'b0000001111101111; // vC= 1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011110; // iC= 1566 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001101; // iC= 1549 
vC = 14'b0000001111100011; // vC=  995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010001; // iC= 1489 
vC = 14'b0000010000111100; // vC= 1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011100; // iC= 1500 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010101; // iC= 1493 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100110; // iC= 1510 
vC = 14'b0000010001001001; // vC= 1097 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001111; // iC= 1423 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110010; // iC= 1458 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000000; // iC= 1408 
vC = 14'b0000010001110000; // vC= 1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011000; // iC= 1496 
vC = 14'b0000010000110111; // vC= 1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111111; // iC= 1535 
vC = 14'b0000010000110000; // vC= 1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100111; // iC= 1511 
vC = 14'b0000010000010010; // vC= 1042 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110000; // iC= 1392 
vC = 14'b0000010000111101; // vC= 1085 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010011; // iC= 1427 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011001; // iC= 1433 
vC = 14'b0000010000001001; // vC= 1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011010; // iC= 1498 
vC = 14'b0000010001101001; // vC= 1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010010; // iC= 1490 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111010; // iC= 1466 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000001; // iC= 1345 
vC = 14'b0000010001110111; // vC= 1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110110; // iC= 1462 
vC = 14'b0000010010010111; // vC= 1175 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001001; // iC= 1481 
vC = 14'b0000010000110100; // vC= 1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010010; // iC= 1490 
vC = 14'b0000010001111010; // vC= 1146 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001110; // iC= 1486 
vC = 14'b0000010001101101; // vC= 1133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011010; // iC= 1370 
vC = 14'b0000010010001111; // vC= 1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101110; // iC= 1326 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110010; // iC= 1458 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000111; // iC= 1351 
vC = 14'b0000010001101101; // vC= 1133 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111001; // iC= 1401 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000110; // iC= 1350 
vC = 14'b0000010001010100; // vC= 1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110100; // iC= 1332 
vC = 14'b0000010010010000; // vC= 1168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100100; // iC= 1380 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000111; // iC= 1287 
vC = 14'b0000010010110101; // vC= 1205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111001; // iC= 1401 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011000; // iC= 1304 
vC = 14'b0000010001001110; // vC= 1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001101; // iC= 1357 
vC = 14'b0000010010001000; // vC= 1160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001010; // iC= 1354 
vC = 14'b0000010001110111; // vC= 1143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110110; // iC= 1270 
vC = 14'b0000010010001110; // vC= 1166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011100; // iC= 1372 
vC = 14'b0000010011001001; // vC= 1225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100111; // iC= 1383 
vC = 14'b0000010011100101; // vC= 1253 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000000; // iC= 1280 
vC = 14'b0000010100000011; // vC= 1283 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100001; // iC= 1313 
vC = 14'b0000010011111010; // vC= 1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010101; // iC= 1365 
vC = 14'b0000010100000101; // vC= 1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001111; // iC= 1359 
vC = 14'b0000010011010011; // vC= 1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101101; // iC= 1389 
vC = 14'b0000010011000110; // vC= 1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000111; // iC= 1223 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110011; // iC= 1331 
vC = 14'b0000010011011111; // vC= 1247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010100; // iC= 1236 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110100; // iC= 1268 
vC = 14'b0000010100001010; // vC= 1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010100; // iC= 1300 
vC = 14'b0000010010100100; // vC= 1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100001; // iC= 1249 
vC = 14'b0000010100010011; // vC= 1299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101101; // iC= 1325 
vC = 14'b0000010100010111; // vC= 1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110010; // iC= 1330 
vC = 14'b0000010011110001; // vC= 1265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011110; // iC= 1246 
vC = 14'b0000010100100111; // vC= 1319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110101; // iC= 1333 
vC = 14'b0000010100110111; // vC= 1335 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000100; // iC= 1220 
vC = 14'b0000010100000110; // vC= 1286 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000111; // iC= 1223 
vC = 14'b0000010100101011; // vC= 1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000010011110100; // vC= 1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001110; // iC= 1166 
vC = 14'b0000010010111111; // vC= 1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100100; // iC= 1316 
vC = 14'b0000010010101111; // vC= 1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111100; // iC= 1212 
vC = 14'b0000010100101111; // vC= 1327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101011; // iC= 1195 
vC = 14'b0000010100111011; // vC= 1339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100110; // iC= 1254 
vC = 14'b0000010100111011; // vC= 1339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100100; // iC= 1252 
vC = 14'b0000010101000101; // vC= 1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100000; // iC= 1248 
vC = 14'b0000010011101000; // vC= 1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000010011010110; // vC= 1238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101000; // iC= 1256 
vC = 14'b0000010101011000; // vC= 1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100100; // iC= 1124 
vC = 14'b0000010100111010; // vC= 1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110000; // iC= 1136 
vC = 14'b0000010011001111; // vC= 1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111101; // iC= 1213 
vC = 14'b0000010101000001; // vC= 1345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101101; // iC= 1197 
vC = 14'b0000010100111101; // vC= 1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101100; // iC= 1196 
vC = 14'b0000010100110001; // vC= 1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000010; // iC= 1154 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001011111; // iC= 1119 
vC = 14'b0000010100011000; // vC= 1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010100; // iC= 1236 
vC = 14'b0000010101001110; // vC= 1358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000010011111001; // vC= 1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010000001; // iC= 1153 
vC = 14'b0000010110001011; // vC= 1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000110; // iC= 1094 
vC = 14'b0000010101111111; // vC= 1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001100; // iC= 1164 
vC = 14'b0000010101011111; // vC= 1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110011; // iC= 1203 
vC = 14'b0000010101000100; // vC= 1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010110100; // iC= 1204 
vC = 14'b0000010100110010; // vC= 1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101011; // iC= 1195 
vC = 14'b0000010110001011; // vC= 1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100001; // iC= 1185 
vC = 14'b0000010101011001; // vC= 1369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011111; // iC= 1183 
vC = 14'b0000010101100000; // vC= 1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000000; // iC= 1088 
vC = 14'b0000010110011111; // vC= 1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010000; // iC= 1040 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011101; // iC= 1053 
vC = 14'b0000010110000101; // vC= 1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000100; // iC= 1028 
vC = 14'b0000010101010100; // vC= 1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111100; // iC= 1148 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111110; // iC= 1022 
vC = 14'b0000010101000011; // vC= 1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110000; // iC= 1072 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010100; // iC= 1044 
vC = 14'b0000010101101100; // vC= 1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110011; // iC= 1075 
vC = 14'b0000010101010011; // vC= 1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100000; // iC= 1120 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111111010; // iC= 1018 
vC = 14'b0000010101010011; // vC= 1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100000; // iC=  992 
vC = 14'b0000010100101100; // vC= 1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010101; // iC=  981 
vC = 14'b0000010110010011; // vC= 1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100101; // iC= 1061 
vC = 14'b0000010111001101; // vC= 1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010010; // iC= 1106 
vC = 14'b0000010101101111; // vC= 1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011110; // iC=  990 
vC = 14'b0000010110110001; // vC= 1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011000; // iC= 1048 
vC = 14'b0000010101101000; // vC= 1384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110100; // iC= 1076 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011011; // iC= 1051 
vC = 14'b0000010110010001; // vC= 1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011110; // iC= 1054 
vC = 14'b0000010101110011; // vC= 1395 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000110000; // iC= 1072 
vC = 14'b0000010110100110; // vC= 1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011011; // iC=  923 
vC = 14'b0000010110010100; // vC= 1428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011100; // iC=  924 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011000; // iC=  984 
vC = 14'b0000010110000001; // vC= 1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000000; // iC=  960 
vC = 14'b0000010101110001; // vC= 1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010001; // iC= 1041 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001011; // iC=  907 
vC = 14'b0000010101111101; // vC= 1405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000100; // iC=  900 
vC = 14'b0000010111001111; // vC= 1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000000; // iC=  960 
vC = 14'b0000010110001011; // vC= 1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011001; // iC=  985 
vC = 14'b0000010101101011; // vC= 1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010110; // iC=  918 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111000; // iC=  952 
vC = 14'b0000010111100111; // vC= 1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011000; // iC=  920 
vC = 14'b0000010111100110; // vC= 1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011111; // iC=  927 
vC = 14'b0000010110000001; // vC= 1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110011; // iC=  947 
vC = 14'b0000010110010111; // vC= 1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110000; // iC=  880 
vC = 14'b0000010111000001; // vC= 1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101101; // iC=  877 
vC = 14'b0000010110110100; // vC= 1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010101; // iC=  917 
vC = 14'b0000010111011000; // vC= 1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011100; // iC=  860 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001111; // iC=  847 
vC = 14'b0000010110110110; // vC= 1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111000011; // iC=  963 
vC = 14'b0000010110001100; // vC= 1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001001; // iC=  905 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010010; // iC=  914 
vC = 14'b0000010110010111; // vC= 1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111100; // iC=  892 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111001; // iC=  825 
vC = 14'b0000010110010110; // vC= 1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001111; // iC=  911 
vC = 14'b0000010111000101; // vC= 1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110001; // iC=  817 
vC = 14'b0000010111010111; // vC= 1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100110100; // iC=  820 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011000; // iC=  856 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010110; // iC=  918 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010100; // iC=  852 
vC = 14'b0000010110011100; // vC= 1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001111; // iC=  783 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011111; // iC=  799 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110110; // iC=  886 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000111; // iC=  839 
vC = 14'b0000010111111001; // vC= 1529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110011; // iC=  755 
vC = 14'b0000011000010111; // vC= 1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101111; // iC=  815 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101001; // iC=  873 
vC = 14'b0000010111111101; // vC= 1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101001011; // iC=  843 
vC = 14'b0000010111000010; // vC= 1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000100; // iC=  772 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000001; // iC=  833 
vC = 14'b0000010110111001; // vC= 1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110111; // iC=  695 
vC = 14'b0000011001001101; // vC= 1613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011011; // iC=  731 
vC = 14'b0000010111011100; // vC= 1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010110; // iC=  726 
vC = 14'b0000011001000010; // vC= 1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000110; // iC=  710 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011100; // iC=  796 
vC = 14'b0000011000111110; // vC= 1598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010011; // iC=  723 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111001; // iC=  761 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111100; // iC=  700 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111010; // iC=  698 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100111; // iC=  679 
vC = 14'b0000010111001000; // vC= 1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000110; // iC=  646 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000111; // iC=  711 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010101000; // iC=  680 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111110; // iC=  766 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001000; // iC=  648 
vC = 14'b0000010111111110; // vC= 1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101010; // iC=  618 
vC = 14'b0000010111111011; // vC= 1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100010; // iC=  674 
vC = 14'b0000011001101000; // vC= 1640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010000; // iC=  656 
vC = 14'b0000010111111011; // vC= 1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110001; // iC=  689 
vC = 14'b0000010111010100; // vC= 1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001000; // iC=  712 
vC = 14'b0000011001101100; // vC= 1644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010011; // iC=  659 
vC = 14'b0000010111011110; // vC= 1502 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011000; // iC=  664 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111110; // iC=  574 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110011; // iC=  691 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010111110; // iC=  702 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011110; // iC=  670 
vC = 14'b0000011001010101; // vC= 1621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101101; // iC=  621 
vC = 14'b0000011001110110; // vC= 1654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001110000; // iC=  624 
vC = 14'b0000010111100010; // vC= 1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010011001; // iC=  665 
vC = 14'b0000011001101101; // vC= 1645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100110; // iC=  614 
vC = 14'b0000011001010010; // vC= 1618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001011; // iC=  587 
vC = 14'b0000011001110000; // vC= 1648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000010; // iC=  642 
vC = 14'b0000011001101000; // vC= 1640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101001; // iC=  553 
vC = 14'b0000011001110011; // vC= 1651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010101; // iC=  597 
vC = 14'b0000011000110001; // vC= 1585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000000; // iC=  576 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000110; // iC=  518 
vC = 14'b0000011010001010; // vC= 1674 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010101; // iC=  597 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010010; // iC=  594 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011010; // iC=  602 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000000000; // iC=  512 
vC = 14'b0000011010001011; // vC= 1675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101100; // iC=  492 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111000; // iC=  504 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001010000; // iC=  592 
vC = 14'b0000011000001110; // vC= 1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001100; // iC=  460 
vC = 14'b0000011010001101; // vC= 1677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001100; // iC=  588 
vC = 14'b0000011000010110; // vC= 1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111110011; // iC=  499 
vC = 14'b0000011000101100; // vC= 1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100100; // iC=  548 
vC = 14'b0000011001111010; // vC= 1658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000000; // iC=  576 
vC = 14'b0000011001000110; // vC= 1606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101100; // iC=  556 
vC = 14'b0000011010010101; // vC= 1685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100100; // iC=  420 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011111; // iC=  415 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100110; // iC=  422 
vC = 14'b0000011001010101; // vC= 1621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010110; // iC=  470 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011010; // iC=  474 
vC = 14'b0000011001100010; // vC= 1634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100110; // iC=  358 
vC = 14'b0000011010100101; // vC= 1701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111000010; // iC=  450 
vC = 14'b0000011000110100; // vC= 1588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011100; // iC=  412 
vC = 14'b0000011000011011; // vC= 1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100110; // iC=  422 
vC = 14'b0000011001110101; // vC= 1653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100000; // iC=  352 
vC = 14'b0000011001001101; // vC= 1613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100110001; // iC=  305 
vC = 14'b0000011010000111; // vC= 1671 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110100100; // iC=  420 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101101100; // iC=  364 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100001001; // iC=  265 
vC = 14'b0000011010100001; // vC= 1697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100000; // iC=  352 
vC = 14'b0000011010010111; // vC= 1687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001101; // iC=  333 
vC = 14'b0000011001110110; // vC= 1654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111011; // iC=  251 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011001101; // iC=  205 
vC = 14'b0000011010001101; // vC= 1677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010110; // iC=  278 
vC = 14'b0000011001111011; // vC= 1659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000111; // iC=  263 
vC = 14'b0000011001011000; // vC= 1624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000111; // iC=  263 
vC = 14'b0000011001111111; // vC= 1663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111011; // iC=  251 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100101; // iC=  293 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001001; // iC=  137 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000011; // iC=  195 
vC = 14'b0000011000010111; // vC= 1559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000001; // iC=  193 
vC = 14'b0000011000111110; // vC= 1598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010011000; // iC=  152 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001010000; // iC=   80 
vC = 14'b0000011001100101; // vC= 1637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000010; // iC=   66 
vC = 14'b0000011010010111; // vC= 1687 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101010; // iC=   42 
vC = 14'b0000011010000000; // vC= 1664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011011; // iC=   27 
vC = 14'b0000011001010111; // vC= 1623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101101; // iC=  109 
vC = 14'b0000011010000000; // vC= 1664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001000011; // iC=   67 
vC = 14'b0000011000100110; // vC= 1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000000; // iC=    0 
vC = 14'b0000011001101111; // vC= 1647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001100011; // iC=   99 
vC = 14'b0000011001100110; // vC= 1638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011010; // iC=   26 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001110; // iC=   14 
vC = 14'b0000011000101101; // vC= 1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011101; // iC=   29 
vC = 14'b0000011010011100; // vC= 1692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110010111; // iC= -105 
vC = 14'b0000011010000011; // vC= 1667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111001; // iC=   -7 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101011000; // iC= -168 
vC = 14'b0000011000111110; // vC= 1598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111000; // iC= -136 
vC = 14'b0000011000111111; // vC= 1599 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101101; // iC= -147 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101110; // iC= -146 
vC = 14'b0000011001010100; // vC= 1620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001111; // iC= -241 
vC = 14'b0000011001010100; // vC= 1620 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100001; // iC= -159 
vC = 14'b0000011000101111; // vC= 1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001101; // iC= -307 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111000; // iC= -200 
vC = 14'b0000011000100000; // vC= 1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001000; // iC= -248 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111011; // iC= -261 
vC = 14'b0000011010001110; // vC= 1678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101110; // iC= -338 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010011010; // iC= -358 
vC = 14'b0000011001001000; // vC= 1608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111011; // iC= -389 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000101; // iC= -443 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100011; // iC= -413 
vC = 14'b0000011001101000; // vC= 1640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101011; // iC= -469 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110111; // iC= -521 
vC = 14'b0000011001101100; // vC= 1644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000000; // iC= -512 
vC = 14'b0000010111110011; // vC= 1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111111110; // iC= -514 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101001; // iC= -535 
vC = 14'b0000011001110101; // vC= 1653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011000; // iC= -616 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111000; // iC= -584 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110010; // iC= -590 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101100; // iC= -596 
vC = 14'b0000011000110011; // vC= 1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100010; // iC= -670 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011111; // iC= -609 
vC = 14'b0000011000110010; // vC= 1586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101000; // iC= -728 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010111; // iC= -809 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100000; // iC= -736 
vC = 14'b0000011000111001; // vC= 1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100000; // iC= -736 
vC = 14'b0000011000111000; // vC= 1592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101010; // iC= -726 
vC = 14'b0000011000101111; // vC= 1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100100; // iC= -860 
vC = 14'b0000011000110111; // vC= 1591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000000; // iC= -768 
vC = 14'b0000011000100111; // vC= 1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001111; // iC= -817 
vC = 14'b0000011001000001; // vC= 1601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110000; // iC= -848 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110110; // iC= -906 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010000; // iC= -944 
vC = 14'b0000010111100001; // vC= 1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010110; // iC= -874 
vC = 14'b0000010111001010; // vC= 1482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000011; // iC= -957 
vC = 14'b0000011000111100; // vC= 1596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010011; // iC=-1005 
vC = 14'b0000010111010100; // vC= 1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101111; // iC= -977 
vC = 14'b0000010111100011; // vC= 1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010001; // iC= -943 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000000; // iC=-1024 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111110; // iC=-1090 
vC = 14'b0000011000100011; // vC= 1571 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110111; // iC=-1033 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001010; // iC=-1142 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010010; // iC=-1134 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101001; // iC=-1111 
vC = 14'b0000010110111110; // vC= 1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110001; // iC=-1167 
vC = 14'b0000010111010111; // vC= 1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111010; // iC=-1222 
vC = 14'b0000010110101101; // vC= 1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110010; // iC=-1230 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101101; // iC=-1107 
vC = 14'b0000010111101111; // vC= 1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001111; // iC=-1265 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b0000010101110100; // vC= 1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111011; // iC=-1285 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100000; // iC=-1184 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000101; // iC=-1275 
vC = 14'b0000010101101110; // vC= 1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111010; // iC=-1350 
vC = 14'b0000010101111100; // vC= 1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010110; // iC=-1258 
vC = 14'b0000010110010011; // vC= 1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b0000010110010000; // vC= 1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110001; // iC=-1359 
vC = 14'b0000010110011100; // vC= 1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100101; // iC=-1307 
vC = 14'b0000010110010110; // vC= 1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110101; // iC=-1419 
vC = 14'b0000010100111111; // vC= 1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001010; // iC=-1398 
vC = 14'b0000010110110011; // vC= 1459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011101; // iC=-1443 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010000; // iC=-1456 
vC = 14'b0000010101010100; // vC= 1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100011; // iC=-1437 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000100; // iC=-1404 
vC = 14'b0000010100011111; // vC= 1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000101; // iC=-1467 
vC = 14'b0000010110011010; // vC= 1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100011; // iC=-1501 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b0000010101000110; // vC= 1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b0000010100000001; // vC= 1281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010111; // iC=-1449 
vC = 14'b0000010101011101; // vC= 1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111101; // iC=-1475 
vC = 14'b0000010110001001; // vC= 1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b0000010101000110; // vC= 1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101010; // iC=-1430 
vC = 14'b0000010101010110; // vC= 1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101001; // iC=-1495 
vC = 14'b0000010101000111; // vC= 1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010101; // iC=-1451 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b0000010100010110; // vC= 1302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001100; // iC=-1460 
vC = 14'b0000010011111011; // vC= 1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100000; // iC=-1568 
vC = 14'b0000010011101011; // vC= 1259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101010; // iC=-1622 
vC = 14'b0000010100010001; // vC= 1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001001; // iC=-1591 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100001; // iC=-1567 
vC = 14'b0000010100000101; // vC= 1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101101; // iC=-1619 
vC = 14'b0000010100111111; // vC= 1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101010; // iC=-1558 
vC = 14'b0000010010110111; // vC= 1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b0000010011100111; // vC= 1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101110; // iC=-1554 
vC = 14'b0000010011100011; // vC= 1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b0000010100110000; // vC= 1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001101; // iC=-1651 
vC = 14'b0000010010101100; // vC= 1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111101; // iC=-1667 
vC = 14'b0000010010010010; // vC= 1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b0000010011101111; // vC= 1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010111; // iC=-1641 
vC = 14'b0000010100001101; // vC= 1293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b0000010010000101; // vC= 1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100000; // iC=-1632 
vC = 14'b0000010010011011; // vC= 1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110101; // iC=-1675 
vC = 14'b0000010011001000; // vC= 1224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000010010101101; // vC= 1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b0000010011110000; // vC= 1264 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000010001101100; // vC= 1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101010; // iC=-1686 
vC = 14'b0000010010111100; // vC= 1212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000010001011100; // vC= 1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000001; // iC=-1663 
vC = 14'b0000010010100100; // vC= 1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101110; // iC=-1618 
vC = 14'b0000010010110100; // vC= 1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000010001010011; // vC= 1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b0000010010000100; // vC= 1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b0000010000011001; // vC= 1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000010010000111; // vC= 1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101100; // iC=-1620 
vC = 14'b0000010000110111; // vC= 1079 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000010001111001; // vC= 1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000010000110011; // vC= 1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111000; // iC=-1736 
vC = 14'b0000010000111011; // vC= 1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000001111100110; // vC=  998 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000010001111001; // vC= 1145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000010000011110; // vC= 1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000010000001001; // vC= 1033 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111010; // iC=-1798 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000010000001000; // vC= 1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b0000001110111110; // vC=  958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111100; // iC=-1668 
vC = 14'b0000010001001111; // vC= 1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000001111101001; // vC= 1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000001111101001; // vC= 1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b0000010000101111; // vC= 1071 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000001111101011; // vC= 1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000001111101000; // vC= 1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000001110010010; // vC=  914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000001110010111; // vC=  919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b0000001111111111; // vC= 1023 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b0000001110111110; // vC=  958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000001110100111; // vC=  935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000001110110111; // vC=  951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b0000001101101000; // vC=  872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000001110011110; // vC=  926 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101101; // iC=-1811 
vC = 14'b0000001110101000; // vC=  936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000001101111011; // vC=  891 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000001110110100; // vC=  948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001110111011; // vC=  955 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100100; // iC=-1820 
vC = 14'b0000001110110111; // vC=  951 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b0000001110111000; // vC=  952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010000; // iC=-1840 
vC = 14'b0000001110101011; // vC=  939 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000001101110100; // vC=  884 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000001101011100; // vC=  860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100100; // iC=-1756 
vC = 14'b0000001101000101; // vC=  837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000001100110110; // vC=  822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001001; // iC=-1783 
vC = 14'b0000001110010100; // vC=  916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101010; // iC=-1750 
vC = 14'b0000001110010100; // vC=  916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000001100000001; // vC=  769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000001011101000; // vC=  744 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b0000001101111101; // vC=  893 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000001100110100; // vC=  820 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000001101010010; // vC=  850 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000001101000110; // vC=  838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000001100000110; // vC=  774 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111010; // iC=-1862 
vC = 14'b0000001100101110; // vC=  814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000001011101010; // vC=  746 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000001011011011; // vC=  731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101010; // iC=-1750 
vC = 14'b0000001011111000; // vC=  760 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000001100110000; // vC=  816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000001011000011; // vC=  707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b0000001011110001; // vC=  753 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000001011011011; // vC=  731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010101; // iC=-1771 
vC = 14'b0000001010110011; // vC=  691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000100; // iC=-1724 
vC = 14'b0000001001111001; // vC=  633 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000001100000111; // vC=  775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000000; // iC=-1792 
vC = 14'b0000001011011101; // vC=  733 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000001011000001; // vC=  705 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111011; // iC=-1861 
vC = 14'b0000001010001100; // vC=  652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010100; // iC=-1836 
vC = 14'b0000001001100110; // vC=  614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000001001010010; // vC=  594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100010; // iC=-1886 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000001011001001; // vC=  713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101011; // iC=-1877 
vC = 14'b0000001000101110; // vC=  558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001001110110; // vC=  630 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b0000001001000100; // vC=  580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011110; // iC=-1890 
vC = 14'b0000001010100001; // vC=  673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000001000010001; // vC=  529 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b0000001010010000; // vC=  656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b0000001001111000; // vC=  632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b0000001010001010; // vC=  650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000001000011110; // vC=  542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110110; // iC=-1866 
vC = 14'b0000000111111001; // vC=  505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001011; // iC=-1781 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000000111111110; // vC=  510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000001000110111; // vC=  567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011010; // iC=-1830 
vC = 14'b0000001001100011; // vC=  611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000001001000011; // vC=  579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101000; // iC=-1816 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011010; // iC=-1894 
vC = 14'b0000000111000100; // vC=  452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001010; // iC=-1846 
vC = 14'b0000000111010001; // vC=  465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110000; // iC=-1872 
vC = 14'b0000000110100010; // vC=  418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000000111111111; // vC=  511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000110111000; // vC=  440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000000110100100; // vC=  420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101010; // iC=-1878 
vC = 14'b0000000110001010; // vC=  394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010010; // iC=-1774 
vC = 14'b0000000111000000; // vC=  448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110000; // iC=-1872 
vC = 14'b0000000111000000; // vC=  448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000000101111010; // vC=  378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b0000000101101001; // vC=  361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011010; // iC=-1894 
vC = 14'b0000000110011101; // vC=  413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110111; // iC=-1737 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000000110110101; // vC=  437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000010; // iC=-1854 
vC = 14'b0000000101111011; // vC=  379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000110100001; // vC=  417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000000101001010; // vC=  330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b0000000110011111; // vC=  415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000000111000111; // vC=  455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000000100111100; // vC=  316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001010; // iC=-1782 
vC = 14'b0000000110000110; // vC=  390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010010101; // iC=-1899 
vC = 14'b0000000110010011; // vC=  403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000000100010110; // vC=  278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111110; // iC=-1858 
vC = 14'b0000000100010101; // vC=  277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001111; // iC=-1841 
vC = 14'b0000000110000011; // vC=  387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000000110000100; // vC=  388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000000101100110; // vC=  358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011111; // iC=-1825 
vC = 14'b0000000101011101; // vC=  349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100010; // iC=-1758 
vC = 14'b0000000110000000; // vC=  384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000000101010010; // vC=  338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000000011100011; // vC=  227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011011; // iC=-1893 
vC = 14'b0000000101101110; // vC=  366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000000101010111; // vC=  343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111011; // iC=-1861 
vC = 14'b0000000100011010; // vC=  282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b0000000101100011; // vC=  355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000011011111; // vC=  223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000000100011001; // vC=  281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b0000000011100010; // vC=  226 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100101; // iC=-1755 
vC = 14'b0000000010110011; // vC=  179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000000100011001; // vC=  281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110010; // iC=-1870 
vC = 14'b0000000011001000; // vC=  200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111111; // iC=-1857 
vC = 14'b0000000100001001; // vC=  265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000000010101000; // vC=  168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110111; // iC=-1865 
vC = 14'b0000000010010001; // vC=  145 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100000; // iC=-1824 
vC = 14'b0000000010100111; // vC=  167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000000011110001; // vC=  241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000000; // iC=-1856 
vC = 14'b0000000100010000; // vC=  272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000000011110101; // vC=  245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000000010100011; // vC=  163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110010; // iC=-1870 
vC = 14'b0000000011110011; // vC=  243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000000011011111; // vC=  223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101001; // iC=-1815 
vC = 14'b0000000010110010; // vC=  178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000000011011001; // vC=  217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b0000000010111110; // vC=  190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010101; // iC=-1835 
vC = 14'b0000000001011110; // vC=   94 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010011; // iC=-1837 
vC = 14'b0000000010000000; // vC=  128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110100; // iC=-1868 
vC = 14'b0000000000101000; // vC=   40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010111; // iC=-1833 
vC = 14'b0000000010010100; // vC=  148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000000010101011; // vC=  171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110100; // iC=-1740 
vC = 14'b0000000010000100; // vC=  132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000000001001100; // vC=   76 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110000; // iC=-1872 
vC = 14'b0000000001010000; // vC=   80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111101; // iC=-1859 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b0000000000011111; // vC=   31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111001; // iC=-1863 
vC = 14'b1111111111100110; // vC=  -26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b0000000000010011; // vC=   19 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000000001001110; // vC=   78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b1111111111001011; // vC=  -53 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001010; // iC=-1846 
vC = 14'b1111111111111001; // vC=   -7 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b1111111111001011; // vC=  -53 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001101; // iC=-1715 
vC = 14'b0000000000000110; // vC=    6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011100; // iC=-1764 
vC = 14'b1111111111000110; // vC=  -58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111110; // iC=-1730 
vC = 14'b1111111111011100; // vC=  -36 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101101; // iC=-1747 
vC = 14'b1111111110100000; // vC=  -96 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b1111111111101100; // vC=  -20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101010; // iC=-1814 
vC = 14'b1111111110111001; // vC=  -71 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b1111111111111101; // vC=   -3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b1111111111111101; // vC=   -3 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b1111111111100110; // vC=  -26 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001011; // iC=-1845 
vC = 14'b1111111111100101; // vC=  -27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b1111111110100011; // vC=  -93 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b1111111111001110; // vC=  -50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001100; // iC=-1844 
vC = 14'b1111111110011001; // vC= -103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b1111111110010100; // vC= -108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b1111111111110100; // vC=  -12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010011; // iC=-1773 
vC = 14'b1111111111100101; // vC=  -27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100000; // iC=-1760 
vC = 14'b1111111110010010; // vC= -110 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b1111111110100111; // vC=  -89 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b1111111100111100; // vC= -196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b1111111110100110; // vC=  -90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b1111111110010101; // vC= -107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010100; // iC=-1708 
vC = 14'b1111111101010100; // vC= -172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100001; // iC=-1823 
vC = 14'b1111111100100010; // vC= -222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b1111111110010110; // vC= -106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b1111111110101010; // vC=  -86 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b1111111101101101; // vC= -147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b1111111101000001; // vC= -191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b1111111100000001; // vC= -255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b1111111100100011; // vC= -221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000010; // iC=-1662 
vC = 14'b1111111100011100; // vC= -228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b1111111100110000; // vC= -208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110111; // iC=-1801 
vC = 14'b1111111011111100; // vC= -260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001101; // iC=-1651 
vC = 14'b1111111101000110; // vC= -186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000001; // iC=-1663 
vC = 14'b1111111101101000; // vC= -152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b1111111100010110; // vC= -234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b1111111011110001; // vC= -271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111001; // iC=-1799 
vC = 14'b1111111011111101; // vC= -259 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b1111111011001100; // vC= -308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b1111111100111101; // vC= -195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b1111111010101010; // vC= -342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b1111111100100110; // vC= -218 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001000; // iC=-1656 
vC = 14'b1111111011011011; // vC= -293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b1111111100001111; // vC= -241 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b1111111011011010; // vC= -294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001010; // iC=-1654 
vC = 14'b1111111100101001; // vC= -215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b1111111010100000; // vC= -352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101010; // iC=-1686 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b1111111011110011; // vC= -269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b1111111011011010; // vC= -294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b1111111100000111; // vC= -249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b1111111011001000; // vC= -312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b1111111011011010; // vC= -294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101110; // iC=-1682 
vC = 14'b1111111001010110; // vC= -426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011101; // iC=-1699 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b1111111001011101; // vC= -419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111110; // iC=-1666 
vC = 14'b1111111011011011; // vC= -293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111000; // iC=-1608 
vC = 14'b1111111010111001; // vC= -327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b1111111010001100; // vC= -372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b1111111000111011; // vC= -453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101001; // iC=-1623 
vC = 14'b1111111010101111; // vC= -337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b1111111010001110; // vC= -370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b1111111001000010; // vC= -446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b1111111000011001; // vC= -487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b1111111000100110; // vC= -474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111001; // iC=-1671 
vC = 14'b1111111001011100; // vC= -420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010100; // iC=-1580 
vC = 14'b1111111010011100; // vC= -356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111110; // iC=-1602 
vC = 14'b1111111001011010; // vC= -422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b1111111010010000; // vC= -368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011000; // iC=-1576 
vC = 14'b1111111000011111; // vC= -481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000100; // iC=-1660 
vC = 14'b1111111000111001; // vC= -455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b1111111000100000; // vC= -480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b1111111000110011; // vC= -461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b1111111000101101; // vC= -467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b1111111000000110; // vC= -506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001001; // iC=-1655 
vC = 14'b1111111001100001; // vC= -415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b1111111001010100; // vC= -428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b1111111000001000; // vC= -504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110101; // iC=-1547 
vC = 14'b1111111000011110; // vC= -482 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b1111111001000100; // vC= -444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b1111111000001011; // vC= -501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111100; // iC=-1604 
vC = 14'b1111110110101110; // vC= -594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b1111110111001111; // vC= -561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b1111111000001000; // vC= -504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000011; // iC=-1533 
vC = 14'b1111110110011111; // vC= -609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110001; // iC=-1551 
vC = 14'b1111110110111101; // vC= -579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000111; // iC=-1529 
vC = 14'b1111110111111111; // vC= -513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b1111111000011100; // vC= -484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110111; // iC=-1609 
vC = 14'b1111110110101000; // vC= -600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b1111110111110100; // vC= -524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b1111110110000001; // vC= -639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101011; // iC=-1621 
vC = 14'b1111110111011010; // vC= -550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110111; // iC=-1609 
vC = 14'b1111111000001111; // vC= -497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010101; // iC=-1643 
vC = 14'b1111110101101111; // vC= -657 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101000; // iC=-1496 
vC = 14'b1111111000000001; // vC= -511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010010; // iC=-1582 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110011; // iC=-1613 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001011; // iC=-1589 
vC = 14'b1111110101101000; // vC= -664 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b1111110111010001; // vC= -559 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011100; // iC=-1508 
vC = 14'b1111110101111100; // vC= -644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b1111110101010100; // vC= -684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b1111110111000110; // vC= -570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111011; // iC=-1477 
vC = 14'b1111110101100010; // vC= -670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b1111110110101111; // vC= -593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111101; // iC=-1475 
vC = 14'b1111110110100000; // vC= -608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001100; // iC=-1524 
vC = 14'b1111110100111111; // vC= -705 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110001; // iC=-1551 
vC = 14'b1111110110010001; // vC= -623 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011010; // iC=-1510 
vC = 14'b1111110101110111; // vC= -649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011101; // iC=-1507 
vC = 14'b1111110110000010; // vC= -638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010000; // iC=-1520 
vC = 14'b1111110101010000; // vC= -688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010101; // iC=-1579 
vC = 14'b1111110100000110; // vC= -762 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100110; // iC=-1434 
vC = 14'b1111110101111000; // vC= -648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001001; // iC=-1463 
vC = 14'b1111110101100101; // vC= -667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100101; // iC=-1563 
vC = 14'b1111110011111111; // vC= -769 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001111; // iC=-1457 
vC = 14'b1111110101010100; // vC= -684 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b1111110100011011; // vC= -741 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b1111110101110111; // vC= -649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100101; // iC=-1499 
vC = 14'b1111110101110011; // vC= -653 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110011; // iC=-1549 
vC = 14'b1111110100011110; // vC= -738 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010001; // iC=-1455 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111010; // iC=-1414 
vC = 14'b1111110100111101; // vC= -707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b1111110011010111; // vC= -809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001000; // iC=-1528 
vC = 14'b1111110011101001; // vC= -791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010111; // iC=-1385 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000100; // iC=-1532 
vC = 14'b1111110011100111; // vC= -793 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110100; // iC=-1420 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100000; // iC=-1504 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100101; // iC=-1371 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100100; // iC=-1372 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b1111110010011010; // vC= -870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010111; // iC=-1449 
vC = 14'b1111110100000100; // vC= -764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111001; // iC=-1351 
vC = 14'b1111110010111111; // vC= -833 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000011; // iC=-1405 
vC = 14'b1111110010010110; // vC= -874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000111; // iC=-1465 
vC = 14'b1111110100000010; // vC= -766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100010; // iC=-1438 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101111; // iC=-1361 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000001; // iC=-1343 
vC = 14'b1111110010110100; // vC= -844 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111110010011110; // vC= -866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001001; // iC=-1399 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001011; // iC=-1397 
vC = 14'b1111110011011011; // vC= -805 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111111; // iC=-1345 
vC = 14'b1111110001011011; // vC= -933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b1111110010000000; // vC= -896 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001101; // iC=-1395 
vC = 14'b1111110010100110; // vC= -858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110110; // iC=-1354 
vC = 14'b1111110010100000; // vC= -864 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010110; // iC=-1322 
vC = 14'b1111110001101000; // vC= -920 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000000; // iC=-1408 
vC = 14'b1111110001101011; // vC= -917 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011100010; // iC=-1310 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100001; // iC=-1439 
vC = 14'b1111110010100111; // vC= -857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010000; // iC=-1392 
vC = 14'b1111110010011110; // vC= -866 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001001; // iC=-1335 
vC = 14'b1111110010010001; // vC= -879 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001011; // iC=-1269 
vC = 14'b1111110000101101; // vC= -979 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010000; // iC=-1328 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111110010000001; // vC= -895 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111001; // iC=-1287 
vC = 14'b1111110001001100; // vC= -948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000010; // iC=-1406 
vC = 14'b1111110001011000; // vC= -936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111100; // iC=-1348 
vC = 14'b1111110001000100; // vC= -956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001111; // iC=-1329 
vC = 14'b1111110000111111; // vC= -961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110111; // iC=-1289 
vC = 14'b1111110001111100; // vC= -900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101011; // iC=-1301 
vC = 14'b1111110001010000; // vC= -944 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001000; // iC=-1272 
vC = 14'b1111110010001101; // vC= -883 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110101; // iC=-1355 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101110; // iC=-1298 
vC = 14'b1111110010001011; // vC= -885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101000; // iC=-1304 
vC = 14'b1111110000110011; // vC= -973 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011000; // iC=-1256 
vC = 14'b1111110000001101; // vC=-1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101100; // iC=-1236 
vC = 14'b1111110001110100; // vC= -908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111010; // iC=-1222 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000011; // iC=-1213 
vC = 14'b1111110000001001; // vC=-1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101001; // iC=-1303 
vC = 14'b1111110001001100; // vC= -948 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011010; // iC=-1190 
vC = 14'b1111101111100111; // vC=-1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010010; // iC=-1326 
vC = 14'b1111101111100010; // vC=-1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011101; // iC=-1187 
vC = 14'b1111101111110010; // vC=-1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100101; // iC=-1243 
vC = 14'b1111110000101100; // vC= -980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011111; // iC=-1249 
vC = 14'b1111101111111000; // vC=-1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101110; // iC=-1234 
vC = 14'b1111101111101001; // vC=-1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001110; // iC=-1202 
vC = 14'b1111101111001110; // vC=-1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011011111; // iC=-1313 
vC = 14'b1111101110110100; // vC=-1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100010; // iC=-1182 
vC = 14'b1111110000111001; // vC= -967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001111; // iC=-1265 
vC = 14'b1111101111011001; // vC=-1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000001; // iC=-1215 
vC = 14'b1111110000110001; // vC= -975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100011; // iC=-1245 
vC = 14'b1111101111111110; // vC=-1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000001; // iC=-1215 
vC = 14'b1111101110110101; // vC=-1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110100; // iC=-1292 
vC = 14'b1111101111100010; // vC=-1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111010; // iC=-1286 
vC = 14'b1111101110011010; // vC=-1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101101; // iC=-1235 
vC = 14'b1111101110010001; // vC=-1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001100; // iC=-1268 
vC = 14'b1111101111011101; // vC=-1059 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001001; // iC=-1271 
vC = 14'b1111101110001010; // vC=-1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100001; // iC=-1183 
vC = 14'b1111101111101000; // vC=-1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111111; // iC=-1217 
vC = 14'b1111110000010100; // vC=-1004 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011101; // iC=-1251 
vC = 14'b1111101111000111; // vC=-1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101000010; // iC=-1214 
vC = 14'b1111101101111101; // vC=-1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101111; // iC=-1105 
vC = 14'b1111110000001000; // vC=-1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100100; // iC=-1180 
vC = 14'b1111101110110100; // vC=-1100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000100; // iC=-1084 
vC = 14'b1111101110011110; // vC=-1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101101110; // iC=-1170 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111101; // iC=-1155 
vC = 14'b1111101101110110; // vC=-1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100101; // iC=-1179 
vC = 14'b1111101110101110; // vC=-1106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101010; // iC=-1110 
vC = 14'b1111101111010000; // vC=-1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001100; // iC=-1076 
vC = 14'b1111101110010111; // vC=-1129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011011; // iC=-1125 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000111; // iC=-1081 
vC = 14'b1111101110011001; // vC=-1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110111; // iC=-1097 
vC = 14'b1111101101001000; // vC=-1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111100; // iC=-1156 
vC = 14'b1111101110001000; // vC=-1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101010; // iC=-1110 
vC = 14'b1111101111001101; // vC=-1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101110; // iC=-1042 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011011; // iC=-1125 
vC = 14'b1111101111001011; // vC=-1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000101; // iC=-1019 
vC = 14'b1111101101110001; // vC=-1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101101; // iC=-1043 
vC = 14'b1111101101000110; // vC=-1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011110; // iC=-1122 
vC = 14'b1111101110011001; // vC=-1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111100; // iC=-1092 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001010; // iC=-1078 
vC = 14'b1111101101000110; // vC=-1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111101; // iC=-1091 
vC = 14'b1111101101101101; // vC=-1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001010; // iC=-1142 
vC = 14'b1111101100100101; // vC=-1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000100; // iC=-1020 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000011001; // iC= -999 
vC = 14'b1111101100111111; // vC=-1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000011; // iC=-1085 
vC = 14'b1111101110011111; // vC=-1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011100; // iC=-1124 
vC = 14'b1111101101010101; // vC=-1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110110; // iC=-1034 
vC = 14'b1111101101011011; // vC=-1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101101; // iC=-1107 
vC = 14'b1111101100000101; // vC=-1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011100; // iC=-1060 
vC = 14'b1111101101101111; // vC=-1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110111; // iC=-1097 
vC = 14'b1111101100010110; // vC=-1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111110; // iC=-1026 
vC = 14'b1111101100001100; // vC=-1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000010; // iC= -958 
vC = 14'b1111101101011010; // vC=-1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101111; // iC=-1041 
vC = 14'b1111101100011101; // vC=-1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000001; // iC= -959 
vC = 14'b1111101101110110; // vC=-1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111111; // iC= -961 
vC = 14'b1111101101111011; // vC=-1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111101; // iC= -963 
vC = 14'b1111101100010110; // vC=-1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100111; // iC=-1049 
vC = 14'b1111101101100100; // vC=-1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011101; // iC= -931 
vC = 14'b1111101100000100; // vC=-1276 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111101011101101; // vC=-1299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000000; // iC= -960 
vC = 14'b1111101101100111; // vC=-1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110011; // iC=-1037 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111001; // iC= -903 
vC = 14'b1111101101011000; // vC=-1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011100; // iC= -932 
vC = 14'b1111101101000011; // vC=-1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110001; // iC= -911 
vC = 14'b1111101100110011; // vC=-1229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111000; // iC=-1032 
vC = 14'b1111101011100010; // vC=-1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110010; // iC= -974 
vC = 14'b1111101101011000; // vC=-1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b1111101011111100; // vC=-1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000000; // iC= -896 
vC = 14'b1111101101001111; // vC=-1201 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101000; // iC= -856 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001111; // iC= -945 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000111000; // iC= -968 
vC = 14'b1111101101001000; // vC=-1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011100; // iC= -932 
vC = 14'b1111101100011001; // vC=-1255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010010; // iC= -942 
vC = 14'b1111101011001010; // vC=-1334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000111; // iC= -825 
vC = 14'b1111101011110100; // vC=-1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101000; // iC= -856 
vC = 14'b1111101011110000; // vC=-1296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001000; // iC= -824 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100000; // iC= -864 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110100; // iC= -844 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010000; // iC= -880 
vC = 14'b1111101011100111; // vC=-1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010010; // iC= -942 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010011; // iC= -813 
vC = 14'b1111101100000010; // vC=-1278 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010110; // iC= -810 
vC = 14'b1111101011011010; // vC=-1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001101; // iC= -883 
vC = 14'b1111101010110111; // vC=-1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010011; // iC= -813 
vC = 14'b1111101100011101; // vC=-1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111011; // iC= -901 
vC = 14'b1111101010010011; // vC=-1389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001010; // iC= -822 
vC = 14'b1111101010110011; // vC=-1357 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000011; // iC= -893 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001010; // iC= -758 
vC = 14'b1111101010111010; // vC=-1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001011; // iC= -821 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011000; // iC= -744 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100000; // iC= -800 
vC = 14'b1111101100001110; // vC=-1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110111; // iC= -777 
vC = 14'b1111101010011001; // vC=-1383 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011110; // iC= -866 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101110; // iC= -786 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011000000; // iC= -832 
vC = 14'b1111101010101100; // vC=-1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010010; // iC= -750 
vC = 14'b1111101010001000; // vC=-1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110101; // iC= -843 
vC = 14'b1111101010111101; // vC=-1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010110; // iC= -810 
vC = 14'b1111101010101010; // vC=-1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100111; // iC= -729 
vC = 14'b1111101011011111; // vC=-1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001001; // iC= -823 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100110; // iC= -794 
vC = 14'b1111101011110001; // vC=-1295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011100; // iC= -676 
vC = 14'b1111101010111101; // vC=-1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111110; // iC= -706 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111100; // iC= -708 
vC = 14'b1111101011010110; // vC=-1322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110001; // iC= -783 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000100; // iC= -764 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110011; // iC= -717 
vC = 14'b1111101010110010; // vC=-1358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100011; // iC= -733 
vC = 14'b1111101001011110; // vC=-1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010100; // iC= -748 
vC = 14'b1111101010110100; // vC=-1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000011; // iC= -701 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000101; // iC= -699 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100100; // iC= -668 
vC = 14'b1111101001000110; // vC=-1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110010; // iC= -718 
vC = 14'b1111101010111001; // vC=-1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010011; // iC= -621 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101011; // iC= -661 
vC = 14'b1111101001111111; // vC=-1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000000; // iC= -704 
vC = 14'b1111101010010100; // vC=-1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100010; // iC= -606 
vC = 14'b1111101001000000; // vC=-1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000000; // iC= -704 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111110; // iC= -578 
vC = 14'b1111101010101000; // vC=-1368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100101; // iC= -731 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101000001; // iC= -703 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100101; // iC= -603 
vC = 14'b1111101010111110; // vC=-1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011010; // iC= -678 
vC = 14'b1111101010100111; // vC=-1369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011010; // iC= -550 
vC = 14'b1111101000101100; // vC=-1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100111101; // iC= -707 
vC = 14'b1111101000011010; // vC=-1510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011010; // iC= -678 
vC = 14'b1111101001011110; // vC=-1442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111010; // iC= -582 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000011; // iC= -573 
vC = 14'b1111101010011101; // vC=-1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101010; // iC= -534 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100110; // iC= -666 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110000; // iC= -656 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000101; // iC= -507 
vC = 14'b1111101001101100; // vC=-1428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011011; // iC= -549 
vC = 14'b1111101010100101; // vC=-1371 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001001; // iC= -503 
vC = 14'b1111101010001110; // vC=-1394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110100111; // iC= -601 
vC = 14'b1111101000100011; // vC=-1501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011001; // iC= -615 
vC = 14'b1111101000110111; // vC=-1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001101; // iC= -499 
vC = 14'b1111101001100111; // vC=-1433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010001; // iC= -623 
vC = 14'b1111100111111100; // vC=-1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101101; // iC= -467 
vC = 14'b1111101001111100; // vC=-1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000010; // iC= -510 
vC = 14'b1111101000011011; // vC=-1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000010; // iC= -574 
vC = 14'b1111101001111010; // vC=-1414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010001; // iC= -495 
vC = 14'b1111101010001001; // vC=-1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000000; // iC= -512 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011110; // iC= -482 
vC = 14'b1111101000111111; // vC=-1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000110; // iC= -570 
vC = 14'b1111101000011011; // vC=-1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010101; // iC= -427 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100000; // iC= -544 
vC = 14'b1111100111101110; // vC=-1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001010011; // iC= -429 
vC = 14'b1111101000100000; // vC=-1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b1111100111111011; // vC=-1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100111; // iC= -473 
vC = 14'b1111101001110111; // vC=-1417 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101110; // iC= -466 
vC = 14'b1111101000000000; // vC=-1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100010; // iC= -414 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000000100; // iC= -508 
vC = 14'b1111101001010100; // vC=-1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001110; // iC= -434 
vC = 14'b1111101000001101; // vC=-1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111100; // iC= -388 
vC = 14'b1111100111100001; // vC=-1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001101; // iC= -499 
vC = 14'b1111101000011101; // vC=-1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000011; // iC= -381 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111101; // iC= -387 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011111; // iC= -481 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001011001; // iC= -423 
vC = 14'b1111100111011001; // vC=-1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000001; // iC= -383 
vC = 14'b1111100111110111; // vC=-1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110101; // iC= -459 
vC = 14'b1111101000101111; // vC=-1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100111; // iC= -409 
vC = 14'b1111101000010111; // vC=-1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001101111; // iC= -401 
vC = 14'b1111101000100011; // vC=-1501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001001; // iC= -375 
vC = 14'b1111101000010001; // vC=-1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111000; // iC= -328 
vC = 14'b1111101000010010; // vC=-1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010101000; // iC= -344 
vC = 14'b1111100111001110; // vC=-1586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111111; // iC= -385 
vC = 14'b1111101001101001; // vC=-1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110111; // iC= -265 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100001; // iC= -287 
vC = 14'b1111101000001100; // vC=-1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011001; // iC= -231 
vC = 14'b1111101000000000; // vC=-1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000001; // iC= -255 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001000; // iC= -248 
vC = 14'b1111100111011110; // vC=-1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010100; // iC= -172 
vC = 14'b1111101001011100; // vC=-1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100001011; // iC= -245 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000011; // iC= -125 
vC = 14'b1111100111010110; // vC=-1578 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111101; // iC= -131 
vC = 14'b1111101000011110; // vC=-1506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100010001; // iC= -239 
vC = 14'b1111100111011111; // vC=-1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011000; // iC= -104 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110000011; // iC= -125 
vC = 14'b1111100111101010; // vC=-1558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101000000; // iC= -192 
vC = 14'b1111100111010100; // vC=-1580 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111110; // iC= -130 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011111; // iC=  -33 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101011; // iC= -149 
vC = 14'b1111101000001001; // vC=-1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000000110; // iC=    6 
vC = 14'b1111101001100001; // vC=-1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011011; // iC= -101 
vC = 14'b1111101000000010; // vC=-1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100111; // iC=  -89 
vC = 14'b1111101001000100; // vC=-1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111101; // iC=   61 
vC = 14'b1111100111000111; // vC=-1593 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111000; // iC=   -8 
vC = 14'b1111100111000011; // vC=-1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111011000; // iC=  -40 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011101; // iC=   29 
vC = 14'b1111100111101011; // vC=-1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000010111; // iC=   23 
vC = 14'b1111100111110011; // vC=-1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001111; // iC=  143 
vC = 14'b1111100111110111; // vC=-1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001111101; // iC=  125 
vC = 14'b1111100111011110; // vC=-1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001101; // iC=  141 
vC = 14'b1111101000110100; // vC=-1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001101; // iC=   77 
vC = 14'b1111101001010010; // vC=-1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001100; // iC=  140 
vC = 14'b1111100111101110; // vC=-1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010010000; // iC=  144 
vC = 14'b1111101001010100; // vC=-1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011110; // iC=  222 
vC = 14'b1111101000110101; // vC=-1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111110; // iC=  254 
vC = 14'b1111101000011011; // vC=-1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100100000; // iC=  288 
vC = 14'b1111100111110001; // vC=-1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000001; // iC=  321 
vC = 14'b1111101000001100; // vC=-1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101101; // iC=  237 
vC = 14'b1111100111110000; // vC=-1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100011; // iC=  355 
vC = 14'b1111100111100101; // vC=-1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000011; // iC=  387 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111110; // iC=  446 
vC = 14'b1111101001001111; // vC=-1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010111; // iC=  407 
vC = 14'b1111100111111100; // vC=-1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110001011; // iC=  395 
vC = 14'b1111101001100101; // vC=-1435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100101; // iC=  485 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111000; // iC=  440 
vC = 14'b1111100111100000; // vC=-1568 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011101; // iC=  477 
vC = 14'b1111100111111101; // vC=-1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111111; // iC=  575 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101100; // iC=  556 
vC = 14'b1111100111111011; // vC=-1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111000; // iC=  632 
vC = 14'b1111101000001000; // vC=-1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111111; // iC=  511 
vC = 14'b1111101001011010; // vC=-1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010110; // iC=  662 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001011; // iC=  651 
vC = 14'b1111101001000000; // vC=-1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010101; // iC=  725 
vC = 14'b1111100111111100; // vC=-1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010000; // iC=  656 
vC = 14'b1111100111110000; // vC=-1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001101; // iC=  781 
vC = 14'b1111101001111110; // vC=-1410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010101; // iC=  789 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001101; // iC=  717 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100110; // iC=  806 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100110; // iC=  870 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101010110; // iC=  854 
vC = 14'b1111101000110000; // vC=-1488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000000; // iC=  896 
vC = 14'b1111101000000100; // vC=-1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100101; // iC=  869 
vC = 14'b1111101000000101; // vC=-1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110100; // iC=  884 
vC = 14'b1111101000010010; // vC=-1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000010; // iC=  834 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101101; // iC=  941 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011101; // iC=  925 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100111; // iC=  935 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101100; // iC= 1068 
vC = 14'b1111101010100010; // vC=-1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111011; // iC=  955 
vC = 14'b1111101000110011; // vC=-1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001011; // iC= 1035 
vC = 14'b1111101001111100; // vC=-1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101100; // iC= 1004 
vC = 14'b1111101010101111; // vC=-1361 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000011; // iC= 1027 
vC = 14'b1111101001001110; // vC=-1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001111; // iC= 1167 
vC = 14'b1111101000111100; // vC=-1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001111; // iC= 1039 
vC = 14'b1111101000111100; // vC=-1476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011111; // iC= 1183 
vC = 14'b1111101000110011; // vC=-1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000011; // iC= 1091 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101001; // iC= 1129 
vC = 14'b1111101010010111; // vC=-1385 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010111; // iC= 1239 
vC = 14'b1111101001100110; // vC=-1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100101; // iC= 1253 
vC = 14'b1111101011010101; // vC=-1323 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010111; // iC= 1303 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100011; // iC= 1187 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111101; // iC= 1277 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001010; // iC= 1290 
vC = 14'b1111101001101000; // vC=-1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011100; // iC= 1372 
vC = 14'b1111101010011101; // vC=-1379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100000; // iC= 1312 
vC = 14'b1111101010011110; // vC=-1378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100111; // iC= 1383 
vC = 14'b1111101011100010; // vC=-1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111000; // iC= 1400 
vC = 14'b1111101011111011; // vC=-1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001111; // iC= 1359 
vC = 14'b1111101010100010; // vC=-1374 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111011; // iC= 1339 
vC = 14'b1111101011000011; // vC=-1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111000111; // iC= 1479 
vC = 14'b1111101001111100; // vC=-1412 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000001; // iC= 1409 
vC = 14'b1111101010111011; // vC=-1349 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010011; // iC= 1491 
vC = 14'b1111101011010111; // vC=-1321 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010011; // iC= 1491 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111001; // iC= 1401 
vC = 14'b1111101011100110; // vC=-1306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110101; // iC= 1525 
vC = 14'b1111101010100100; // vC=-1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011100; // iC= 1564 
vC = 14'b1111101010101011; // vC=-1365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111001; // iC= 1593 
vC = 14'b1111101011101100; // vC=-1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101011; // iC= 1515 
vC = 14'b1111101100100101; // vC=-1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111010; // iC= 1530 
vC = 14'b1111101011000000; // vC=-1344 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100000; // iC= 1504 
vC = 14'b1111101011001111; // vC=-1329 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110111; // iC= 1591 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000100; // iC= 1604 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011011; // iC= 1563 
vC = 14'b1111101011000011; // vC=-1341 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011111; // iC= 1567 
vC = 14'b1111101011101111; // vC=-1297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101001; // iC= 1641 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010111; // iC= 1687 
vC = 14'b1111101100001110; // vC=-1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111011; // iC= 1659 
vC = 14'b1111101101101110; // vC=-1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111111; // iC= 1599 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100011; // iC= 1699 
vC = 14'b1111101100111111; // vC=-1217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000000; // iC= 1664 
vC = 14'b1111101100101101; // vC=-1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011111; // iC= 1759 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111001; // iC= 1657 
vC = 14'b1111101101011001; // vC=-1191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b1111101101101000; // vC=-1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000100; // iC= 1668 
vC = 14'b1111101100000011; // vC=-1277 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000011; // iC= 1795 
vC = 14'b1111101101000011; // vC=-1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000101; // iC= 1797 
vC = 14'b1111101100101100; // vC=-1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b1111101110110010; // vC=-1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b1111101101001110; // vC=-1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b1111101100100100; // vC=-1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101011; // iC= 1771 
vC = 14'b1111101110011110; // vC=-1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b1111101101101100; // vC=-1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b1111101101011011; // vC=-1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100111; // iC= 1767 
vC = 14'b1111101111000001; // vC=-1087 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011001; // iC= 1881 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111101; // iC= 1789 
vC = 14'b1111101110110001; // vC=-1103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111101110011110; // vC=-1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011000; // iC= 1880 
vC = 14'b1111101111100101; // vC=-1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b1111110000000011; // vC=-1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010000; // iC= 1872 
vC = 14'b1111101101111100; // vC=-1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010101; // iC= 1877 
vC = 14'b1111101110010101; // vC=-1131 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000111; // iC= 1799 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010000; // iC= 1808 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000111; // iC= 1799 
vC = 14'b1111101110110110; // vC=-1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111101110011100; // vC=-1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b1111101110101001; // vC=-1111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111101111110000; // vC=-1040 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b1111101110111111; // vC=-1089 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111110000011101; // vC= -995 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b1111101110111101; // vC=-1091 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111101111101010; // vC=-1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111101111110011; // vC=-1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b1111101111111100; // vC=-1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b1111101111011010; // vC=-1062 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001110; // iC= 1934 
vC = 14'b1111110000110001; // vC= -975 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b1111110000111111; // vC= -961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001101; // iC= 1869 
vC = 14'b1111101111101010; // vC=-1046 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b1111110001101010; // vC= -918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111101111111000; // vC=-1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111101111111111; // vC=-1025 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b1111110000101011; // vC= -981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111010; // iC= 1914 
vC = 14'b1111110000110010; // vC= -974 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000111; // iC= 1863 
vC = 14'b1111110000010111; // vC=-1001 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111110001110111; // vC= -905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011100; // iC= 1948 
vC = 14'b1111110000100001; // vC= -991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001010; // iC= 1866 
vC = 14'b1111110001110111; // vC= -905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b1111110010111000; // vC= -840 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111110001111100; // vC= -900 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110001000110; // vC= -954 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011110; // iC= 1886 
vC = 14'b1111110011001000; // vC= -824 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b1111110001100110; // vC= -922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011001; // iC= 2009 
vC = 14'b1111110001111111; // vC= -897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b1111110001011100; // vC= -932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111110011000100; // vC= -828 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111110010010110; // vC= -874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b1111110100010001; // vC= -751 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111110011100010; // vC= -798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b1111110010001011; // vC= -885 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b1111110011011000; // vC= -808 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000100; // iC= 1988 
vC = 14'b1111110011100010; // vC= -798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011100; // iC= 1948 
vC = 14'b1111110011000000; // vC= -832 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b1111110011100001; // vC= -799 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111110011110001; // vC= -783 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b1111110101010110; // vC= -682 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b1111110011110011; // vC= -781 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b1111110101000111; // vC= -697 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111110011010111; // vC= -809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111101; // iC= 2045 
vC = 14'b1111110011011111; // vC= -801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111110101001110; // vC= -690 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001001; // iC= 1993 
vC = 14'b1111110101100010; // vC= -670 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001111; // iC= 2063 
vC = 14'b1111110101011001; // vC= -679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b1111110100010010; // vC= -750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111110100011100; // vC= -740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111110110000001; // vC= -639 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100000; // iC= 2016 
vC = 14'b1111110100100110; // vC= -730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b1111110100111110; // vC= -706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110111; // iC= 1975 
vC = 14'b1111110101011011; // vC= -677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001011; // iC= 1995 
vC = 14'b1111110101100101; // vC= -667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100010; // iC= 2018 
vC = 14'b1111110110010000; // vC= -624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111110111011010; // vC= -550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b1111110101110001; // vC= -655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001110; // iC= 2062 
vC = 14'b1111110110010000; // vC= -624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b1111110111000110; // vC= -570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111110110100010; // vC= -606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110101111100; // vC= -644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000000; // iC= 1984 
vC = 14'b1111110110110110; // vC= -586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111110110111111; // vC= -577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b1111110101111101; // vC= -643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b1111110111101001; // vC= -535 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b1111110110100110; // vC= -602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001100; // iC= 1996 
vC = 14'b1111110110110111; // vC= -585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111110111110100; // vC= -524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000101; // iC= 2053 
vC = 14'b1111110110101101; // vC= -595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b1111110111000100; // vC= -572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111110111101010; // vC= -534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111110110110011; // vC= -589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001111; // iC= 2063 
vC = 14'b1111111000001001; // vC= -503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111111000101010; // vC= -470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b1111111000011011; // vC= -485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111110111001010; // vC= -566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011111; // iC= 2079 
vC = 14'b1111110111010111; // vC= -553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111111000000111; // vC= -505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111111000111101; // vC= -451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111111001110110; // vC= -394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111111000111100; // vC= -452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111111000110100; // vC= -460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111111; // iC= 2047 
vC = 14'b1111111000010010; // vC= -494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010010; // iC= 2066 
vC = 14'b1111111001101010; // vC= -406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111111001001111; // vC= -433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111111000100111; // vC= -473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011001; // iC= 2073 
vC = 14'b1111111001100111; // vC= -409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000101001; // iC= 2089 
vC = 14'b1111111010100110; // vC= -346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000101010; // iC= 2090 
vC = 14'b1111111000110010; // vC= -462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010011; // iC= 1939 
vC = 14'b1111111010111001; // vC= -327 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111111010001110; // vC= -370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111111001100000; // vC= -416 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b1111111001010011; // vC= -429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101101; // iC= 2029 
vC = 14'b1111111001101000; // vC= -408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100111; // iC= 2087 
vC = 14'b1111111010110011; // vC= -333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111001100010; // vC= -414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000100000; // iC= 2080 
vC = 14'b1111111010011000; // vC= -360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110100; // iC= 1972 
vC = 14'b1111111011000000; // vC= -320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b1111111010011101; // vC= -355 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111111010100111; // vC= -345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011011; // iC= 2011 
vC = 14'b1111111010110100; // vC= -332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010001; // iC= 2065 
vC = 14'b1111111100001100; // vC= -244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011000; // iC= 2072 
vC = 14'b1111111010011110; // vC= -354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110000; // iC= 2032 
vC = 14'b1111111100100000; // vC= -224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010101; // iC= 2005 
vC = 14'b1111111010110000; // vC= -336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110101; // iC= 2037 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b1111111011000111; // vC= -313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111100; // iC= 2044 
vC = 14'b1111111010111011; // vC= -325 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111011100100; // vC= -284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b1111111101001110; // vC= -178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111100; // iC= 2044 
vC = 14'b1111111011110101; // vC= -267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001000; // iC= 2056 
vC = 14'b1111111100100011; // vC= -221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010100; // iC= 2004 
vC = 14'b1111111011010111; // vC= -297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000100; // iC= 1924 
vC = 14'b1111111101100111; // vC= -153 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001101; // iC= 2061 
vC = 14'b1111111101000010; // vC= -190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111111101011100; // vC= -164 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111101100011; // vC= -157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010011; // iC= 2067 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000010; // iC= 1986 
vC = 14'b1111111100000111; // vC= -249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010010; // iC= 2002 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111111101100100; // vC= -156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111111100100010; // vC= -222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011100; // iC= 1948 
vC = 14'b1111111110100101; // vC=  -91 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101110; // iC= 2030 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011010; // iC= 2074 
vC = 14'b1111111101101001; // vC= -151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111111110110101; // vC=  -75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001011; // iC= 2059 
vC = 14'b1111111110000001; // vC= -127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011000; // iC= 2008 
vC = 14'b1111111101100110; // vC= -154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111111110011001; // vC= -103 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b1111111101111010; // vC= -134 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111111101101101; // vC= -147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111111110110010; // vC=  -78 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110100; // iC= 2036 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010011; // iC= 2067 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111111110000001; // vC= -127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110111; // iC= 1975 
vC = 14'b0000000000010100; // vC=   20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b1111111110111111; // vC=  -65 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000000; // iC= 2048 
vC = 14'b1111111110101110; // vC=  -82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001000; // iC= 2056 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b1111111111110100; // vC=  -12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b0000000000110110; // vC=   54 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100010; // iC= 2018 
vC = 14'b0000000000110001; // vC=   49 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b1111111111110010; // vC=  -14 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100110; // iC= 2022 
vC = 14'b0000000000110111; // vC=   55 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111111111001110; // vC=  -50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b0000000001000011; // vC=   67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000001; // iC= 2049 
vC = 14'b0000000000100000; // vC=   32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111111111000110; // vC=  -58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b1111111111111010; // vC=   -6 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b0000000000011000; // vC=   24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011111; // iC= 2015 
vC = 14'b1111111111101010; // vC=  -22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b0000000000100001; // vC=   33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b0000000000100000; // vC=   32 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b0000000000110000; // vC=   48 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b0000000001111100; // vC=  124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b0000000001010000; // vC=   80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101100; // iC= 1900 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000001011100; // vC=   92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b0000000001100101; // vC=  101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000110; // iC= 1926 
vC = 14'b0000000000011011; // vC=   27 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b0000000010011010; // vC=  154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b0000000001011111; // vC=   95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110011; // iC= 1907 
vC = 14'b0000000001101111; // vC=  111 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100011; // iC= 2019 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111110; // iC= 1982 
vC = 14'b0000000011010101; // vC=  213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b0000000001101011; // vC=  107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011100; // iC= 1948 
vC = 14'b0000000010101101; // vC=  173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b0000000010101011; // vC=  171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110000; // iC= 1904 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b0000000010111011; // vC=  187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000000010011111; // vC=  159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b0000000010001111; // vC=  143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b0000000010110010; // vC=  178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b0000000010100111; // vC=  167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b0000000011100001; // vC=  225 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011101; // iC= 2013 
vC = 14'b0000000011100000; // vC=  224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b0000000011100000; // vC=  224 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110101; // iC= 1973 
vC = 14'b0000000011010010; // vC=  210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b0000000010100010; // vC=  162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010100; // iC= 1940 
vC = 14'b0000000011111000; // vC=  248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001100; // iC= 1932 
vC = 14'b0000000010101101; // vC=  173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b0000000011100111; // vC=  231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111010; // iC= 1850 
vC = 14'b0000000011110100; // vC=  244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000100; // iC= 1924 
vC = 14'b0000000011110011; // vC=  243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b0000000011000010; // vC=  194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b0000000100100000; // vC=  288 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b0000000011111000; // vC=  248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001101; // iC= 1997 
vC = 14'b0000000011100101; // vC=  229 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101000; // iC= 1832 
vC = 14'b0000000101101011; // vC=  363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b0000000101110111; // vC=  375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b0000000101010010; // vC=  338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b0000000101100001; // vC=  353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000000100000100; // vC=  260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010111; // iC= 1943 
vC = 14'b0000000101010100; // vC=  340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b0000000101100100; // vC=  356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b0000000110010100; // vC=  404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b0000000110001111; // vC=  399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b0000000101111011; // vC=  379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000000100100111; // vC=  295 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b0000000101110101; // vC=  373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b0000000110001110; // vC=  398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b0000000110001001; // vC=  393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000110001000; // vC=  392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101110; // iC= 1838 
vC = 14'b0000000101011110; // vC=  350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b0000000110110000; // vC=  432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b0000000110111110; // vC=  446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b0000000111011101; // vC=  477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011101; // iC= 1885 
vC = 14'b0000000111001010; // vC=  458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111000; // iC= 1848 
vC = 14'b0000000111111110; // vC=  510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b0000000101111110; // vC=  382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100000; // iC= 1888 
vC = 14'b0000000110110001; // vC=  433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101111; // iC= 1839 
vC = 14'b0000000110000010; // vC=  386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000100; // iC= 1860 
vC = 14'b0000000111101011; // vC=  491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001011; // iC= 1867 
vC = 14'b0000000110000100; // vC=  388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000011; // iC= 1859 
vC = 14'b0000001000000111; // vC=  519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b0000000111100110; // vC=  486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000001000110000; // vC=  560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b0000000110110111; // vC=  439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110011; // iC= 1843 
vC = 14'b0000001000100001; // vC=  545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b0000000111110010; // vC=  498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000001001001100; // vC=  588 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b0000001000100001; // vC=  545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b0000000110111010; // vC=  442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001101; // iC= 1869 
vC = 14'b0000001000001101; // vC=  525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100001; // iC= 1825 
vC = 14'b0000000111011101; // vC=  477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011001; // iC= 1753 
vC = 14'b0000000111100100; // vC=  484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101001; // iC= 1897 
vC = 14'b0000001001100100; // vC=  612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b0000001001100111; // vC=  615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b0000001001000101; // vC=  581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010010; // iC= 1874 
vC = 14'b0000001001100110; // vC=  614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010110; // iC= 1878 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011011; // iC= 1819 
vC = 14'b0000001000111001; // vC=  569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b0000001010010111; // vC=  663 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001010; // iC= 1866 
vC = 14'b0000001010010110; // vC=  662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b0000001000101101; // vC=  557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101101; // iC= 1773 
vC = 14'b0000001001100110; // vC=  614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b0000001000100110; // vC=  550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000001001110011; // vC=  627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b0000001001110011; // vC=  627 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111011; // iC= 1723 
vC = 14'b0000001000110001; // vC=  561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000001010001011; // vC=  651 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110010; // iC= 1714 
vC = 14'b0000001001100000; // vC=  608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101100; // iC= 1772 
vC = 14'b0000001011000011; // vC=  707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100000; // iC= 1760 
vC = 14'b0000001001111000; // vC=  632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000011; // iC= 1731 
vC = 14'b0000001010000001; // vC=  641 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011100; // iC= 1820 
vC = 14'b0000001010111010; // vC=  698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b0000001001110001; // vC=  625 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b0000001010110011; // vC=  691 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001000; // iC= 1672 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000101; // iC= 1797 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b0000001011101110; // vC=  750 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b0000001011001111; // vC=  719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010010110; // iC= 1686 
vC = 14'b0000001100010000; // vC=  784 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001001; // iC= 1801 
vC = 14'b0000001011100111; // vC=  743 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b0000001010001000; // vC=  648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001100; // iC= 1740 
vC = 14'b0000001010111011; // vC=  699 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110110; // iC= 1654 
vC = 14'b0000001010111111; // vC=  703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b0000001011010110; // vC=  726 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b0000001010011011; // vC=  667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101101; // iC= 1645 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000100; // iC= 1668 
vC = 14'b0000001100101110; // vC=  814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b0000001011001011; // vC=  715 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011011; // iC= 1691 
vC = 14'b0000001011110011; // vC=  755 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101001; // iC= 1769 
vC = 14'b0000001100100001; // vC=  801 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b0000001010111100; // vC=  700 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001010; // iC= 1610 
vC = 14'b0000001100111010; // vC=  826 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011100; // iC= 1692 
vC = 14'b0000001100000011; // vC=  771 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010100; // iC= 1748 
vC = 14'b0000001100101001; // vC=  809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110100; // iC= 1716 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111101; // iC= 1725 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011011; // iC= 1755 
vC = 14'b0000001101011100; // vC=  860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001101; // iC= 1677 
vC = 14'b0000001100111110; // vC=  830 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b0000001100001110; // vC=  782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111100; // iC= 1724 
vC = 14'b0000001110001001; // vC=  905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000110; // iC= 1670 
vC = 14'b0000001110001001; // vC=  905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000101; // iC= 1605 
vC = 14'b0000001101101010; // vC=  874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100101; // iC= 1573 
vC = 14'b0000001100011100; // vC=  796 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000111; // iC= 1607 
vC = 14'b0000001100111011; // vC=  827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111011; // iC= 1659 
vC = 14'b0000001110010010; // vC=  914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111010; // iC= 1722 
vC = 14'b0000001101001001; // vC=  841 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001010; // iC= 1610 
vC = 14'b0000001100100111; // vC=  807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100010; // iC= 1570 
vC = 14'b0000001101011001; // vC=  857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101110; // iC= 1646 
vC = 14'b0000001101010100; // vC=  852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000110; // iC= 1606 
vC = 14'b0000001110010010; // vC=  914 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b0000001100111001; // vC=  825 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111001; // iC= 1657 
vC = 14'b0000001100101111; // vC=  815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101111; // iC= 1583 
vC = 14'b0000001100111011; // vC=  827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b0000001110110001; // vC=  945 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001010; // iC= 1674 
vC = 14'b0000001101100101; // vC=  869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000000; // iC= 1536 
vC = 14'b0000001101101101; // vC=  877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b0000001110001100; // vC=  908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001000; // iC= 1608 
vC = 14'b0000001110101010; // vC=  938 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111010; // iC= 1658 
vC = 14'b0000001110100101; // vC=  933 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110000; // iC= 1520 
vC = 14'b0000001111011110; // vC=  990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000111; // iC= 1607 
vC = 14'b0000001110100110; // vC=  934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001000; // iC= 1608 
vC = 14'b0000001111000001; // vC=  961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111101; // iC= 1597 
vC = 14'b0000001110000001; // vC=  897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100011; // iC= 1635 
vC = 14'b0000010000000010; // vC= 1026 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010000; // iC= 1488 
vC = 14'b0000001110101100; // vC=  940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000001110001000; // vC=  904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b0000001111111100; // vC= 1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100001; // iC= 1569 
vC = 14'b0000001111010001; // vC=  977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011000; // iC= 1496 
vC = 14'b0000001110001001; // vC=  905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111110; // iC= 1534 
vC = 14'b0000010000011010; // vC= 1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000010; // iC= 1602 
vC = 14'b0000001110011010; // vC=  922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010101; // iC= 1493 
vC = 14'b0000010000010101; // vC= 1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010111; // iC= 1495 
vC = 14'b0000010000010011; // vC= 1043 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010011; // iC= 1555 
vC = 14'b0000001111001100; // vC=  972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001011; // iC= 1483 
vC = 14'b0000001111111001; // vC= 1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111101; // iC= 1597 
vC = 14'b0000001111101000; // vC= 1000 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101100; // iC= 1452 
vC = 14'b0000010000101110; // vC= 1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b0000010000010101; // vC= 1045 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001010; // iC= 1546 
vC = 14'b0000001111001010; // vC=  970 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101110; // iC= 1454 
vC = 14'b0000010001001110; // vC= 1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011011; // iC= 1435 
vC = 14'b0000001111100010; // vC=  994 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001011; // iC= 1419 
vC = 14'b0000010000010100; // vC= 1044 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110101; // iC= 1525 
vC = 14'b0000010000110011; // vC= 1075 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010101; // iC= 1429 
vC = 14'b0000010001010010; // vC= 1106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011101; // iC= 1501 
vC = 14'b0000010000001011; // vC= 1035 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011001; // iC= 1433 
vC = 14'b0000010001000100; // vC= 1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111111; // iC= 1471 
vC = 14'b0000010000110010; // vC= 1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101011; // iC= 1515 
vC = 14'b0000010001010011; // vC= 1107 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100011; // iC= 1443 
vC = 14'b0000001111101011; // vC= 1003 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101010; // iC= 1514 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110101; // iC= 1525 
vC = 14'b0000010001101100; // vC= 1132 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111001; // iC= 1401 
vC = 14'b0000010000110000; // vC= 1072 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101111; // iC= 1519 
vC = 14'b0000010010000011; // vC= 1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011101; // iC= 1501 
vC = 14'b0000010001100110; // vC= 1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101110; // iC= 1454 
vC = 14'b0000010001011000; // vC= 1112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010011; // iC= 1363 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010110; // iC= 1494 
vC = 14'b0000010000010111; // vC= 1047 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010101; // iC= 1493 
vC = 14'b0000010001011100; // vC= 1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000100; // iC= 1412 
vC = 14'b0000010001100010; // vC= 1122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111100; // iC= 1340 
vC = 14'b0000010001011011; // vC= 1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101101; // iC= 1389 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001101; // iC= 1357 
vC = 14'b0000010010100100; // vC= 1188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110011; // iC= 1459 
vC = 14'b0000010000110101; // vC= 1077 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100100; // iC= 1316 
vC = 14'b0000010010111000; // vC= 1208 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001000; // iC= 1416 
vC = 14'b0000010010010110; // vC= 1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101011; // iC= 1451 
vC = 14'b0000010001001010; // vC= 1098 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101100; // iC= 1388 
vC = 14'b0000010011001100; // vC= 1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011100; // iC= 1436 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001010; // iC= 1418 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001100; // iC= 1356 
vC = 14'b0000010010101101; // vC= 1197 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010011; // iC= 1363 
vC = 14'b0000010011100001; // vC= 1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100001; // iC= 1377 
vC = 14'b0000010010110111; // vC= 1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111001; // iC= 1401 
vC = 14'b0000010001111100; // vC= 1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001111; // iC= 1359 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000110; // iC= 1286 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101011; // iC= 1323 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111100; // iC= 1276 
vC = 14'b0000010001111111; // vC= 1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100011; // iC= 1251 
vC = 14'b0000010010011010; // vC= 1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100000; // iC= 1376 
vC = 14'b0000010010110010; // vC= 1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011011; // iC= 1307 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011110; // iC= 1310 
vC = 14'b0000010010101010; // vC= 1194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011010; // iC= 1370 
vC = 14'b0000010010010110; // vC= 1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010110; // iC= 1366 
vC = 14'b0000010010010001; // vC= 1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000111; // iC= 1287 
vC = 14'b0000010011000101; // vC= 1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011111; // iC= 1247 
vC = 14'b0000010011011100; // vC= 1244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110111; // iC= 1335 
vC = 14'b0000010011001100; // vC= 1228 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100110; // iC= 1318 
vC = 14'b0000010011101010; // vC= 1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101000; // iC= 1256 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011110100; // iC= 1268 
vC = 14'b0000010010101011; // vC= 1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100000011; // iC= 1283 
vC = 14'b0000010011101001; // vC= 1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111110; // iC= 1342 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001100; // iC= 1292 
vC = 14'b0000010100100101; // vC= 1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000010011110110; // vC= 1270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011010; // iC= 1242 
vC = 14'b0000010101000010; // vC= 1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100110011; // iC= 1331 
vC = 14'b0000010011110010; // vC= 1266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111101; // iC= 1277 
vC = 14'b0000010100111001; // vC= 1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010011011; // iC= 1179 
vC = 14'b0000010100001001; // vC= 1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011111010; // iC= 1274 
vC = 14'b0000010011011011; // vC= 1243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011101001; // iC= 1257 
vC = 14'b0000010100001110; // vC= 1294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001100; // iC= 1164 
vC = 14'b0000010011101001; // vC= 1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111000; // iC= 1208 
vC = 14'b0000010011001110; // vC= 1230 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110111; // iC= 1143 
vC = 14'b0000010011010011; // vC= 1235 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001000; // iC= 1288 
vC = 14'b0000010011100100; // vC= 1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011011; // iC= 1243 
vC = 14'b0000010100100110; // vC= 1318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011011011; // iC= 1243 
vC = 14'b0000010100011000; // vC= 1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111101; // iC= 1149 
vC = 14'b0000010101001010; // vC= 1354 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101110; // iC= 1134 
vC = 14'b0000010011111010; // vC= 1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111000; // iC= 1208 
vC = 14'b0000010101111010; // vC= 1402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010111010; // iC= 1210 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001111010; // iC= 1146 
vC = 14'b0000010100011110; // vC= 1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011010111; // iC= 1239 
vC = 14'b0000010100110000; // vC= 1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001100001; // iC= 1121 
vC = 14'b0000010011110101; // vC= 1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001110; // iC= 1102 
vC = 14'b0000010100010111; // vC= 1303 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000100; // iC= 1092 
vC = 14'b0000010100111011; // vC= 1339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010100111; // iC= 1191 
vC = 14'b0000010100110010; // vC= 1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011000001; // iC= 1217 
vC = 14'b0000010101100100; // vC= 1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101001; // iC= 1129 
vC = 14'b0000010101111110; // vC= 1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010010; // iC= 1106 
vC = 14'b0000010110001101; // vC= 1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001001; // iC= 1161 
vC = 14'b0000010101110111; // vC= 1399 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001101100; // iC= 1132 
vC = 14'b0000010101100000; // vC= 1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001111; // iC= 1167 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000010101111100; // vC= 1404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111000; // iC= 1080 
vC = 14'b0000010100100001; // vC= 1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000100; // iC= 1092 
vC = 14'b0000010110011111; // vC= 1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101010; // iC= 1066 
vC = 14'b0000010110111100; // vC= 1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001110110; // iC= 1142 
vC = 14'b0000010101110000; // vC= 1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000111110; // iC= 1086 
vC = 14'b0000010110101011; // vC= 1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001000; // iC= 1096 
vC = 14'b0000010110111001; // vC= 1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010111; // iC= 1047 
vC = 14'b0000010110010111; // vC= 1431 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000101; // iC= 1093 
vC = 14'b0000010101110001; // vC= 1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000110; // iC= 1094 
vC = 14'b0000010101011100; // vC= 1372 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100110; // iC= 1062 
vC = 14'b0000010101111011; // vC= 1403 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110010; // iC= 1010 
vC = 14'b0000010101101100; // vC= 1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010110; // iC= 1110 
vC = 14'b0000010110001100; // vC= 1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001000; // iC= 1032 
vC = 14'b0000010111010110; // vC= 1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000101; // iC= 1029 
vC = 14'b0000010110010011; // vC= 1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000000010; // iC= 1026 
vC = 14'b0000010101101110; // vC= 1390 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001100; // iC= 1036 
vC = 14'b0000010101001100; // vC= 1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001001111; // iC= 1103 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101101; // iC= 1005 
vC = 14'b0000010110101111; // vC= 1455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110111; // iC=  951 
vC = 14'b0000010111100101; // vC= 1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011000; // iC=  984 
vC = 14'b0000010110000000; // vC= 1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101010; // iC= 1066 
vC = 14'b0000010110000011; // vC= 1411 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000001001; // iC= 1033 
vC = 14'b0000010101110001; // vC= 1393 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000011111; // iC= 1055 
vC = 14'b0000010101110110; // vC= 1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111010010; // iC=  978 
vC = 14'b0000010101100110; // vC= 1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010111; // iC= 1047 
vC = 14'b0000010111001001; // vC= 1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111000; // iC=  952 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111100101; // iC=  997 
vC = 14'b0000010110111001; // vC= 1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011110; // iC=  926 
vC = 14'b0000010110001011; // vC= 1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001001; // iC=  905 
vC = 14'b0000010110001101; // vC= 1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110000; // iC=  944 
vC = 14'b0000010110111011; // vC= 1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101010; // iC=  938 
vC = 14'b0000010111000111; // vC= 1479 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111011; // iC=  955 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101101111; // iC=  879 
vC = 14'b0000010111110011; // vC= 1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110110001; // iC=  945 
vC = 14'b0000010111000000; // vC= 1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111101010; // iC= 1002 
vC = 14'b0000010111001001; // vC= 1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110111011; // iC=  955 
vC = 14'b0000011000001100; // vC= 1548 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000110; // iC=  838 
vC = 14'b0000010110100100; // vC= 1444 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010100; // iC=  916 
vC = 14'b0000010110101100; // vC= 1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110100; // iC=  884 
vC = 14'b0000010110100111; // vC= 1447 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101100101; // iC=  869 
vC = 14'b0000011000001101; // vC= 1549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111010; // iC=  890 
vC = 14'b0000010111001011; // vC= 1483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101110101; // iC=  885 
vC = 14'b0000011000101111; // vC= 1583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110100001; // iC=  929 
vC = 14'b0000010110110101; // vC= 1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110001011; // iC=  907 
vC = 14'b0000011000101000; // vC= 1576 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010010; // iC=  914 
vC = 14'b0000010110011101; // vC= 1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100011100; // iC=  796 
vC = 14'b0000010111110110; // vC= 1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101111100; // iC=  892 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000101; // iC=  773 
vC = 14'b0000011000010001; // vC= 1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000010; // iC=  898 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010001; // iC=  913 
vC = 14'b0000010110110110; // vC= 1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110101; // iC=  757 
vC = 14'b0000010111110111; // vC= 1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010000; // iC=  784 
vC = 14'b0000010111110010; // vC= 1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000111; // iC=  839 
vC = 14'b0000010111011010; // vC= 1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111110; // iC=  766 
vC = 14'b0000010111100100; // vC= 1508 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000111; // iC=  775 
vC = 14'b0000011000011001; // vC= 1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000100; // iC=  772 
vC = 14'b0000011000101001; // vC= 1577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100111110; // iC=  830 
vC = 14'b0000010111110011; // vC= 1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100101010; // iC=  810 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011111; // iC=  863 
vC = 14'b0000010111000000; // vC= 1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100100001; // iC=  801 
vC = 14'b0000010111010100; // vC= 1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000111; // iC=  775 
vC = 14'b0000010111101000; // vC= 1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011101; // iC=  733 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011110101; // iC=  757 
vC = 14'b0000011000001001; // vC= 1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000010; // iC=  706 
vC = 14'b0000010111111011; // vC= 1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101110; // iC=  750 
vC = 14'b0000010111010100; // vC= 1492 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001111; // iC=  719 
vC = 14'b0000011001100010; // vC= 1634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011111000; // iC=  760 
vC = 14'b0000011001010001; // vC= 1617 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100000001; // iC=  769 
vC = 14'b0000011000010100; // vC= 1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011011000; // iC=  728 
vC = 14'b0000011001001101; // vC= 1613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011101001; // iC=  745 
vC = 14'b0000011000000010; // vC= 1538 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010001100; // iC=  652 
vC = 14'b0000010111011100; // vC= 1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011000010; // iC=  706 
vC = 14'b0000011001001111; // vC= 1615 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010001; // iC=  785 
vC = 14'b0000010111100111; // vC= 1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100001011; // iC=  779 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001100; // iC=  716 
vC = 14'b0000011001111010; // vC= 1658 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100100; // iC=  612 
vC = 14'b0000010111100111; // vC= 1511 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100010; // iC=  738 
vC = 14'b0000010111100000; // vC= 1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100101; // iC=  741 
vC = 14'b0000010111011111; // vC= 1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001111010; // iC=  634 
vC = 14'b0000011001111011; // vC= 1659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101001; // iC=  617 
vC = 14'b0000010111111110; // vC= 1534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011010110; // iC=  726 
vC = 14'b0000011001111110; // vC= 1662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000010; // iC=  578 
vC = 14'b0000011001111110; // vC= 1662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001010; // iC=  586 
vC = 14'b0000011001110010; // vC= 1650 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000001; // iC=  577 
vC = 14'b0000011000010011; // vC= 1555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110110; // iC=  566 
vC = 14'b0000011001010101; // vC= 1621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000101111; // iC=  559 
vC = 14'b0000010111101110; // vC= 1518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100010; // iC=  546 
vC = 14'b0000010111111101; // vC= 1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010110100; // iC=  692 
vC = 14'b0000010111111010; // vC= 1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001001011; // iC=  587 
vC = 14'b0000011001001100; // vC= 1612 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100111; // iC=  679 
vC = 14'b0000010111110101; // vC= 1525 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100001; // iC=  673 
vC = 14'b0000011000000111; // vC= 1543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100111; // iC=  679 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001011110; // iC=  606 
vC = 14'b0000011000111010; // vC= 1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101000; // iC=  616 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010000111; // iC=  647 
vC = 14'b0000011001110100; // vC= 1652 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000111011; // iC=  571 
vC = 14'b0000011000001011; // vC= 1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101100; // iC=  492 
vC = 14'b0000011001101000; // vC= 1640 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101011; // iC=  619 
vC = 14'b0000011001011010; // vC= 1626 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000010001; // iC=  529 
vC = 14'b0000011010001110; // vC= 1678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100010; // iC=  482 
vC = 14'b0000011001000001; // vC= 1601 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111111001; // iC=  505 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011010; // iC=  474 
vC = 14'b0000011001010110; // vC= 1622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001000110; // iC=  582 
vC = 14'b0000011010001111; // vC= 1679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110101; // iC=  565 
vC = 14'b0000011010000101; // vC= 1669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111011; // iC=  443 
vC = 14'b0000011010011101; // vC= 1693 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011010; // iC=  538 
vC = 14'b0000011001001011; // vC= 1611 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110100; // iC=  564 
vC = 14'b0000011000110000; // vC= 1584 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101100; // iC=  492 
vC = 14'b0000011010000001; // vC= 1665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001000; // iC=  456 
vC = 14'b0000011001110001; // vC= 1649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000110000; // iC=  560 
vC = 14'b0000011001100110; // vC= 1638 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100011; // iC=  483 
vC = 14'b0000011010001001; // vC= 1673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111100; // iC=  444 
vC = 14'b0000011001101110; // vC= 1646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110011111; // iC=  415 
vC = 14'b0000011010000011; // vC= 1667 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111100111; // iC=  487 
vC = 14'b0000011010110001; // vC= 1713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111101001; // iC=  489 
vC = 14'b0000011010100010; // vC= 1698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111110; // iC=  446 
vC = 14'b0000011001100010; // vC= 1634 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111010011; // iC=  467 
vC = 14'b0000011001011000; // vC= 1624 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110111110; // iC=  446 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101100011; // iC=  355 
vC = 14'b0000011000011000; // vC= 1560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001001; // iC=  457 
vC = 14'b0000011001000100; // vC= 1604 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110001; // iC=  433 
vC = 14'b0000011001000000; // vC= 1600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110000000; // iC=  384 
vC = 14'b0000011010111001; // vC= 1721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111101; // iC=  317 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100111100; // iC=  316 
vC = 14'b0000011010101010; // vC= 1706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110010010; // iC=  402 
vC = 14'b0000011010011100; // vC= 1692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110000; // iC=  368 
vC = 14'b0000011001010010; // vC= 1618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101011010; // iC=  346 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001000; // iC=  328 
vC = 14'b0000011010111001; // vC= 1721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000001; // iC=  321 
vC = 14'b0000011010001000; // vC= 1672 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101001001; // iC=  329 
vC = 14'b0000011010100111; // vC= 1703 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100000010; // iC=  258 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011000100; // iC=  196 
vC = 14'b0000011010001101; // vC= 1677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010111100; // iC=  188 
vC = 14'b0000011010110011; // vC= 1715 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100010001; // iC=  273 
vC = 14'b0000011010100010; // vC= 1698 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011010011; // iC=  211 
vC = 14'b0000011011000000; // vC= 1728 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110000; // iC=  240 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011111110; // iC=  254 
vC = 14'b0000011001010011; // vC= 1619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011011110; // iC=  222 
vC = 14'b0000011001000111; // vC= 1607 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011011; // iC=   91 
vC = 14'b0000011000011111; // vC= 1567 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001001111; // iC=   79 
vC = 14'b0000011001011100; // vC= 1628 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001010; // iC=  138 
vC = 14'b0000011001011111; // vC= 1631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110010; // iC=   50 
vC = 14'b0000011000100101; // vC= 1573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111101; // iC=   61 
vC = 14'b0000011001101011; // vC= 1643 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001011111; // iC=   95 
vC = 14'b0000011010101110; // vC= 1710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001110101; // iC=  117 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111101; // iC=   61 
vC = 14'b0000011010011000; // vC= 1688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011111; // iC=   31 
vC = 14'b0000011001101111; // vC= 1647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101101; // iC=   45 
vC = 14'b0000011001101111; // vC= 1647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001010; // iC=  -54 
vC = 14'b0000011001000101; // vC= 1605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110100110; // iC=  -90 
vC = 14'b0000011001110000; // vC= 1648 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011001; // iC= -103 
vC = 14'b0000011000100001; // vC= 1569 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000001; // iC=  -63 
vC = 14'b0000011010000010; // vC= 1666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011111; // iC=  -97 
vC = 14'b0000011010001100; // vC= 1676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100111; // iC= -153 
vC = 14'b0000011001111110; // vC= 1662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110001; // iC= -143 
vC = 14'b0000011010101100; // vC= 1708 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000101; // iC=  -59 
vC = 14'b0000011010010101; // vC= 1685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100100; // iC= -156 
vC = 14'b0000011000101110; // vC= 1582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100110; // iC= -218 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101001000; // iC= -184 
vC = 14'b0000011010001001; // vC= 1673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100011; // iC= -157 
vC = 14'b0000011001001101; // vC= 1613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110011; // iC= -269 
vC = 14'b0000011010100000; // vC= 1696 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100011101; // iC= -227 
vC = 14'b0000011001100000; // vC= 1632 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100010; // iC= -350 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111000; // iC= -264 
vC = 14'b0000011001000010; // vC= 1602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011100010; // iC= -286 
vC = 14'b0000011000111110; // vC= 1598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011010101; // iC= -299 
vC = 14'b0000011010001110; // vC= 1678 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111000; // iC= -392 
vC = 14'b0000011000010101; // vC= 1557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000011; // iC= -381 
vC = 14'b0000011010000001; // vC= 1665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110010; // iC= -462 
vC = 14'b0000011000000000; // vC= 1536 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000011; // iC= -381 
vC = 14'b0000011000001010; // vC= 1546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000101100; // iC= -468 
vC = 14'b0000011010001100; // vC= 1676 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010011; // iC= -557 
vC = 14'b0000011000100010; // vC= 1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100011; // iC= -541 
vC = 14'b0000011010000001; // vC= 1665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111111; // iC= -577 
vC = 14'b0000011000111101; // vC= 1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101111; // iC= -529 
vC = 14'b0000010111111011; // vC= 1531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011111; // iC= -545 
vC = 14'b0000011010001111; // vC= 1679 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110100; // iC= -652 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111111; // iC= -641 
vC = 14'b0000011001111011; // vC= 1659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011011; // iC= -613 
vC = 14'b0000011001010000; // vC= 1616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110110; // iC= -586 
vC = 14'b0000011001111000; // vC= 1656 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110000111; // iC= -633 
vC = 14'b0000010111100001; // vC= 1505 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001000; // iC= -696 
vC = 14'b0000011000111101; // vC= 1597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001000; // iC= -760 
vC = 14'b0000011001001110; // vC= 1614 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101000; // iC= -728 
vC = 14'b0000011001101111; // vC= 1647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111010; // iC= -774 
vC = 14'b0000010111011011; // vC= 1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001111; // iC= -817 
vC = 14'b0000010111110010; // vC= 1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010011; // iC= -877 
vC = 14'b0000011000111011; // vC= 1595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111101; // iC= -899 
vC = 14'b0000010111001100; // vC= 1484 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101011; // iC= -853 
vC = 14'b0000011000010000; // vC= 1552 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001011; // iC= -885 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010111100; // iC= -836 
vC = 14'b0000010111110001; // vC= 1521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001000101; // iC= -955 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101010; // iC= -854 
vC = 14'b0000010111110000; // vC= 1520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111100; // iC= -900 
vC = 14'b0000010111101101; // vC= 1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110111; // iC= -905 
vC = 14'b0000011000001111; // vC= 1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010101; // iC= -939 
vC = 14'b0000011000011010; // vC= 1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001111; // iC= -945 
vC = 14'b0000011000011100; // vC= 1564 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100010; // iC= -990 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000110; // iC=-1082 
vC = 14'b0000010110110010; // vC= 1458 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010010; // iC=-1006 
vC = 14'b0000011000000101; // vC= 1541 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000101; // iC=-1083 
vC = 14'b0000010111100101; // vC= 1509 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110011011; // iC=-1125 
vC = 14'b0000011000011110; // vC= 1566 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110110; // iC=-1098 
vC = 14'b0000011000100100; // vC= 1572 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001001; // iC=-1143 
vC = 14'b0000010111110100; // vC= 1524 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111111; // iC=-1153 
vC = 14'b0000011000000011; // vC= 1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101110; // iC=-1106 
vC = 14'b0000011000001001; // vC= 1545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110001; // iC=-1103 
vC = 14'b0000010111010001; // vC= 1489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111011; // iC=-1221 
vC = 14'b0000010111111100; // vC= 1532 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110001001; // iC=-1143 
vC = 14'b0000010110010011; // vC= 1427 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111011; // iC=-1221 
vC = 14'b0000010110000001; // vC= 1409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101010; // iC=-1302 
vC = 14'b0000010110101110; // vC= 1454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100000; // iC=-1248 
vC = 14'b0000010110010010; // vC= 1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101011101; // iC=-1187 
vC = 14'b0000010111101001; // vC= 1513 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100011001; // iC=-1255 
vC = 14'b0000010101101100; // vC= 1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101111; // iC=-1361 
vC = 14'b0000010110010110; // vC= 1430 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111111; // iC=-1345 
vC = 14'b0000010110010010; // vC= 1426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000100; // iC=-1340 
vC = 14'b0000010101000100; // vC= 1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110111; // iC=-1417 
vC = 14'b0000010110011110; // vC= 1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001001; // iC=-1271 
vC = 14'b0000010110000111; // vC= 1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010100; // iC=-1388 
vC = 14'b0000010111000010; // vC= 1474 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010100; // iC=-1388 
vC = 14'b0000010101111000; // vC= 1400 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100111; // iC=-1433 
vC = 14'b0000010110100101; // vC= 1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b0000010101101100; // vC= 1388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010001011; // iC=-1397 
vC = 14'b0000010100111100; // vC= 1340 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111010; // iC=-1478 
vC = 14'b0000010101111110; // vC= 1406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110111; // iC=-1481 
vC = 14'b0000010100101000; // vC= 1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101001; // iC=-1431 
vC = 14'b0000010110000101; // vC= 1413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b0000010110101010; // vC= 1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111101; // iC=-1411 
vC = 14'b0000010100011110; // vC= 1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001100101; // iC=-1435 
vC = 14'b0000010101110000; // vC= 1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011110; // iC=-1506 
vC = 14'b0000010110001101; // vC= 1421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b0000010101100100; // vC= 1380 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110100; // iC=-1548 
vC = 14'b0000010100010010; // vC= 1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b0000010100100001; // vC= 1313 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111101; // iC=-1603 
vC = 14'b0000010100110010; // vC= 1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001010100; // iC=-1452 
vC = 14'b0000010100001011; // vC= 1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101100; // iC=-1556 
vC = 14'b0000010100100010; // vC= 1314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100100; // iC=-1500 
vC = 14'b0000010101000111; // vC= 1351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b0000010101010100; // vC= 1364 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b0000010100011110; // vC= 1310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010111; // iC=-1577 
vC = 14'b0000010100001100; // vC= 1292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011001; // iC=-1575 
vC = 14'b0000010011111001; // vC= 1273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011110; // iC=-1634 
vC = 14'b0000010011101010; // vC= 1258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b0000010010101011; // vC= 1195 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010011; // iC=-1645 
vC = 14'b0000010011011101; // vC= 1245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101011; // iC=-1557 
vC = 14'b0000010011000000; // vC= 1216 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101011; // iC=-1621 
vC = 14'b0000010011100010; // vC= 1250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000010; // iC=-1662 
vC = 14'b0000010011001011; // vC= 1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011101; // iC=-1635 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b0000010010100011; // vC= 1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000110; // iC=-1594 
vC = 14'b0000010010111010; // vC= 1210 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100011; // iC=-1629 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011000; // iC=-1704 
vC = 14'b0000010001101010; // vC= 1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100000; // iC=-1632 
vC = 14'b0000010001100101; // vC= 1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b0000010011011110; // vC= 1246 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b0000010001100111; // vC= 1127 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000011; // iC=-1725 
vC = 14'b0000010010101111; // vC= 1199 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b0000010010111111; // vC= 1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b0000010010000110; // vC= 1158 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000110; // iC=-1658 
vC = 14'b0000010001110101; // vC= 1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110111; // iC=-1609 
vC = 14'b0000010011000110; // vC= 1222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b0000010001011100; // vC= 1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011001; // iC=-1639 
vC = 14'b0000010010100001; // vC= 1185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000010000011101; // vC= 1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b0000010001001110; // vC= 1102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000010000110110; // vC= 1078 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010010; // iC=-1646 
vC = 14'b0000010010000010; // vC= 1154 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b0000010001110001; // vC= 1137 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000010001011010; // vC= 1114 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011110; // iC=-1698 
vC = 14'b0000010010001011; // vC= 1163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b0000010010000011; // vC= 1155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111011; // iC=-1669 
vC = 14'b0000010001011100; // vC= 1116 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000100; // iC=-1724 
vC = 14'b0000010000001000; // vC= 1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010010; // iC=-1710 
vC = 14'b0000010001001011; // vC= 1099 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101011; // iC=-1685 
vC = 14'b0000010001000110; // vC= 1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001000; // iC=-1784 
vC = 14'b0000010000011101; // vC= 1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111010; // iC=-1734 
vC = 14'b0000010000111011; // vC= 1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b0000010001001101; // vC= 1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000001111100100; // vC=  996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011110; // iC=-1698 
vC = 14'b0000010000001100; // vC= 1036 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b0000010000011101; // vC= 1053 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010000; // iC=-1712 
vC = 14'b0000001110101100; // vC=  940 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000001110010110; // vC=  918 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100001; // iC=-1695 
vC = 14'b0000001110100100; // vC=  932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011000; // iC=-1768 
vC = 14'b0000001111001000; // vC=  968 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000001110100111; // vC=  935 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000101; // iC=-1659 
vC = 14'b0000001110101001; // vC=  937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100001; // iC=-1759 
vC = 14'b0000001111010001; // vC=  977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b0000001111100111; // vC=  999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100010; // iC=-1694 
vC = 14'b0000001110101000; // vC=  936 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110101; // iC=-1803 
vC = 14'b0000001111110110; // vC= 1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011100; // iC=-1700 
vC = 14'b0000001111110011; // vC= 1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011011; // iC=-1701 
vC = 14'b0000001111010001; // vC=  977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000001101010110; // vC=  854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b0000001101010100; // vC=  852 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b0000001101100011; // vC=  867 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100111; // iC=-1817 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000001100110111; // vC=  823 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000001; // iC=-1791 
vC = 14'b0000001111000100; // vC=  964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010011; // iC=-1837 
vC = 14'b0000001110001010; // vC=  906 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b0000001100101111; // vC=  815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101111; // iC=-1809 
vC = 14'b0000001110010100; // vC=  916 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000001100010011; // vC=  787 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101011; // iC=-1813 
vC = 14'b0000001101110001; // vC=  881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000001101100110; // vC=  870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000001110001001; // vC=  905 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110010; // iC=-1742 
vC = 14'b0000001100010010; // vC=  786 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b0000001100001001; // vC=  777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101001; // iC=-1815 
vC = 14'b0000001100001001; // vC=  777 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000101; // iC=-1787 
vC = 14'b0000001101000100; // vC=  836 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000001011110110; // vC=  758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101100; // iC=-1748 
vC = 14'b0000001011001110; // vC=  718 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000011; // iC=-1853 
vC = 14'b0000001100111101; // vC=  829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001111; // iC=-1713 
vC = 14'b0000001101000110; // vC=  838 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010100; // iC=-1836 
vC = 14'b0000001100010001; // vC=  785 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000001100000000; // vC=  768 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000001010111101; // vC=  701 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111101; // iC=-1859 
vC = 14'b0000001010111110; // vC=  702 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011110; // iC=-1826 
vC = 14'b0000001100001011; // vC=  779 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000001100011110; // vC=  798 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000010; // iC=-1726 
vC = 14'b0000001011001111; // vC=  719 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010100; // iC=-1836 
vC = 14'b0000001011011011; // vC=  731 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b0000001010001111; // vC=  655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000001011110100; // vC=  756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000001011000011; // vC=  707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000001011000111; // vC=  711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000001001110111; // vC=  631 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000001010101000; // vC=  680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000001011001001; // vC=  713 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000001011001000; // vC=  712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010010; // iC=-1838 
vC = 14'b0000001001100101; // vC=  613 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000001010010100; // vC=  660 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001110; // iC=-1842 
vC = 14'b0000001001010101; // vC=  597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001101; // iC=-1843 
vC = 14'b0000001001000110; // vC=  582 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000100; // iC=-1724 
vC = 14'b0000001000101010; // vC=  554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000001001001010; // vC=  586 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001100; // iC=-1780 
vC = 14'b0000001000011110; // vC=  542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001110; // iC=-1842 
vC = 14'b0000001001011011; // vC=  603 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110101; // iC=-1739 
vC = 14'b0000001001010100; // vC=  596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011001; // iC=-1831 
vC = 14'b0000001010000111; // vC=  647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000001000001001; // vC=  521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111001; // iC=-1735 
vC = 14'b0000001001100001; // vC=  609 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101101; // iC=-1875 
vC = 14'b0000001000101001; // vC=  553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101011; // iC=-1877 
vC = 14'b0000001000101101; // vC=  557 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100000; // iC=-1824 
vC = 14'b0000001000101011; // vC=  555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000000111111010; // vC=  506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000000111110100; // vC=  500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001111; // iC=-1777 
vC = 14'b0000001001101011; // vC=  619 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111111; // iC=-1857 
vC = 14'b0000000111111000; // vC=  504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000001000101011; // vC=  555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101011; // iC=-1749 
vC = 14'b0000001000011100; // vC=  540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011010; // iC=-1766 
vC = 14'b0000000111101110; // vC=  494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000010; // iC=-1854 
vC = 14'b0000000111110010; // vC=  498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111011; // iC=-1861 
vC = 14'b0000000111110010; // vC=  498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b0000000110111011; // vC=  443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100101; // iC=-1819 
vC = 14'b0000000110100011; // vC=  419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111111; // iC=-1793 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100111; // iC=-1881 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000001000100101; // vC=  549 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100110; // iC=-1818 
vC = 14'b0000001000000100; // vC=  516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010001; // iC=-1775 
vC = 14'b0000000111101000; // vC=  488 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000000110000111; // vC=  391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000000110010110; // vC=  406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000000110000100; // vC=  388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000000110111010; // vC=  442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110110; // iC=-1802 
vC = 14'b0000000111100110; // vC=  486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001010; // iC=-1846 
vC = 14'b0000000111000110; // vC=  454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111011; // iC=-1733 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101110; // iC=-1810 
vC = 14'b0000000110011001; // vC=  409 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000000101010110; // vC=  342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000000101100110; // vC=  358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010001; // iC=-1839 
vC = 14'b0000000111001111; // vC=  463 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010100001; // iC=-1887 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110001; // iC=-1743 
vC = 14'b0000000100101000; // vC=  296 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000000110000010; // vC=  386 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b0000000110111000; // vC=  440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010011100; // iC=-1892 
vC = 14'b0000000100101001; // vC=  297 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010100; // iC=-1836 
vC = 14'b0000000100010010; // vC=  274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000000101101010; // vC=  362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000000100100101; // vC=  293 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111101; // iC=-1731 
vC = 14'b0000000011111000; // vC=  248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000110; // iC=-1850 
vC = 14'b0000000100001001; // vC=  265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b0000000100100100; // vC=  292 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011011101; // iC=-1827 
vC = 14'b0000000011101101; // vC=  237 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000110; // iC=-1786 
vC = 14'b0000000100111100; // vC=  316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000100; // iC=-1852 
vC = 14'b0000000011101100; // vC=  236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000101; // iC=-1851 
vC = 14'b0000000100100010; // vC=  290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111000; // iC=-1864 
vC = 14'b0000000011011110; // vC=  222 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110001; // iC=-1871 
vC = 14'b0000000011110101; // vC=  245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011010110; // iC=-1834 
vC = 14'b0000000100110100; // vC=  308 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110011; // iC=-1741 
vC = 14'b0000000011110100; // vC=  244 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101111; // iC=-1873 
vC = 14'b0000000010110110; // vC=  182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000000100010111; // vC=  279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111011; // iC=-1861 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000010; // iC=-1790 
vC = 14'b0000000010111100; // vC=  188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000000011111100; // vC=  252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000000010111100; // vC=  188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110001; // iC=-1807 
vC = 14'b0000000011001101; // vC=  205 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010111; // iC=-1769 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010101000; // iC=-1880 
vC = 14'b0000000011011101; // vC=  221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100000; // iC=-1824 
vC = 14'b0000000010100010; // vC=  162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101000; // iC=-1752 
vC = 14'b0000000011011001; // vC=  217 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000000; // iC=-1728 
vC = 14'b0000000010010000; // vC=  144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101001; // iC=-1751 
vC = 14'b0000000011001110; // vC=  206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000000; // iC=-1792 
vC = 14'b0000000001110000; // vC=  112 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111101; // iC=-1795 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000000010110011; // vC=  179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000000011000110; // vC=  198 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b0000000001000000; // vC=   64 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010110110; // iC=-1866 
vC = 14'b0000000010011100; // vC=  156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b0000000010100011; // vC=  163 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011101; // iC=-1763 
vC = 14'b0000000000101101; // vC=   45 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000111; // iC=-1785 
vC = 14'b0000000001101010; // vC=  106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000100; // iC=-1788 
vC = 14'b0000000010101110; // vC=  174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110100; // iC=-1804 
vC = 14'b0000000010100000; // vC=  160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011000001; // iC=-1855 
vC = 14'b0000000000001101; // vC=   13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111101; // iC=-1859 
vC = 14'b0000000010100001; // vC=  161 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110000; // iC=-1744 
vC = 14'b0000000000000001; // vC=    1 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b0000000001010001; // vC=   81 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100010111100; // iC=-1860 
vC = 14'b0000000010000000; // vC=  128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001001; // iC=-1847 
vC = 14'b0000000000011111; // vC=   31 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000110; // iC=-1722 
vC = 14'b1111111111100010; // vC=  -30 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001000; // iC=-1848 
vC = 14'b0000000000110010; // vC=   50 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000000000100101; // vC=   37 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b0000000001010000; // vC=   80 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b0000000000101110; // vC=   46 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101110; // iC=-1746 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011101100; // iC=-1812 
vC = 14'b1111111111110101; // vC=  -11 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b0000000001001011; // vC=   75 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b0000000001000100; // vC=   68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001110; // iC=-1714 
vC = 14'b0000000001001000; // vC=   72 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000101; // iC=-1723 
vC = 14'b1111111111000110; // vC=  -58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b1111111110011011; // vC= -101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011111; // iC=-1761 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100101111; // iC=-1745 
vC = 14'b1111111111010001; // vC=  -47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b1111111110011110; // vC=  -98 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011001010; // iC=-1846 
vC = 14'b0000000000001100; // vC=   12 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b1111111111011000; // vC=  -40 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110011; // iC=-1805 
vC = 14'b1111111110011000; // vC= -104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001000; // iC=-1720 
vC = 14'b1111111110001000; // vC= -120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b1111111110000110; // vC= -122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100001101; // iC=-1779 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b1111111110111101; // vC=  -67 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011110000; // iC=-1808 
vC = 14'b1111111101001100; // vC= -180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100011; // iC=-1757 
vC = 14'b1111111111010001; // vC=  -47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111110; // iC=-1794 
vC = 14'b1111111101001101; // vC= -179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000111; // iC=-1721 
vC = 14'b1111111101010011; // vC= -173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011100010; // iC=-1822 
vC = 14'b1111111101110101; // vC= -139 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011011; // iC=-1765 
vC = 14'b1111111110011101; // vC=  -99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111111; // iC=-1729 
vC = 14'b1111111110100001; // vC=  -95 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b1111111100110010; // vC= -206 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101101; // iC=-1683 
vC = 14'b1111111101101101; // vC= -147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100011111100; // iC=-1796 
vC = 14'b1111111101000000; // vC= -192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001001; // iC=-1719 
vC = 14'b1111111110011101; // vC=  -99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b1111111101000001; // vC= -191 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101000001; // iC=-1727 
vC = 14'b1111111101110100; // vC= -140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100100111; // iC=-1753 
vC = 14'b1111111101100000; // vC= -160 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010100; // iC=-1772 
vC = 14'b1111111101111111; // vC= -129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100000011; // iC=-1789 
vC = 14'b1111111011101101; // vC= -275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001010; // iC=-1718 
vC = 14'b1111111110000110; // vC= -122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100011001; // iC=-1767 
vC = 14'b1111111011111110; // vC= -258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110011; // iC=-1677 
vC = 14'b1111111100000110; // vC= -250 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101111; // iC=-1681 
vC = 14'b1111111011010011; // vC= -301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100000; // iC=-1696 
vC = 14'b1111111011111110; // vC= -258 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100101; // iC=-1691 
vC = 14'b1111111011110010; // vC= -270 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011111; // iC=-1697 
vC = 14'b1111111100111110; // vC= -194 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010110; // iC=-1770 
vC = 14'b1111111011000101; // vC= -315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b1111111100001011; // vC= -245 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000000; // iC=-1664 
vC = 14'b1111111100100100; // vC= -220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100100; // iC=-1692 
vC = 14'b1111111100100101; // vC= -219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b1111111010110101; // vC= -331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b1111111100000000; // vC= -256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b1111111011101001; // vC= -279 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010001; // iC=-1711 
vC = 14'b1111111010010000; // vC= -368 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101100110; // iC=-1690 
vC = 14'b1111111011010011; // vC= -301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100010000; // iC=-1776 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110101011; // iC=-1621 
vC = 14'b1111111011111001; // vC= -263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010101; // iC=-1707 
vC = 14'b1111111010000110; // vC= -378 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011110; // iC=-1698 
vC = 14'b1111111010000000; // vC= -384 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100110110; // iC=-1738 
vC = 14'b1111111011000010; // vC= -318 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100100; // iC=-1628 
vC = 14'b1111111001111101; // vC= -387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110000; // iC=-1616 
vC = 14'b1111111010010101; // vC= -363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111010; // iC=-1606 
vC = 14'b1111111011000100; // vC= -316 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111011; // iC=-1605 
vC = 14'b1111111010101010; // vC= -342 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100010; // iC=-1630 
vC = 14'b1111111010101001; // vC= -343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100100111100; // iC=-1732 
vC = 14'b1111111010111110; // vC= -322 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101111000; // iC=-1672 
vC = 14'b1111111010000010; // vC= -382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011010; // iC=-1638 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001011; // iC=-1653 
vC = 14'b1111111011001010; // vC= -310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110100; // iC=-1676 
vC = 14'b1111111010011010; // vC= -358 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100101; // iC=-1627 
vC = 14'b1111111010100001; // vC= -351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101011001; // iC=-1703 
vC = 14'b1111111010010011; // vC= -365 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001011; // iC=-1717 
vC = 14'b1111111001000110; // vC= -442 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101110010; // iC=-1678 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101010111; // iC=-1705 
vC = 14'b1111111001000000; // vC= -448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100001; // iC=-1631 
vC = 14'b1111111001001001; // vC= -439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101001; // iC=-1687 
vC = 14'b1111111000111001; // vC= -455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110010100; // iC=-1644 
vC = 14'b1111111010000011; // vC= -381 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101001100; // iC=-1716 
vC = 14'b1111111001110110; // vC= -394 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b1111111001110010; // vC= -398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011101; // iC=-1571 
vC = 14'b1111111001000011; // vC= -445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010111; // iC=-1577 
vC = 14'b1111111000111001; // vC= -455 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100111; // iC=-1625 
vC = 14'b1111111001011101; // vC= -419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000111; // iC=-1593 
vC = 14'b1111111001101011; // vC= -405 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110001100; // iC=-1652 
vC = 14'b1111110111111101; // vC= -515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111100; // iC=-1540 
vC = 14'b1111110111110000; // vC= -528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110001; // iC=-1615 
vC = 14'b1111111001001101; // vC= -435 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100010; // iC=-1566 
vC = 14'b1111110111011111; // vC= -545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000010; // iC=-1662 
vC = 14'b1111111000000000; // vC= -512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011111; // iC=-1569 
vC = 14'b1111111001001111; // vC= -433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110000111; // iC=-1657 
vC = 14'b1111111000111010; // vC= -454 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100101101100; // iC=-1684 
vC = 14'b1111110110110101; // vC= -587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000000; // iC=-1600 
vC = 14'b1111110110110000; // vC= -592 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000101; // iC=-1531 
vC = 14'b1111110111010010; // vC= -558 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001111; // iC=-1585 
vC = 14'b1111110110111001; // vC= -583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110100; // iC=-1612 
vC = 14'b1111110110101110; // vC= -594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110111111; // iC=-1601 
vC = 14'b1111110111111100; // vC= -516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110011111; // iC=-1633 
vC = 14'b1111110110011110; // vC= -610 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111000; // iC=-1544 
vC = 14'b1111110111111010; // vC= -518 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111001; // iC=-1543 
vC = 14'b1111110110010010; // vC= -622 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b1111111000010011; // vC= -493 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010010; // iC=-1582 
vC = 14'b1111111000001111; // vC= -497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101011; // iC=-1557 
vC = 14'b1111110110100110; // vC= -602 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110110010; // iC=-1614 
vC = 14'b1111110111011001; // vC= -551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100110100110; // iC=-1626 
vC = 14'b1111110110010110; // vC= -618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111110010; // iC=-1550 
vC = 14'b1111110111111000; // vC= -520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000011; // iC=-1597 
vC = 14'b1111110111010101; // vC= -555 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111010; // iC=-1542 
vC = 14'b1111110111011110; // vC= -546 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001101; // iC=-1587 
vC = 14'b1111110110100011; // vC= -605 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101001; // iC=-1559 
vC = 14'b1111110101100100; // vC= -668 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101010; // iC=-1494 
vC = 14'b1111110110101101; // vC= -595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001110; // iC=-1586 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001001101; // iC=-1459 
vC = 14'b1111110101101101; // vC= -659 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b1111110101101011; // vC= -661 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111111111; // iC=-1537 
vC = 14'b1111110101111010; // vC= -646 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b1111110101111011; // vC= -645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111001000; // iC=-1592 
vC = 14'b1111110110000011; // vC= -637 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000001; // iC=-1471 
vC = 14'b1111110101111001; // vC= -647 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000101100; // iC=-1492 
vC = 14'b1111110101011011; // vC= -677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111000100; // iC=-1596 
vC = 14'b1111110101011111; // vC= -673 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000110; // iC=-1530 
vC = 14'b1111110101001010; // vC= -694 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000010; // iC=-1470 
vC = 14'b1111110101001100; // vC= -692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111010010; // iC=-1582 
vC = 14'b1111110011111110; // vC= -770 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111100111; // iC=-1561 
vC = 14'b1111110100000010; // vC= -766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011110; // iC=-1442 
vC = 14'b1111110100111101; // vC= -707 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001011; // iC=-1525 
vC = 14'b1111110101111100; // vC= -644 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111011110; // iC=-1570 
vC = 14'b1111110011100101; // vC= -795 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001001; // iC=-1527 
vC = 14'b1111110101011011; // vC= -677 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110011; // iC=-1485 
vC = 14'b1111110101011101; // vC= -675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111100111101000; // iC=-1560 
vC = 14'b1111110100110100; // vC= -716 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000011; // iC=-1405 
vC = 14'b1111110011010111; // vC= -809 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001000110; // iC=-1466 
vC = 14'b1111110011100011; // vC= -797 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000000001; // iC=-1535 
vC = 14'b1111110011011110; // vC= -802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000100110; // iC=-1498 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000011011; // iC=-1509 
vC = 14'b1111110011011110; // vC= -802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000001110; // iC=-1522 
vC = 14'b1111110011011010; // vC= -806 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000100; // iC=-1404 
vC = 14'b1111110011001110; // vC= -818 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010110; // iC=-1514 
vC = 14'b1111110100111010; // vC= -710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000010111; // iC=-1513 
vC = 14'b1111110011010001; // vC= -815 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b1111110100100010; // vC= -734 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000110001; // iC=-1487 
vC = 14'b1111110100101111; // vC= -721 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011000; // iC=-1384 
vC = 14'b1111110010011001; // vC= -871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001111110; // iC=-1410 
vC = 14'b1111110100010011; // vC= -749 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011101; // iC=-1379 
vC = 14'b1111110010110010; // vC= -846 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010101110; // iC=-1362 
vC = 14'b1111110011100000; // vC= -800 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011100; // iC=-1380 
vC = 14'b1111110011011001; // vC= -807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101000111000; // iC=-1480 
vC = 14'b1111110010100001; // vC= -863 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011011; // iC=-1381 
vC = 14'b1111110010010100; // vC= -876 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111110011000001; // vC= -831 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001101; // iC=-1331 
vC = 14'b1111110010101001; // vC= -855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011010; // iC=-1382 
vC = 14'b1111110010000010; // vC= -894 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010011101; // iC=-1379 
vC = 14'b1111110011000101; // vC= -827 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101000; // iC=-1432 
vC = 14'b1111110011010010; // vC= -814 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000111; // iC=-1401 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101000; // iC=-1432 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001011010; // iC=-1446 
vC = 14'b1111110011010000; // vC= -816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001001; // iC=-1335 
vC = 14'b1111110001000111; // vC= -953 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b1111110011001010; // vC= -822 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001110; // iC=-1330 
vC = 14'b1111110010010000; // vC= -880 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101101; // iC=-1427 
vC = 14'b1111110001110001; // vC= -911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001101; // iC=-1331 
vC = 14'b1111110001011110; // vC= -930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001110001; // iC=-1423 
vC = 14'b1111110001110010; // vC= -910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101001101111; // iC=-1425 
vC = 14'b1111110010011001; // vC= -871 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110110; // iC=-1290 
vC = 14'b1111110010011011; // vC= -869 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010011; // iC=-1389 
vC = 14'b1111110010010110; // vC= -874 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101110; // iC=-1298 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111011; // iC=-1349 
vC = 14'b1111110000100101; // vC= -987 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010010100; // iC=-1388 
vC = 14'b1111110000100010; // vC= -990 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101010; // iC=-1302 
vC = 14'b1111110000110000; // vC= -976 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010000101; // iC=-1403 
vC = 14'b1111110001110011; // vC= -909 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101000; // iC=-1304 
vC = 14'b1111110001111000; // vC= -904 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010110010; // iC=-1358 
vC = 14'b1111110000000100; // vC=-1020 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011110001; // iC=-1295 
vC = 14'b1111110001000110; // vC= -954 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000001; // iC=-1279 
vC = 14'b1111110001110010; // vC= -910 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011010001; // iC=-1327 
vC = 14'b1111110000010010; // vC=-1006 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010100100; // iC=-1372 
vC = 14'b1111110001011100; // vC= -932 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011000110; // iC=-1338 
vC = 14'b1111110000100011; // vC= -989 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111110; // iC=-1282 
vC = 14'b1111110000010000; // vC=-1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100001110; // iC=-1266 
vC = 14'b1111110000101001; // vC= -983 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000110; // iC=-1274 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011001001; // iC=-1335 
vC = 14'b1111101111111000; // vC=-1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001111; // iC=-1201 
vC = 14'b1111110001100001; // vC= -927 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111101; // iC=-1283 
vC = 14'b1111110000111010; // vC= -966 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010111; // iC=-1257 
vC = 14'b1111110000011001; // vC= -999 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101010111110; // iC=-1346 
vC = 14'b1111101111011100; // vC=-1060 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b1111110000001111; // vC=-1009 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110010; // iC=-1230 
vC = 14'b1111101111100110; // vC=-1050 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101010; // iC=-1238 
vC = 14'b1111110000001101; // vC=-1011 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101001010; // iC=-1206 
vC = 14'b1111110001000001; // vC= -959 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100101010; // iC=-1238 
vC = 14'b1111110000001000; // vC=-1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011111000; // iC=-1288 
vC = 14'b1111110001001000; // vC= -952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101011101110; // iC=-1298 
vC = 14'b1111101111111001; // vC=-1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100000000; // iC=-1280 
vC = 14'b1111110000010011; // vC=-1005 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010011; // iC=-1197 
vC = 14'b1111101111111000; // vC=-1032 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100111100; // iC=-1220 
vC = 14'b1111101110100101; // vC=-1115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100110; // iC=-1242 
vC = 14'b1111101111100111; // vC=-1049 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100010100; // iC=-1260 
vC = 14'b1111110000000111; // vC=-1017 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110010; // iC=-1166 
vC = 14'b1111101110110011; // vC=-1101 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100010; // iC=-1246 
vC = 14'b1111110000010001; // vC=-1007 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100100100; // iC=-1244 
vC = 14'b1111101111011000; // vC=-1064 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000000; // iC=-1152 
vC = 14'b1111101110011011; // vC=-1125 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010000; // iC=-1200 
vC = 14'b1111101111111001; // vC=-1031 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101110110; // iC=-1162 
vC = 14'b1111101110110000; // vC=-1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100101; // iC=-1179 
vC = 14'b1111101101111100; // vC=-1156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110101011; // iC=-1109 
vC = 14'b1111101111010111; // vC=-1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110111; // iC=-1225 
vC = 14'b1111101110111100; // vC=-1092 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100000; // iC=-1184 
vC = 14'b1111101110011101; // vC=-1123 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101100110001; // iC=-1231 
vC = 14'b1111101110010001; // vC=-1135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110111100; // iC=-1092 
vC = 14'b1111101111001000; // vC=-1080 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000011; // iC=-1085 
vC = 14'b1111101101111001; // vC=-1159 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110111; // iC=-1097 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101010100; // iC=-1196 
vC = 14'b1111101110011100; // vC=-1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111001110; // iC=-1074 
vC = 14'b1111101101011101; // vC=-1187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111010000; // iC=-1072 
vC = 14'b1111101110100010; // vC=-1118 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110010011; // iC=-1133 
vC = 14'b1111101111000000; // vC=-1088 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100000; // iC=-1184 
vC = 14'b1111101110011111; // vC=-1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110000000; // iC=-1152 
vC = 14'b1111101101100000; // vC=-1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101111001; // iC=-1159 
vC = 14'b1111101101000111; // vC=-1209 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110100; // iC=-1100 
vC = 14'b1111101111001110; // vC=-1074 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101101100011; // iC=-1181 
vC = 14'b1111101110000100; // vC=-1148 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111000; // iC=-1032 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000100; // iC=-1084 
vC = 14'b1111101101101000; // vC=-1176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100110; // iC=-1050 
vC = 14'b1111101100110001; // vC=-1231 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001001; // iC=-1015 
vC = 14'b1111101101010111; // vC=-1193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000101; // iC=-1019 
vC = 14'b1111101101101010; // vC=-1174 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111000; // iC=-1032 
vC = 14'b1111101110000010; // vC=-1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000001; // iC=-1087 
vC = 14'b1111101101010100; // vC=-1196 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111101101; // iC=-1043 
vC = 14'b1111101101110001; // vC=-1167 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100111; // iC=-1049 
vC = 14'b1111101110101100; // vC=-1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100011; // iC=-1053 
vC = 14'b1111101101101101; // vC=-1171 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111111011; // iC=-1029 
vC = 14'b1111101110000001; // vC=-1151 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001001; // iC=-1015 
vC = 14'b1111101110010110; // vC=-1130 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111000111; // iC=-1081 
vC = 14'b1111101100000110; // vC=-1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101110110000; // iC=-1104 
vC = 14'b1111101100100110; // vC=-1242 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000000111; // iC=-1017 
vC = 14'b1111101100010111; // vC=-1257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111011110; // iC=-1058 
vC = 14'b1111101100001000; // vC=-1272 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000010111; // iC=-1001 
vC = 14'b1111101101111011; // vC=-1157 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010100; // iC= -940 
vC = 14'b1111101101101011; // vC=-1173 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b1111101011111100; // vC=-1284 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111100100; // iC=-1052 
vC = 14'b1111101101000011; // vC=-1213 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011011; // iC= -933 
vC = 14'b1111101101011000; // vC=-1192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001101010; // iC= -918 
vC = 14'b1111101101000101; // vC=-1211 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100101; // iC= -987 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110100; // iC=-1036 
vC = 14'b1111101011111110; // vC=-1282 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111101111110000; // iC=-1040 
vC = 14'b1111101100001100; // vC=-1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001110010; // iC= -910 
vC = 14'b1111101101101111; // vC=-1169 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000100; // iC= -892 
vC = 14'b1111101011100111; // vC=-1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011000; // iC= -936 
vC = 14'b1111101101100000; // vC=-1184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100000; // iC= -992 
vC = 14'b1111101011000110; // vC=-1338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101101; // iC= -979 
vC = 14'b1111101011011011; // vC=-1317 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010110; // iC= -938 
vC = 14'b1111101011101101; // vC=-1299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000001110; // iC=-1010 
vC = 14'b1111101101000010; // vC=-1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010010; // iC= -942 
vC = 14'b1111101010111010; // vC=-1350 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010001001; // iC= -887 
vC = 14'b1111101011011101; // vC=-1315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001001000; // iC= -952 
vC = 14'b1111101100011100; // vC=-1252 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010000011; // iC= -893 
vC = 14'b1111101011101101; // vC=-1299 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000101110; // iC= -978 
vC = 14'b1111101100101100; // vC=-1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000100001; // iC= -991 
vC = 14'b1111101100111101; // vC=-1219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110000110110; // iC= -970 
vC = 14'b1111101100011111; // vC=-1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010010000; // iC= -880 
vC = 14'b1111101100001100; // vC=-1268 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001011110; // iC= -930 
vC = 14'b1111101011110111; // vC=-1289 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010101011; // iC= -853 
vC = 14'b1111101011001000; // vC=-1336 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011101; // iC= -867 
vC = 14'b1111101011100101; // vC=-1307 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110001; // iC= -847 
vC = 14'b1111101100000110; // vC=-1274 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001100110; // iC= -922 
vC = 14'b1111101100011000; // vC=-1256 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010110001; // iC= -847 
vC = 14'b1111101011110101; // vC=-1291 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001010; // iC= -822 
vC = 14'b1111101010010000; // vC=-1392 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001010100; // iC= -940 
vC = 14'b1111101100100000; // vC=-1248 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011001110; // iC= -818 
vC = 14'b1111101100000000; // vC=-1280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011010111; // iC= -809 
vC = 14'b1111101011101110; // vC=-1298 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010011111; // iC= -865 
vC = 14'b1111101011010100; // vC=-1324 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110001111001; // iC= -903 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011000; // iC= -808 
vC = 14'b1111101011100111; // vC=-1305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000100; // iC= -764 
vC = 14'b1111101011000111; // vC=-1337 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011111101; // iC= -771 
vC = 14'b1111101011110110; // vC=-1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010001; // iC= -751 
vC = 14'b1111101010111101; // vC=-1347 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000111; // iC= -761 
vC = 14'b1111101010010101; // vC=-1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100110; // iC= -858 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110010100010; // iC= -862 
vC = 14'b1111101011011000; // vC=-1320 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100110; // iC= -794 
vC = 14'b1111101011111011; // vC=-1285 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110001; // iC= -783 
vC = 14'b1111101001100001; // vC=-1439 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011110; // iC= -738 
vC = 14'b1111101001110101; // vC=-1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011101000; // iC= -792 
vC = 14'b1111101010001010; // vC=-1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011011; // iC= -805 
vC = 14'b1111101001110101; // vC=-1419 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010000; // iC= -752 
vC = 14'b1111101001110010; // vC=-1422 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000110; // iC= -762 
vC = 14'b1111101010111110; // vC=-1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011110111; // iC= -777 
vC = 14'b1111101010110000; // vC=-1360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011011001; // iC= -807 
vC = 14'b1111101011101100; // vC=-1300 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100001101; // iC= -755 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101001000; // iC= -696 
vC = 14'b1111101001100110; // vC=-1434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100010001; // iC= -751 
vC = 14'b1111101011001101; // vC=-1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011010; // iC= -678 
vC = 14'b1111101010111100; // vC=-1348 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100101001; // iC= -727 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100100110; // iC= -730 
vC = 14'b1111101011001110; // vC=-1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110011100111; // iC= -793 
vC = 14'b1111101001100100; // vC=-1436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110111; // iC= -713 
vC = 14'b1111101010001010; // vC=-1398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100000101; // iC= -763 
vC = 14'b1111101011001101; // vC=-1331 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101011011; // iC= -677 
vC = 14'b1111101010111110; // vC=-1346 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100011; // iC= -669 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001000; // iC= -632 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010110; // iC= -682 
vC = 14'b1111101001001011; // vC=-1461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100110101; // iC= -715 
vC = 14'b1111101010010101; // vC=-1387 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101101111; // iC= -657 
vC = 14'b1111101010110111; // vC=-1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111111; // iC= -641 
vC = 14'b1111101011000001; // vC=-1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110100011111; // iC= -737 
vC = 14'b1111101010100001; // vC=-1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001100; // iC= -628 
vC = 14'b1111101010100001; // vC=-1375 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001011; // iC= -629 
vC = 14'b1111101000101101; // vC=-1491 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110101011; // iC= -597 
vC = 14'b1111101000110011; // vC=-1485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111011; // iC= -645 
vC = 14'b1111101010010001; // vC=-1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101010101; // iC= -683 
vC = 14'b1111101001000011; // vC=-1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011000; // iC= -552 
vC = 14'b1111101000011101; // vC=-1507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110011101; // iC= -611 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101100010; // iC= -670 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101110010; // iC= -654 
vC = 14'b1111101001011010; // vC=-1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010000; // iC= -560 
vC = 14'b1111101001101000; // vC=-1432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110001011; // iC= -629 
vC = 14'b1111101001001100; // vC=-1460 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110110001; // iC= -591 
vC = 14'b1111101010001011; // vC=-1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010001; // iC= -559 
vC = 14'b1111101000001110; // vC=-1522 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110101111001; // iC= -647 
vC = 14'b1111101010011010; // vC=-1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010101; // iC= -619 
vC = 14'b1111101000100001; // vC=-1503 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110111100; // iC= -580 
vC = 14'b1111101000010101; // vC=-1515 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110010; // iC= -526 
vC = 14'b1111101000011000; // vC=-1512 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000001100; // iC= -500 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110110010000; // iC= -624 
vC = 14'b1111101001111001; // vC=-1415 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b1111100111111101; // vC=-1539 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101101; // iC= -531 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111000101; // iC= -571 
vC = 14'b1111101000010110; // vC=-1514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100111; // iC= -473 
vC = 14'b1111101001001010; // vC=-1462 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011000; // iC= -552 
vC = 14'b1111101010000000; // vC=-1408 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111110000; // iC= -528 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011010; // iC= -550 
vC = 14'b1111100111101110; // vC=-1554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000010001; // iC= -495 
vC = 14'b1111101001101111; // vC=-1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001001; // iC= -439 
vC = 14'b1111101000100100; // vC=-1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111010111; // iC= -553 
vC = 14'b1111100111110101; // vC=-1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011000; // iC= -488 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111100111; // iC= -537 
vC = 14'b1111100111101111; // vC=-1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111011001; // iC= -551 
vC = 14'b1111100111110101; // vC=-1547 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111110111101111; // iC= -529 
vC = 14'b1111101000100100; // vC=-1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001001111; // iC= -433 
vC = 14'b1111101001000111; // vC=-1465 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000011000; // iC= -488 
vC = 14'b1111101001000010; // vC=-1470 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000100; // iC= -380 
vC = 14'b1111101000010011; // vC=-1517 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001000111; // iC= -441 
vC = 14'b1111101001110000; // vC=-1424 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000110000; // iC= -464 
vC = 14'b1111101001011101; // vC=-1443 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001100101; // iC= -411 
vC = 14'b1111101001110100; // vC=-1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100111; // iC= -345 
vC = 14'b1111101000001010; // vC=-1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111000100100; // iC= -476 
vC = 14'b1111101000001101; // vC=-1523 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010001100; // iC= -372 
vC = 14'b1111101000001010; // vC=-1526 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111110; // iC= -322 
vC = 14'b1111100111110001; // vC=-1551 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111001111000; // iC= -392 
vC = 14'b1111101000100111; // vC=-1497 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010000100; // iC= -380 
vC = 14'b1111101001000110; // vC=-1466 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010111100; // iC= -324 
vC = 14'b1111100111011010; // vC=-1574 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011110111; // iC= -265 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001111; // iC= -305 
vC = 14'b1111101000111000; // vC=-1480 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010010111; // iC= -361 
vC = 14'b1111100111101100; // vC=-1556 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011111010; // iC= -262 
vC = 14'b1111101001000101; // vC=-1467 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111010100111; // iC= -345 
vC = 14'b1111101000100100; // vC=-1500 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100100001; // iC= -223 
vC = 14'b1111100111001011; // vC=-1589 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111011001110; // iC= -306 
vC = 14'b1111101001010111; // vC=-1449 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101101010; // iC= -150 
vC = 14'b1111101001010101; // vC=-1451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101111101; // iC= -131 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100000111; // iC= -249 
vC = 14'b1111100111010011; // vC=-1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101010010; // iC= -174 
vC = 14'b1111101000101110; // vC=-1490 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100111001; // iC= -199 
vC = 14'b1111101001011000; // vC=-1448 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111100101111; // iC= -209 
vC = 14'b1111100111000110; // vC=-1594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001111; // iC= -113 
vC = 14'b1111100111010011; // vC=-1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101110000; // iC= -144 
vC = 14'b1111101001100010; // vC=-1438 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111101100111; // iC= -153 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110001010; // iC= -118 
vC = 14'b1111100111111010; // vC=-1542 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110011111; // iC=  -97 
vC = 14'b1111101000111011; // vC=-1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001110; // iC=  -50 
vC = 14'b1111101000110001; // vC=-1487 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111000101; // iC=  -59 
vC = 14'b1111101000010001; // vC=-1519 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101000; // iC=   40 
vC = 14'b1111101000101001; // vC=-1495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111001100; // iC=  -52 
vC = 14'b1111101001100011; // vC=-1437 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111110111101; // iC=  -67 
vC = 14'b1111100111010011; // vC=-1581 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000110110; // iC=   54 
vC = 14'b1111100111011001; // vC=-1575 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000011001; // iC=   25 
vC = 14'b1111101000001000; // vC=-1528 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b1111111111111011; // iC=   -5 
vC = 14'b1111101001011111; // vC=-1441 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000001111; // iC=   15 
vC = 14'b1111101001010110; // vC=-1450 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000111010; // iC=   58 
vC = 14'b1111101001000000; // vC=-1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000000101010; // iC=   42 
vC = 14'b1111100111011110; // vC=-1570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000010001111; // iC=  143 
vC = 14'b1111101000000011; // vC=-1533 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000001101100; // iC=  108 
vC = 14'b1111101000100110; // vC=-1498 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101011; // iC=  235 
vC = 14'b1111101000100011; // vC=-1501 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101110; // iC=  238 
vC = 14'b1111100111100111; // vC=-1561 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011110111; // iC=  247 
vC = 14'b1111101000111011; // vC=-1477 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000011101011; // iC=  235 
vC = 14'b1111100111110010; // vC=-1550 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100101001; // iC=  297 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000100011001; // iC=  281 
vC = 14'b1111100111001101; // vC=-1587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101000001; // iC=  321 
vC = 14'b1111100111111000; // vC=-1544 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101010110; // iC=  342 
vC = 14'b1111101001100000; // vC=-1440 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101110011; // iC=  371 
vC = 14'b1111101000110010; // vC=-1486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110110110; // iC=  438 
vC = 14'b1111101001010011; // vC=-1453 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111001111; // iC=  463 
vC = 14'b1111101000000110; // vC=-1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000101111101; // iC=  381 
vC = 14'b1111101001101111; // vC=-1425 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000111011011; // iC=  475 
vC = 14'b1111100111111100; // vC=-1540 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000000110101111; // iC=  431 
vC = 14'b1111101000110111; // vC=-1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000100111; // iC=  551 
vC = 14'b1111100111100101; // vC=-1563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000011111; // iC=  543 
vC = 14'b1111101001000100; // vC=-1468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100110; // iC=  614 
vC = 14'b1111101000111101; // vC=-1475 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001000001111; // iC=  527 
vC = 14'b1111100111101111; // vC=-1553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100100; // iC=  612 
vC = 14'b1111101010000001; // vC=-1407 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100001; // iC=  673 
vC = 14'b1111101000101010; // vC=-1494 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001101110; // iC=  622 
vC = 14'b1111100111100110; // vC=-1562 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001001100100; // iC=  612 
vC = 14'b1111101001000011; // vC=-1469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010100000; // iC=  672 
vC = 14'b1111101010001100; // vC=-1396 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001111; // iC=  719 
vC = 14'b1111101001110001; // vC=-1423 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001010010101; // iC=  661 
vC = 14'b1111101000001001; // vC=-1527 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001100010001; // iC=  785 
vC = 14'b1111101000111010; // vC=-1478 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011001001; // iC=  713 
vC = 14'b1111101000110111; // vC=-1481 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001011100000; // iC=  736 
vC = 14'b1111101010001011; // vC=-1397 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101000000; // iC=  832 
vC = 14'b1111101000000110; // vC=-1530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110010010; // iC=  914 
vC = 14'b1111101000100101; // vC=-1499 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001101011110; // iC=  862 
vC = 14'b1111101000101000; // vC=-1496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110000001; // iC=  897 
vC = 14'b1111101010100000; // vC=-1376 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110101110; // iC=  942 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111110110; // iC= 1014 
vC = 14'b1111101001110100; // vC=-1420 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111011001; // iC=  985 
vC = 14'b1111101001001000; // vC=-1464 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001110011101; // iC=  925 
vC = 14'b1111101001011010; // vC=-1446 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000001111001100; // iC=  972 
vC = 14'b1111101000100000; // vC=-1504 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000010110; // iC= 1046 
vC = 14'b1111101010110111; // vC=-1353 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010011; // iC= 1107 
vC = 14'b1111101001001111; // vC=-1457 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001010101; // iC= 1109 
vC = 14'b1111101000111111; // vC=-1473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100100; // iC= 1060 
vC = 14'b1111101001101011; // vC=-1429 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000100011; // iC= 1059 
vC = 14'b1111101010010001; // vC=-1391 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010000101110; // iC= 1070 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101001; // iC= 1193 
vC = 14'b1111101001000000; // vC=-1472 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010001000111; // iC= 1095 
vC = 14'b1111101001011011; // vC=-1445 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010001111; // iC= 1167 
vC = 14'b1111101011001011; // vC=-1333 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010010011; // iC= 1171 
vC = 14'b1111101010101101; // vC=-1363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010010101000; // iC= 1192 
vC = 14'b1111101010100110; // vC=-1370 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011100010; // iC= 1250 
vC = 14'b1111101010100011; // vC=-1373 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111001; // iC= 1337 
vC = 14'b1111101001010100; // vC=-1452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100001000; // iC= 1288 
vC = 14'b1111101011100001; // vC=-1311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010011001111; // iC= 1231 
vC = 14'b1111101010101010; // vC=-1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100011000; // iC= 1304 
vC = 14'b1111101010101010; // vC=-1366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101101; // iC= 1325 
vC = 14'b1111101011000101; // vC=-1339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101111000; // iC= 1400 
vC = 14'b1111101010111000; // vC=-1352 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100010110; // iC= 1302 
vC = 14'b1111101011001100; // vC=-1332 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100100110; // iC= 1318 
vC = 14'b1111101010011010; // vC=-1382 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101110; // iC= 1390 
vC = 14'b1111101011010000; // vC=-1328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101011000; // iC= 1368 
vC = 14'b1111101011111001; // vC=-1287 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110000; // iC= 1456 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010101; // iC= 1493 
vC = 14'b1111101100010001; // vC=-1263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110000; // iC= 1520 
vC = 14'b1111101010110100; // vC=-1356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100001; // iC= 1505 
vC = 14'b1111101010011111; // vC=-1377 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010011; // iC= 1427 
vC = 14'b1111101011100000; // vC=-1312 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111101; // iC= 1533 
vC = 14'b1111101100001001; // vC=-1271 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010110; // iC= 1494 
vC = 14'b1111101011000001; // vC=-1343 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001000; // iC= 1544 
vC = 14'b1111101011001110; // vC=-1330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000111111; // iC= 1599 
vC = 14'b1111101100011101; // vC=-1251 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001101; // iC= 1613 
vC = 14'b1111101101001100; // vC=-1204 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100111; // iC= 1511 
vC = 14'b1111101011101000; // vC=-1304 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100110; // iC= 1638 
vC = 14'b1111101100000101; // vC=-1275 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000001; // iC= 1665 
vC = 14'b1111101100110101; // vC=-1227 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001101; // iC= 1549 
vC = 14'b1111101011000101; // vC=-1339 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101110; // iC= 1646 
vC = 14'b1111101100101100; // vC=-1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110110; // iC= 1654 
vC = 14'b1111101100011010; // vC=-1254 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101110; // iC= 1710 
vC = 14'b1111101011101010; // vC=-1302 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001100100; // iC= 1636 
vC = 14'b1111101101001001; // vC=-1207 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000100; // iC= 1604 
vC = 14'b1111101100101111; // vC=-1233 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001001; // iC= 1673 
vC = 14'b1111101100011111; // vC=-1249 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000000; // iC= 1728 
vC = 14'b1111101110001010; // vC=-1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011110; // iC= 1694 
vC = 14'b1111101100001011; // vC=-1269 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110001; // iC= 1713 
vC = 14'b1111101011110110; // vC=-1290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101100; // iC= 1708 
vC = 14'b1111101101011011; // vC=-1189 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010110; // iC= 1750 
vC = 14'b1111101100111011; // vC=-1221 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110000; // iC= 1776 
vC = 14'b1111101110011000; // vC=-1128 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011101; // iC= 1693 
vC = 14'b1111101110001011; // vC=-1141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110100; // iC= 1716 
vC = 14'b1111101100101100; // vC=-1236 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b1111101100111100; // vC=-1220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b1111101110001000; // vC=-1144 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b1111101110100000; // vC=-1120 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011010; // iC= 1754 
vC = 14'b1111101101100111; // vC=-1177 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100011; // iC= 1827 
vC = 14'b1111101101101110; // vC=-1170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b1111101101011110; // vC=-1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001010; // iC= 1802 
vC = 14'b1111101110111110; // vC=-1090 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001101; // iC= 1741 
vC = 14'b1111101101101100; // vC=-1172 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110010; // iC= 1778 
vC = 14'b1111101111000111; // vC=-1081 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b1111101110000101; // vC=-1147 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b1111101101100001; // vC=-1183 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b1111101110011010; // vC=-1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001100; // iC= 1868 
vC = 14'b1111101111011001; // vC=-1063 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110000; // iC= 1776 
vC = 14'b1111101110011010; // vC=-1126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101011; // iC= 1899 
vC = 14'b1111110000001110; // vC=-1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b1111101111010010; // vC=-1070 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000000; // iC= 1792 
vC = 14'b1111101110100011; // vC=-1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001110; // iC= 1806 
vC = 14'b1111110000010000; // vC=-1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111101111000101; // vC=-1083 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100000001; // iC= 1793 
vC = 14'b1111101111001100; // vC=-1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001101; // iC= 1933 
vC = 14'b1111101111110010; // vC=-1038 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011100; // iC= 1884 
vC = 14'b1111101110100111; // vC=-1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111110000100100; // vC= -988 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b1111101111001100; // vC=-1076 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b1111110001010111; // vC= -937 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b1111101111100010; // vC=-1054 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101111; // iC= 1839 
vC = 14'b1111101111011110; // vC=-1058 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100100; // iC= 1892 
vC = 14'b1111101111111100; // vC=-1028 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011001; // iC= 1945 
vC = 14'b1111110000111100; // vC= -964 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001001; // iC= 1865 
vC = 14'b1111110000011011; // vC= -997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b1111110000011100; // vC= -996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011011; // iC= 1883 
vC = 14'b1111110000111001; // vC= -967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111110001011010; // vC= -934 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b1111110001010011; // vC= -941 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111110001101001; // vC= -919 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b1111110001000010; // vC= -958 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100101; // iC= 1893 
vC = 14'b1111110001110101; // vC= -907 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b1111110001111010; // vC= -902 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011010; // iC= 1882 
vC = 14'b1111110010001111; // vC= -881 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b1111110001000011; // vC= -957 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010010; // iC= 1938 
vC = 14'b1111110000111000; // vC= -968 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b1111110001001000; // vC= -952 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111100; // iC= 1916 
vC = 14'b1111110010010111; // vC= -873 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000110; // iC= 1862 
vC = 14'b1111110001111111; // vC= -897 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000110; // iC= 1990 
vC = 14'b1111110011000011; // vC= -829 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001111; // iC= 1999 
vC = 14'b1111110011001101; // vC= -819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111110; // iC= 1982 
vC = 14'b1111110010111011; // vC= -837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000100; // iC= 1924 
vC = 14'b1111110011010011; // vC= -813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011000; // iC= 1880 
vC = 14'b1111110010010000; // vC= -880 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111000; // iC= 1912 
vC = 14'b1111110001100111; // vC= -921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111110010101001; // vC= -855 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111110010100100; // vC= -860 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110001; // iC= 1905 
vC = 14'b1111110011011001; // vC= -807 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011001; // iC= 1881 
vC = 14'b1111110011110010; // vC= -782 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000000; // iC= 1920 
vC = 14'b1111110010111101; // vC= -835 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111110; // iC= 1918 
vC = 14'b1111110010101111; // vC= -849 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000100; // iC= 1924 
vC = 14'b1111110010111001; // vC= -839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111110010101010; // vC= -854 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111110010111110; // vC= -834 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111110100001010; // vC= -758 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111110010110001; // vC= -847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100100; // iC= 2020 
vC = 14'b1111110011001111; // vC= -817 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111011; // iC= 1979 
vC = 14'b1111110100000100; // vC= -764 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111110011101001; // vC= -791 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111110011111001; // vC= -775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001010; // iC= 1994 
vC = 14'b1111110100111000; // vC= -712 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110011; // iC= 1971 
vC = 14'b1111110100011100; // vC= -740 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111110101001111; // vC= -689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111110100001100; // vC= -756 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b1111110101100000; // vC= -672 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111110100001011; // vC= -757 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b1111110100011101; // vC= -739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100101; // iC= 2021 
vC = 14'b1111110101011000; // vC= -680 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011110; // iC= 2014 
vC = 14'b1111110100111011; // vC= -709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000000; // iC= 2048 
vC = 14'b1111110110101101; // vC= -595 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b1111110101111011; // vC= -645 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000001; // iC= 1985 
vC = 14'b1111110101100111; // vC= -665 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111110110101011; // vC= -597 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111110100111011; // vC= -709 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101101; // iC= 1965 
vC = 14'b1111110111001011; // vC= -565 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111010; // iC= 2042 
vC = 14'b1111110101101010; // vC= -662 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111110111000011; // vC= -573 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011110; // iC= 1950 
vC = 14'b1111110101100011; // vC= -669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111110101111110; // vC= -642 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b1111110111010111; // vC= -553 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011010; // iC= 1946 
vC = 14'b1111110110101010; // vC= -598 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111110111010110; // vC= -554 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000111; // iC= 1991 
vC = 14'b1111110101110001; // vC= -655 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b1111110111101101; // vC= -531 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111110110100010; // vC= -606 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111110110101100; // vC= -596 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101011; // iC= 1963 
vC = 14'b1111110111010000; // vC= -560 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111110; // iC= 2046 
vC = 14'b1111111000010000; // vC= -496 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111110111111000; // vC= -520 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111111000110101; // vC= -459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111111000111000; // vC= -456 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111000110011; // vC= -461 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011010; // iC= 2010 
vC = 14'b1111110111011111; // vC= -545 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100111; // iC= 1959 
vC = 14'b1111111001011110; // vC= -418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000010001; // iC= 2065 
vC = 14'b1111111000011010; // vC= -486 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011000; // iC= 2072 
vC = 14'b1111111000010111; // vC= -489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001110; // iC= 2062 
vC = 14'b1111111000110101; // vC= -459 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111001100110; // vC= -410 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b1111110111101110; // vC= -530 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000110; // iC= 2054 
vC = 14'b1111111000000010; // vC= -510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011000; // iC= 2072 
vC = 14'b1111111001011110; // vC= -418 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001000; // iC= 2056 
vC = 14'b1111111000011101; // vC= -483 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001010; // iC= 1930 
vC = 14'b1111111001100010; // vC= -414 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111111001001111; // vC= -433 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011101; // iC= 2077 
vC = 14'b1111111001101100; // vC= -404 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111001; // iC= 1977 
vC = 14'b1111111000011011; // vC= -485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111111001101010; // vC= -406 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100101; // iC= 1957 
vC = 14'b1111111001001100; // vC= -436 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111111001010000; // vC= -432 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101001; // iC= 2025 
vC = 14'b1111111010001111; // vC= -369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101000; // iC= 1960 
vC = 14'b1111111010010101; // vC= -363 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b1111111011001010; // vC= -310 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b1111111001011011; // vC= -421 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b1111111010111000; // vC= -328 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110110; // iC= 1974 
vC = 14'b1111111010101110; // vC= -338 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111010010010; // vC= -366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111010110110; // vC= -330 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b1111111010000101; // vC= -379 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111011; // iC= 2043 
vC = 14'b1111111010011100; // vC= -356 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001001; // iC= 2057 
vC = 14'b1111111100000001; // vC= -255 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101101; // iC= 2029 
vC = 14'b1111111011001001; // vC= -311 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111111011101111; // vC= -273 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101100; // iC= 2028 
vC = 14'b1111111011111011; // vC= -261 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b1111111011110111; // vC= -265 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b1111111011110110; // vC= -266 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001011; // iC= 1931 
vC = 14'b1111111011111111; // vC= -257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b1111111011111100; // vC= -260 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000001; // iC= 1921 
vC = 14'b1111111101000111; // vC= -185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011011; // iC= 1947 
vC = 14'b1111111100010010; // vC= -238 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101000; // iC= 2024 
vC = 14'b1111111101010000; // vC= -176 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100011; // iC= 1955 
vC = 14'b1111111101000000; // vC= -192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010011; // iC= 2003 
vC = 14'b1111111101100100; // vC= -156 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000011; // iC= 2051 
vC = 14'b1111111100101001; // vC= -215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011000; // iC= 1944 
vC = 14'b1111111100111000; // vC= -200 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b1111111101000100; // vC= -188 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000011000; // iC= 2072 
vC = 14'b1111111011011110; // vC= -290 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111101; // iC= 1917 
vC = 14'b1111111100001101; // vC= -243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110110; // iC= 2038 
vC = 14'b1111111100100001; // vC= -223 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100001; // iC= 1953 
vC = 14'b1111111110001001; // vC= -119 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b1111111110010110; // vC= -106 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000000; // iC= 2048 
vC = 14'b1111111100001101; // vC= -243 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001110; // iC= 1998 
vC = 14'b1111111101001100; // vC= -180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111111110010111; // vC= -105 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111111000; // iC= 2040 
vC = 14'b1111111101000101; // vC= -187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000101; // iC= 2053 
vC = 14'b1111111101010110; // vC= -170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000001001; // iC= 2057 
vC = 14'b1111111100100100; // vC= -220 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000011; // iC= 1923 
vC = 14'b1111111101011000; // vC= -168 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110001; // iC= 2033 
vC = 14'b1111111110000111; // vC= -121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111001000; // iC= 1992 
vC = 14'b1111111111001100; // vC=  -52 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111111101000101; // vC= -187 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b1111111110001101; // vC= -115 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110111; // iC= 1911 
vC = 14'b1111111111101011; // vC=  -21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111100011; // iC= 2019 
vC = 14'b1111111101101000; // vC= -152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101010; // iC= 2026 
vC = 14'b1111111101110011; // vC= -141 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b1111111110000110; // vC= -122 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b0000000000000101; // vC=    5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001111; // iC= 1935 
vC = 14'b1111111111010001; // vC=  -47 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000010; // iC= 1922 
vC = 14'b1111111111100011; // vC=  -29 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111100; // iC= 1980 
vC = 14'b0000000000010101; // vC=   21 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010000; // iC= 2000 
vC = 14'b0000000000001101; // vC=   13 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b0000000000010111; // vC=   23 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b0000000000010110; // vC=   22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111111111100100; // vC=  -28 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010001; // iC= 2001 
vC = 14'b1111111111011111; // vC=  -33 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111111; // iC= 1983 
vC = 14'b1111111111010000; // vC=  -48 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101110; // iC= 1902 
vC = 14'b0000000000101010; // vC=   42 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100110; // iC= 1958 
vC = 14'b0000000000010100; // vC=   20 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000100000000011; // iC= 2051 
vC = 14'b1111111111110111; // vC=   -9 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111111111000110; // vC=  -58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b0000000001001010; // vC=   74 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b1111111111110111; // vC=   -9 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101010; // iC= 1962 
vC = 14'b1111111111111100; // vC=   -4 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110000; // iC= 1968 
vC = 14'b1111111111111011; // vC=   -5 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b0000000001000100; // vC=   68 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111011; // iC= 1915 
vC = 14'b0000000001100011; // vC=   99 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111101111; // iC= 2031 
vC = 14'b0000000000010110; // vC=   22 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b0000000000011000; // vC=   24 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001000; // iC= 1928 
vC = 14'b0000000000000000; // vC=    0 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000101; // iC= 1989 
vC = 14'b0000000000111010; // vC=   58 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010111; // iC= 2007 
vC = 14'b0000000010100110; // vC=  166 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010000; // iC= 1936 
vC = 14'b0000000001011100; // vC=   92 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000000010000001; // vC=  129 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011111; // iC= 1951 
vC = 14'b0000000001000110; // vC=   70 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111110010; // iC= 2034 
vC = 14'b0000000010111010; // vC=  186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b0000000001010010; // vC=   82 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111011100; // iC= 2012 
vC = 14'b0000000010101010; // vC=  170 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110110; // iC= 1910 
vC = 14'b0000000001100100; // vC=  100 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101111111; // iC= 1919 
vC = 14'b0000000001111110; // vC=  126 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101111; // iC= 1967 
vC = 14'b0000000010001111; // vC=  143 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110111101; // iC= 1981 
vC = 14'b0000000001100110; // vC=  102 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100110; // iC= 1894 
vC = 14'b0000000011000000; // vC=  192 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010110; // iC= 1942 
vC = 14'b0000000001011010; // vC=   90 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111010110; // iC= 2006 
vC = 14'b0000000010111000; // vC=  184 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100011; // iC= 1891 
vC = 14'b0000000010011011; // vC=  155 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011110; // iC= 1886 
vC = 14'b0000000011101010; // vC=  234 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000101; // iC= 1925 
vC = 14'b0000000010110110; // vC=  182 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b0000000011011011; // vC=  219 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011111000000; // iC= 1984 
vC = 14'b0000000010000111; // vC=  135 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110001; // iC= 1969 
vC = 14'b0000000100000111; // vC=  263 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b0000000011010100; // vC=  212 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000000011000001; // vC=  193 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101110; // iC= 1966 
vC = 14'b0000000100110001; // vC=  305 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b0000000011110111; // vC=  247 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000100; // iC= 1860 
vC = 14'b0000000100100110; // vC=  294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b0000000100110010; // vC=  306 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110101001; // iC= 1961 
vC = 14'b0000000100011001; // vC=  281 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100010; // iC= 1954 
vC = 14'b0000000100111011; // vC=  315 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110000; // iC= 1840 
vC = 14'b0000000101001110; // vC=  334 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101011000; // iC= 1880 
vC = 14'b0000000100000001; // vC=  257 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100100; // iC= 1828 
vC = 14'b0000000101101000; // vC=  360 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100111; // iC= 1895 
vC = 14'b0000000100111010; // vC=  314 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111111; // iC= 1855 
vC = 14'b0000000100011000; // vC=  280 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010011; // iC= 1875 
vC = 14'b0000000100100110; // vC=  294 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110110100; // iC= 1972 
vC = 14'b0000000101101110; // vC=  366 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101000; // iC= 1896 
vC = 14'b0000000100111111; // vC=  319 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100100; // iC= 1956 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110100; // iC= 1844 
vC = 14'b0000000100101101; // vC=  301 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101101; // iC= 1837 
vC = 14'b0000000110000100; // vC=  388 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b0000000101011001; // vC=  345 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110011101; // iC= 1949 
vC = 14'b0000000110000101; // vC=  389 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111100; // iC= 1852 
vC = 14'b0000000101101010; // vC=  362 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011010; // iC= 1818 
vC = 14'b0000000110010001; // vC=  401 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100101; // iC= 1829 
vC = 14'b0000000101011111; // vC=  351 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110010001; // iC= 1937 
vC = 14'b0000000110110010; // vC=  434 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110100000; // iC= 1952 
vC = 14'b0000000110011101; // vC=  413 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110010; // iC= 1842 
vC = 14'b0000000111011001; // vC=  473 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010100; // iC= 1876 
vC = 14'b0000000111010100; // vC=  468 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100111110; // iC= 1854 
vC = 14'b0000000101101111; // vC=  367 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b0000000110001110; // vC=  398 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001111; // iC= 1807 
vC = 14'b0000000111000100; // vC=  452 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101110100; // iC= 1908 
vC = 14'b0000000111100101; // vC=  485 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001011; // iC= 1803 
vC = 14'b0000000110010010; // vC=  402 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101001011; // iC= 1867 
vC = 14'b0000000111111011; // vC=  507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110000111; // iC= 1927 
vC = 14'b0000000111111011; // vC=  507 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011110001001; // iC= 1929 
vC = 14'b0000000101110001; // vC=  369 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011101; // iC= 1821 
vC = 14'b0000000111101001; // vC=  489 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101101101; // iC= 1901 
vC = 14'b0000000110101100; // vC=  428 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000001; // iC= 1857 
vC = 14'b0000000111111110; // vC=  510 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100011; // iC= 1763 
vC = 14'b0000000110101010; // vC=  426 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011001; // iC= 1817 
vC = 14'b0000001000000010; // vC=  514 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b0000000111010101; // vC=  469 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100100111; // iC= 1831 
vC = 14'b0000000111010111; // vC=  471 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001000; // iC= 1800 
vC = 14'b0000001000110011; // vC=  563 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b0000001001000111; // vC=  583 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101111; // iC= 1775 
vC = 14'b0000000111111010; // vC=  506 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100101; // iC= 1765 
vC = 14'b0000000111000011; // vC=  451 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100010; // iC= 1890 
vC = 14'b0000001000000100; // vC=  516 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101100; // iC= 1836 
vC = 14'b0000001001001111; // vC=  591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101100001; // iC= 1889 
vC = 14'b0000001000011111; // vC=  543 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100110000; // iC= 1840 
vC = 14'b0000001001001111; // vC=  591 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100001101; // iC= 1805 
vC = 14'b0000001000010110; // vC=  534 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101010111; // iC= 1879 
vC = 14'b0000000111011100; // vC=  476 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000111; // iC= 1735 
vC = 14'b0000001001101010; // vC=  618 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b0000000111101111; // vC=  495 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011101000100; // iC= 1860 
vC = 14'b0000001001000001; // vC=  577 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010100; // iC= 1812 
vC = 14'b0000001000001001; // vC=  521 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011110; // iC= 1822 
vC = 14'b0000001001001001; // vC=  585 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000001001010010; // vC=  594 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100011100; // iC= 1820 
vC = 14'b0000001001000011; // vC=  579 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b0000001000111010; // vC=  570 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010111; // iC= 1751 
vC = 14'b0000001010101001; // vC=  681 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101011; // iC= 1707 
vC = 14'b0000001001011000; // vC=  600 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110110; // iC= 1718 
vC = 14'b0000001010001001; // vC=  649 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b0000001010101110; // vC=  686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011010; // iC= 1690 
vC = 14'b0000001010011010; // vC=  666 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100101011; // iC= 1835 
vC = 14'b0000001010110100; // vC=  692 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b0000001010101101; // vC=  685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011100001; // iC= 1761 
vC = 14'b0000001001100000; // vC=  608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000001001101000; // vC=  616 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011100010010; // iC= 1810 
vC = 14'b0000001001001011; // vC=  587 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011101; // iC= 1757 
vC = 14'b0000001011011010; // vC=  730 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101110; // iC= 1710 
vC = 14'b0000001010101110; // vC=  686 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100011; // iC= 1699 
vC = 14'b0000001001100000; // vC=  608 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011101010; // iC= 1770 
vC = 14'b0000001010011101; // vC=  669 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011111011; // iC= 1787 
vC = 14'b0000001011000110; // vC=  710 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011011100; // iC= 1756 
vC = 14'b0000001001101101; // vC=  621 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110011; // iC= 1651 
vC = 14'b0000001010100011; // vC=  675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000001010100011; // vC=  675 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b0000001010001110; // vC=  654 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000001010110000; // vC=  688 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110000; // iC= 1712 
vC = 14'b0000001011111110; // vC=  766 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011110011; // iC= 1779 
vC = 14'b0000001011100011; // vC=  739 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010001100; // iC= 1676 
vC = 14'b0000001011010111; // vC=  727 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011010000; // iC= 1744 
vC = 14'b0000001011000010; // vC=  706 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010111001; // iC= 1721 
vC = 14'b0000001010110001; // vC=  689 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111110; // iC= 1662 
vC = 14'b0000001010101101; // vC=  685 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100010; // iC= 1698 
vC = 14'b0000001011101001; // vC=  745 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111101; // iC= 1661 
vC = 14'b0000001101000111; // vC=  839 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101100; // iC= 1644 
vC = 14'b0000001011000111; // vC=  711 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011001111; // iC= 1743 
vC = 14'b0000001100100011; // vC=  803 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001000111; // iC= 1607 
vC = 14'b0000001011100001; // vC=  737 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000011; // iC= 1667 
vC = 14'b0000001101010011; // vC=  851 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010110111; // iC= 1719 
vC = 14'b0000001100101101; // vC=  813 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011011000001; // iC= 1729 
vC = 14'b0000001101011110; // vC=  862 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111100; // iC= 1660 
vC = 14'b0000001101011001; // vC=  857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110111; // iC= 1655 
vC = 14'b0000001100000111; // vC=  775 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010101010; // iC= 1706 
vC = 14'b0000001100110011; // vC=  819 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010100100; // iC= 1700 
vC = 14'b0000001011011111; // vC=  735 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001100; // iC= 1612 
vC = 14'b0000001101101000; // vC=  872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111111; // iC= 1663 
vC = 14'b0000001101101101; // vC=  877 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000001; // iC= 1665 
vC = 14'b0000001100110000; // vC=  816 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000110010; // iC= 1586 
vC = 14'b0000001100100010; // vC=  802 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010000010; // iC= 1666 
vC = 14'b0000001101000101; // vC=  837 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011100; // iC= 1628 
vC = 14'b0000001101001111; // vC=  847 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001010; // iC= 1610 
vC = 14'b0000001100011000; // vC=  792 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001110; // iC= 1614 
vC = 14'b0000001101011010; // vC=  858 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001111110; // iC= 1662 
vC = 14'b0000001101011101; // vC=  861 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110010; // iC= 1650 
vC = 14'b0000001100100100; // vC=  804 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010111; // iC= 1623 
vC = 14'b0000001101011001; // vC=  857 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100110; // iC= 1574 
vC = 14'b0000001101001110; // vC=  846 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011010011101; // iC= 1693 
vC = 14'b0000001101101000; // vC=  872 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001000; // iC= 1544 
vC = 14'b0000001110100010; // vC=  930 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111101; // iC= 1533 
vC = 14'b0000001101110110; // vC=  886 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001101101; // iC= 1645 
vC = 14'b0000001101001011; // vC=  843 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110010; // iC= 1650 
vC = 14'b0000001101100110; // vC=  870 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001001000; // iC= 1608 
vC = 14'b0000001110011001; // vC=  921 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111100111; // iC= 1511 
vC = 14'b0000001111010101; // vC=  981 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010111; // iC= 1623 
vC = 14'b0000001111100100; // vC=  996 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001010001; // iC= 1617 
vC = 14'b0000001111000001; // vC=  961 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001110011; // iC= 1651 
vC = 14'b0000001111010001; // vC=  977 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011111; // iC= 1503 
vC = 14'b0000001110111100; // vC=  956 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011001011011; // iC= 1627 
vC = 14'b0000001111110000; // vC= 1008 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000100000; // iC= 1568 
vC = 14'b0000001111011001; // vC=  985 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111011000; // iC= 1496 
vC = 14'b0000001111010100; // vC=  980 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111110000; // iC= 1520 
vC = 14'b0000001111110101; // vC= 1013 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000101; // iC= 1541 
vC = 14'b0000001110011010; // vC=  922 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001110; // iC= 1486 
vC = 14'b0000001110001100; // vC=  908 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101001; // iC= 1513 
vC = 14'b0000001110001111; // vC=  911 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010001; // iC= 1553 
vC = 14'b0000001111011111; // vC=  991 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111010110; // iC= 1494 
vC = 14'b0000010000011000; // vC= 1048 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011100; // iC= 1564 
vC = 14'b0000010000101011; // vC= 1067 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101110; // iC= 1518 
vC = 14'b0000001110101111; // vC=  943 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000011101; // iC= 1565 
vC = 14'b0000001111001011; // vC=  971 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110110; // iC= 1462 
vC = 14'b0000001111111101; // vC= 1021 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001110; // iC= 1486 
vC = 14'b0000001111110111; // vC= 1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000000101; // iC= 1541 
vC = 14'b0000001111000111; // vC=  967 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010101; // iC= 1557 
vC = 14'b0000010000100101; // vC= 1061 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000101001; // iC= 1577 
vC = 14'b0000001111001100; // vC=  972 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001100; // iC= 1420 
vC = 14'b0000010000010001; // vC= 1041 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111111011; // iC= 1531 
vC = 14'b0000010000111100; // vC= 1084 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101000; // iC= 1448 
vC = 14'b0000010000011011; // vC= 1051 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000001001; // iC= 1545 
vC = 14'b0000001111110010; // vC= 1010 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000011000010111; // iC= 1559 
vC = 14'b0000001111101010; // vC= 1002 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110110000; // iC= 1456 
vC = 14'b0000001111110110; // vC= 1014 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111000; // iC= 1464 
vC = 14'b0000010000001101; // vC= 1037 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001010; // iC= 1482 
vC = 14'b0000010001000110; // vC= 1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101000; // iC= 1512 
vC = 14'b0000010001000110; // vC= 1094 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110001100; // iC= 1420 
vC = 14'b0000001111110111; // vC= 1015 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100110; // iC= 1382 
vC = 14'b0000010001010000; // vC= 1104 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111001110; // iC= 1486 
vC = 14'b0000001111100101; // vC=  997 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010111101101; // iC= 1517 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010101; // iC= 1365 
vC = 14'b0000010000101001; // vC= 1065 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101101; // iC= 1389 
vC = 14'b0000001111111000; // vC= 1016 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100110; // iC= 1446 
vC = 14'b0000010000111110; // vC= 1086 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100010; // iC= 1442 
vC = 14'b0000010010011011; // vC= 1179 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010000; // iC= 1360 
vC = 14'b0000010000101101; // vC= 1069 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000101; // iC= 1349 
vC = 14'b0000010001010100; // vC= 1108 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101010110; // iC= 1366 
vC = 14'b0000010010100010; // vC= 1186 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100111101; // iC= 1341 
vC = 14'b0000010000111010; // vC= 1082 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100111; // iC= 1447 
vC = 14'b0000010010100110; // vC= 1190 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111000; // iC= 1464 
vC = 14'b0000010000011111; // vC= 1055 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101100010; // iC= 1378 
vC = 14'b0000010010001010; // vC= 1162 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101000010; // iC= 1346 
vC = 14'b0000010010011010; // vC= 1178 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110111101; // iC= 1469 
vC = 14'b0000010010100001; // vC= 1185 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011000; // iC= 1432 
vC = 14'b0000010010111110; // vC= 1214 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110101001; // iC= 1449 
vC = 14'b0000010001100100; // vC= 1124 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011100; // iC= 1436 
vC = 14'b0000010001110110; // vC= 1142 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110100001; // iC= 1441 
vC = 14'b0000010001011101; // vC= 1117 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101110101; // iC= 1397 
vC = 14'b0000010001110100; // vC= 1140 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000000; // iC= 1408 
vC = 14'b0000010010111111; // vC= 1215 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110011110; // iC= 1438 
vC = 14'b0000010001110000; // vC= 1136 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110000000; // iC= 1408 
vC = 14'b0000010001011001; // vC= 1113 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010110010010; // iC= 1426 
vC = 14'b0000010010110010; // vC= 1202 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101011; // iC= 1387 
vC = 14'b0000010001111110; // vC= 1150 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101111; // iC= 1391 
vC = 14'b0000010011110011; // vC= 1267 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001100; // iC= 1356 
vC = 14'b0000010010000000; // vC= 1152 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010100101111; // iC= 1327 
vC = 14'b0000010001100001; // vC= 1121 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101001100; // iC= 1356 
vC = 14'b0000010010011100; // vC= 1180 
#5;
clk_100M = 1'b0;
#5;
clk_100M = 1'b1;
iC = 14'b0000010101101100; // iC= 1388 
vC = 14'b0000010010111011; // vC= 1211 
#5;
clk_100M = 1'b0;
#5;




end





endmodule