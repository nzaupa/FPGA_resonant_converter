��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m���ҫ�_���fW�������e4���S�7$�%a/�J�}/���|�跞*rK��1�`ʑ�Fq�5���:�.�v�>���]����@��L>-��o�N|6��Ү;��F*F����!PC�u�#Q�b��Ap��lĳ��gY@0�L�$�$�E�?�EC0����D�#2�����[����?VB[�2 u ��eY,�&�$���"�!���L�c;��ֵ��f�L
�u��o�J�j�t
�ܻ��R�4��\�zA�李xsH�#d�q���CM7G�t������l�J{ j~�u^����N�a;�����Qv��_�����#<��u���8�Z'�@Q|1��h%PT���b���Z��$x��/>d��~�w�#Lc��v�ڀ��`r��T,�h�➆�Co�������i���=Ɏ25[1�9ο��$:�T�����:�V|˔Dg �:v/~X�1h%<^M�Ë㸏��?e$�F�8w�"�@���]E s	��ݑ��X�ڮ�����?���Y*�V��I�4��	�2c�މ}�
TX82$Oל�ga.�.�Y�~��#�Ɇ��³��iچgf�U�B�ej�R�2���(�r��&è�YW)�2bF.[�GԎ��F�7� �A�^���C�B*W�axV��h䜼*7���ܕ%�J��ǰc��<J_IHF�����6���R�W���r��b�:�}�ޥ���tm��8R�� ����d\���D>Oj�a���j`�����K��h��Y��f�����#��)i�uh<�`���$zչ�T���~�؊�/Gq` �`�O՜k��3�kz��}�
N	�Q&e�����9;��M���b���Ls�}qcR���ׅ�
���"�����R�����~&7�iǁ���_.�;b���m ʖ�+o�ҽ(*KzUz�جm�u���\Z�@x�ڽ@N�����C���N��	{���r��Uu�&dYۺQ�dD}���5懈��Z����yw@�p>OoW�z��n���P�0Z�gY.f�e�����<�V3�����6dWm"�4^�!�"=�ĳi���3k�z�ژLZ�k&���'Vɫ񈎲���B��殩�4�u������,��r�A��a�6�v�[��]�8�	qv�g�	���uY@��ӛC�I�����8��ÏJߡ����RF���4H��U#]��-��Jf��ӱR��`�'�KEq	�7oE\��H;445�뺊��P�Ԙ�Kl=�o�N���K�:�����X�!���f�,�FZ��_n��?��Dk��A-�L[��9髠��4�)rg--f-*��o|Wg������n�����4���W�c�,[]��K@�c�ƿ&j��=L[ù���Q�*fI7�*�/���p�s[Ic�b��<N)8'd��c-I���pq��ID@!_�n2�\���Mj�$`�d	0�(=��ڷz�� �]縩}������t=_�;����~���0�<!�����4�©>�f�sk��,�KN鈇a������Ұp1=�(F��Q�MD��O2 �,ǳ��*G��,��-���]�yT��b+��0��y�Ѓ�K�'��8L�VI����&���n��SԳI����M
G6i�}jj��ԅIr7��>�47?�8 �h��S�|K�͂�Z5��WiN~'�w�"A쵛E�r8�����2��ޡ�_� ���-��`6f��0ke�Xʯp�yq&��w�������;?I��}����-�Q3Q)�k��f�A�A��9 "M@0�<-ڗ���Y����ߡ:�b$M�C��a������'d��y �2����=5T�T�Z�eW[�&�}�`�L���b���!��R�6�X�7�0�]tդE{�vg"�=w��c��*����kzU����X�4@,���L+[~�+��´��%���4n��J�����E����r��G��r�
�\Oc�&�����)?T�P�O=��Ղ�v+��8[8H'�W���whs�ig� �gB
�w�dҘ�{�t�W�V"�4�O��ǰ���ldʤd<+���ɓ`3 #���d�t��:�>Xփ����ܜ	�2��o
y�%��{�/m�������3qkޒ=�+��������Nw�4[������.<�B[l8y�>=����+��7�;�����1K�>�ĀY7�04P�*V%�<o�q���Ų�E����(�םo��|�xF�Q>�������;gN�����
CZ�&��z�"�����1�q�0R���Y��%������?�d��=%V��t����';�+�A��ά�� :����;~���%�- F&�s'���	�c]��w���❩����x)��a�G�t���$�x��)p����e���.�T��	��	�4BXY��U��6��H5�pԶG�u۩��(�܀)�������#�mǩ]���2*�G!𙄣l`�X���lLD)P�<�����VS�Ʈt3Tף�Aj���]���G5'�o�UEd*����뛓��2��,� )��,#dGj�Y��s��'-���=	��*Z�R'�k��.`y�D�'wr!�
)J.Қ[�N:?Ǿ� ��M�3�����Â!P]Jr4��/����D��QaH��7��>�y��R�P�lѸM�f c�s��+�-Ŗ�>����������r�'�X������T��n-3[S�/�*a��%��7�� 8�R����`l=�5��yZ0ժ�z��9̵�.e���u`�#�z����t������|�9��F��V:��~2����NJӋ	9��}0�Fb��ԧ-�I(J����?��J���a;Z�xH����|�Ӄ3�*N�w�ޒ%�P���y�{,�h�3�!]֋�|^.W��GQBꮱ^���Z�)h�n;	ߑ��h�?T�᤼E��\��x�޴(Sɘ�v�����ƣc�cL�/�_�R�.��2l.�뭑�yU<I�?# 
6T�x6��8;J����;�ƙB?"�xd�v�����;EZ2����h�iش�D�l0�6!AwK��܂�>t_L�a�quf=lf�4�R�W0�`�Nl��k9�	Z��p��N��x�O�R�1��k�B�?4��̻�^�$�ʉ�,�� �:\D��Dm1�΄�/oJ�L�Q��O�lC7
�5��1͇wYu�[��	�3ŐҌ� hMM(���|,[ �A���C�9�
�gD���7s(ǃA6o��� �Γ�y@�%�d�,	���jv�A����gsk9m��/�5�Z�]�H?�'�����]�?����r5BA�� ��;{��&8��l�!��rI��=T�7��B�y���(c��d��R)+*��j[_��9)	V�(���^R M��nҀ=����y��s٥d�D�=52�۵�s
s܉�T{컼�0��	�S'���(��\���4{�č����.*�Q���5�RJG<T@��b�j�r�Y��c�]��~�����yti&�|�_J�p��+D���O�����㸽ߣ��bs��|!���m  0�J�O�	�A�c��ؕ����/	,P�8S�⮂�c����I���A����3ey��V`�u��_|���WZH�*▏#������,]��$�F<I&&_�E��I=����W��ˑ^�WK ~w�I�p��Øne�1�5�=�6�&b���Q� Q�|r�;���>6�-�a���4�!�r3�����:� �ع�S��9�a���i��y�=����X�D�)�?�!⫊(1�)�Ј�Y�;���>��
&M�qh��p�cc���TQ�F��r�*�fV�?���V��J��Ale�� BEX_�;1�D�@��Fd^[��S#� ���Dy�r����L���cH��\�kB��`�UͿT2��3#��1�b���=R,�h%}��z���~/\�|-^[6+I��Tt������#%&��|ʿ�o�-��<]`Yv��~�O~{���(7[A��oQo�q�w����4���,�t<�=�I0�'��1���:�pVh���. wG�g�?t��ٛ�M�k8��6��E6���Ӡ��R����b�\��g��j4 hE����D�
���j�����c˦8�C��e�O�eg��U��[ +�!ǧ3�������D�RقB/Ӂ��ᨆ���[@�@��Sb�9n7�x�����"]
g��J��2�9Ơ�����2��]��gc#�
s -�D/�U�!NA�`Ixzs.A��qz��ݍ؝K�45!R<?�<�n���w�ڳ��os�#�"�v2rCˆ*�ui_�X:����K��e,|�� ��J^���l��r[<v��}& �7&̘�ݰX���gp���%�V��Vk��H���l��T��<�&�?B+�Al��^��E�:�����п66����8�1�s>�o��})r�)
�!�x~�x�*��a����}]��=�>ɛ�|&��h�uW'����"�<�Jg�I��-�!��f�r�~.R� lY�^Dұ u��V����O����i���%��A�& av�b��@E�;%'mU�4g��of�рk�ϭ�V�I�� ?Z�`�q`�'W h��~�����
e�*Nz��u�ǭ O�����-U�j��0�\���p�,k����~������!۶T�����6K�^5���2J�N�uf�U�s��l�F�#!mZ�`�R:���$��[�q���_�g{�q(�������,�`��x��0]76��{ݜ� ��L�;=�w'*}tQ�v� r��jg)�*��B��֣.ͫ�Ν)�!�R��������l�4ܚ}]��/8��l칄ܼ�f+yG�'�m�8g�]>rL���'͉^�1��5�q�B�x�-s�h�{-\	��=��{������UB��k���	u��e��]7n������U6���Exh9x a�R�~�n�}��}:I8a�N��J3 L�&�o=��T�ii���-�sL$EG�,�y+6����t��C���"@D}ciAv�P�c�sC1LT�dV��}�����ͷ)�O9]vU +h~�ջ�N�B?q��h�o!�վ�m�~ձo�ƂZN�Y) �1��D���ᇊлOS�D�:'�OTI���7��[T^��Я����~?=ݫ"�����ATV�Yl4�<��{���֯kMQt,�J4�-ά�֌6��NP1��Y�#>Y��)�������D��_�'͇�?�〠�/>��z��j��1$�I٩TA>۾���;�l�B9�JSW���+$0�U"<CT��!�]��Vyh2Ĕ�t�Z lǙ�>�|)�\J�y�,/su�l�):�=.3Q�ӌ�� A�7e�'�#Qǈ�,2�H�@������'���9R�NU��s <��`X�{�!�=�	J�5� ���mSժ��U<z����/z��fϏoL��|v��fOvsnc����tҰk��<ƣ7���!Xv?�&�5F��;B��O�U�HX�h����
+�J���G��`�%h6p��̱5[/��P������S�,���~�L���M=�O�X�
BMi�f�
�~>t�^�c/�P��NShH���J%{�%���@	���@�Q� 5�O|>��7�1��#�X�rl5����juɃ0�:��H\dZ8���q��c"��F�rP�݅����L_{ܬ����FU�]��Ke�	���]v��t��̫���f�+yAG��,����uW*Xн'.�,P�H6J@���7;�!�i 1���VY)hw|5(���b	��oo�,���x0�kJ�i���0�^0�Z���z	���/t�ÚK�É`�3�wZ�Î��H�[ ��%�e� ���j؝�rn���s��^���A��~H��2��ӊҩ)�dm�FIq&�`*�����L�����G���JTC/^��nJ�h?F���RW��V�a�����S�� ��}���nu�p�;�&���IˠTst� ��$���oN��/oavS��'UGd����#��@b�Ex�5l�ʭ���dh_�\�\$9�Q�;| �8 ��ai�y00>/���*��7v�-g�'���z6E�t�N#�Z��D�%�fT�S� �ۆ��0ځ�z���pAp��Acx/�@"�B��4��@S6ٵF�&纬+H�|ὄH.6�Lɹ-f�[�ML���s�t��0�J9�B�s����T��Sd�Y!���N��wr�X���q�(�ij_�R��A��wUr���K;2T���J;��+Qb�%�B9��3��y���<Etp��ʁ����xdh)R��qT���61�4�
���]ă�>D�޹�9�z����r���N�}T/1Zb�6a��I��B?�4�mV*�0�aP�>��I�GN� io|o����	ft$��Gvn!�h���b�i;i��z�O�=�^"=;_�n�V���nt�����bv�,��t3Q��l��^�rP>(�X3Y�?��J)�	J/3�k��L�ǫ���8�J���`Zݼb&����ݲ�Ϋy�^�X[X.��#|�	CV�nf�y� ȗO�T����m���'"�pY\uZUћ��$e��a0@����R(�z[�؉���ϡU&$t��h�e��N�N�@R�/�����o�hvՕO�fi�*ϸp�f>�����������)c���$[ۣqJ��܇to�B�0o����.Eį���7}���O��������P���5n�Vz!Иʁ������z� HbV=�,��P9�p^))��R2�.�8<­�T�:�LC��\p�Ӫ��
���`Y `�px�L�_�6�� q���՗�Њ�q
&�%7�j�[��G	{d�Q@X
���ԪHj��7y�9�﫸�s�Bh�}T�X��w�U�8�M�7W��������W`<`6�̀C˝]<���s����y���k�J�E���/�j@\��u�m0�~B��C÷3E�W pV�:��Lu���C"�����0iV� �6cCuz�k ����א�I�-�YI�����!ۗ���LxjxL s�{z��h�5�p�C �O!%@*�������S����B����&��\2TK^K�ae�K5V:�ș�,���ǿaAh
�
˷Yn�ol�ǛL�YN��&$!�R����O;^�CX�ZysO�I�5!�*�4�]��}k{i�w	�����MtJQ��/���Qf*o�{oV���ڢ}s�˟=�]s$�iA�x��ֻ�Ok�ē8\Xcb�hЖM*�Ή�w~Y�~�s�Y	���O�a#�����,��G�8�g��#�Ř�=��fW%M��y�=�ˁں�,<	@00x"N�ʨ�Gb?�8�7;���_��k���Y��tva�u������;u�~\IH2zxP��B��L��⼵>�����"A*��m'׫�@��fOt�1ܻ�v��U'�(��^!�����h�Y�N#A��TʲX���?��f��uv�M��{^�Q��eA�����q�,6W�r�'�[�)dY��s��?l�5׹���ҷi�<��:���u">XJ��g.~�J�Asί j��4-��ohd���r��^E�t��\�1˒�r:Kq���$����^9>��|��9ҟ@�ףC�����9�ef�u��[&��v|�^������Z���y�׮w�jl��J5��'�Ebw���X�����#7��2T �l�#aA�t<��B��$y"�#@l1u܍�JU�[x�^N���[}jݖ����M���%/��GvGnK0Lo�V~a�K��k��l�6����_}��L��`Vy�%�t��BdX����7ӌ�9
 Z�T] ���
#�SG+��4��UH��U�s�p��ﷶ�/�uֵ�&�G-��^�n�-��V�{Lop����R������n1�u+lD��9�^�]�pV.��w�oV��c���I�������Jא�T�W%��ǳ�ff�Q�wU~�G 3�IBzڬ�9s�r�H�m�$�hfBW�w�eh|���Sِ�N�zY$ٍU1aA��$�֥ ,���x�OeOF�v�0.���!�賺�ڕ� u @V�2d9J��L*S�$��k{uM��9d�v�4v:�����7[U~qq��*{��e �ùE��P㖷`�E����3ʡ��5��v�d���;��=���}�m8Bg]�
׿�b����Ob<��\�=�9M:$�2 �Ka��\���r	�A���3cأ9��j'6>�0&�̐���t܈�)v@��%����)6�5��wk/���Vs;b�4Ƶ��Be�KV�ko0dq��>��N�@Θ�;|!d6̟������`\�|1)ئ� �Bi��g[�0�p-+	r�)2ZF�H����������=	r&�wg(��G�RF�s����Rl�߁ˤ TNô6��(��o��.�k'���=�>M��ٌi��,(d��Ydq����e����E\�t��ѽ����Ok;���dX��Hv�p�,�_��p�l^���5�4�Vȁ�ʆD��A�y�WbA�wd����\	��(��4���c<cʚa\�PIp��m��L� �AC���m:�v��W伂Me񭷱{�J@��8��m	��N��H�o���S�8��S�>t���t��#��	�ě��m��!c_�Zȣ�\ö�$ލlӑ�7�+�R�U
��tw5Ɗ#A���V/,���S{�뛰�g@��k}��=�}b����YK�0F�^���&߅U��Ձhn�g9I_���
Ϣ���*�<$Uc�8ڭwZ�"����5���;���P��o&)�.��1i��K�/���/�֕J�o)�6�����3]'�ԑ��`W�p��=���7����1SA)KZ�F��D�klZ'�S}^o��k\��w�6-�42�2�f�V�*ؙ������p�5������]q0s(D�ǳE똺�<�j>�O��5�`4�9�$1��cY�Ò�j�)���@`�U�m.���������ZH�o��eݒ���;���bV�8 7������)b��K�>Z	[;�p)1)s|-N�, g��r[�ܶeR�ah~�F{�Y��o_���[a���|��Gq�N��7���,�K�y�V������(��Ck��x�Ѵ4��;܃^8�*��-�q�x�WD�6��X��6�/>��)��xENVΙ���ݩ���]t��M����_�(U����VO�w�cry$���T'�᱓=�C-�J�a���/��~���R�Oӗ<?u��y>X�����?8�C���N��=W������c|�^
�+�����9�[5[��N�vP��>��Ѣ	���M��&��}4�D��� �meZ����O�.��Gc��'`�O'����,,S�b;�a���ȸJ,S�#>����O�R<4�Ŏȃ�"0�����I�E,�%��ݩJz�+�1T8t�F�fe�7-Q_oU#���uB�����Sz��λ��6f�A�C*`_
e�cO�Sj"�u7g5F|�	ػ�~1�S�������5��G�����.�@�Gy?�wH�I��p����^�M
����L����iƗ4)���d�bmZ}��f��u�Hy�bHK����b������Z-V����6��I������7�}�d�	�]��)ǐʅ��&*�r���4#�&��1��RS~B�ԉ���@�ޣ�ps]پ�|q�� �ث�HHweuM�4�zM�q���@	%�����;���������	��Yjψ����2!k`���}`��f��*�_Ϣ�}������%��6!a�_�i�T9=�PY��#�Yw����eޜ]�]ĐAP<�hB��؆4�m~��p���3?����<1h����ɹ �M䣶7 l����i�L��L�&�\U���ף��3�{}�݇�'���3�HC�P���,5F�I'pL*�G.Q�w����sF�7���>��lɭ4.��>���&��(B����%WS|��B�i+*�$�>���A����CoM%,���S]��p&�E��ȤO�ɘ֘�]+���B��Q7�n���a9�;�?��[e���([��_KcM���S{��� =n�3��:}�8���{pk"U�MP����7���L���`W��(
4Y��Ar�o��n�ew�t44j�����D�r0sEl�z�@�� H+I�����hH^�������j�鮖�%��p�!�Ak����I�&�eu������-�S�R�?���lm}�f��3P"���Q�8$�[v�
��L88�]�|��7��m���afc@���b�l'>��ſ�}v��#z,����
aP�`��n�PѨ��%-sK6Xu������MD&�E��8�2��p�&��ܞIbx�f�����"�F�7�U��'����rȰ�O�~q� )Iw�Y����mr�E�����[:SH���6U��ϸ l+ls7�6��Ks�gj�E=w����[��ɜ�9�[�Lca�\%���4�ü���EeL<�#i?"2|B��-Y[��P�L����A�ҶL���S�3'u5T����ݎ���xT�Kͱ�m;&b��z_:7ۙFoFӳHq�
�Ze���v�|J�IZw�ĿJLҕ`�Γ�G�ȽIj���w􊰋jS�$�6r�'���γ�(�xr���<��K�,�����!�	ȍܭ*�?k�/jjɫ��x�q5�U5��!�gVV�z��ڟ5nQ��ۣ�:@"^����3�s`]+D�Ɋc;�x�Z��<��N���޻��3��}Uj."C�ᕀ��ϔG�5�MnR(ߝα�u��H�Ҵ�c��ɶ"/�+���H��;W1�,�������=-$Q�q�4_�Oh��I��h��������.�������7�[b�"�e.��U+�~��wy�%����������h�-!Zy:�������`��̚��+BJ@F޾�Q�N��A,\���o�deֈ������ņi���#8���.�J�&���y��ޞ;�0����J�q`Z� ߞW��ᅉ�<��i��G�ʤ�.�����jf�K���H���dj��)�0����&Gý)�?���-��/_R�F���� Q�F��_�rү��CK����E�kc�����έ��j�w�HFCw�
e�钷^�5uYɞ(�#?�-঍R��c	��ج*c��`�����yٕ�p�o�ȣ�aL�����Y���7sj�������^?�;A�MӥaFY���	}naYnv������8hg�>R�����~	���
�8T��0;le��܉��s���Ց�� F�LZc[چS�B��I�Hp��u�l����E�E�U��l�%.�w��bw�����Da�����.��S�ͳ������ �bE�K.��)ɢ <�=�'Aɀ�1��ߟ�����
��..0v�ӣ��A��ڊ׼Ʋ����8 \b�=��k�����H��u>O��H��C����;�rm�P�XR�.|�(7ym.>�|	�v�嚝#��n��m�\K&�����E7�3���|�MS:оW��:l���#y�5ߜ����N-�	!��	>D��R��7��~*�.9���#�$�/&�r�H������Z���E5:v�h.�ν��;^�d�N�2e�(d�2e�L�d��T�,\������!8!-���Z�7c���#ն��o<r���M�d�}����7u?���'W��6��F#q|"��{/��y�G��|�"�&O��\��"״�y�c��$_Uμw{:PEm�c���k�����	�쾫l˴�:�u;��tx�Gv������QӀ(�o�-����k�j,�0ꢃ�F�JdtJ,oG������}���x�2��8b�'Y���I~C��.��yф�L��sa2ˍ��:���?ͽg��9>�Pm�ۜ!/��R�fX��
�yx5��Q1���̾����!��!9�b�ݲ���	ʥ�&�A���W�$� ���n6���#Z�?�\2k���87"^�b��Þ�F��+��n����F���X��l��\Pn�e}���/5��p*I��L��p?����~� ���ei��ww�,!h�(�%>�����u���Ǯ�L���ʪ|f�
ڣR(��NX���R���!2bW���%1'N�	��<V8t�t�C��@o�4a&�����*ᔃ)�������mK���AW���8)���t�����`���/f;�p���$�gʩ V B�&T˰��K�o�[���D3���l	ޥ��[k��y~< o�nh��>�F��U��ۮGR;������ן����ͭȴ�OaB4������OC��#�F��ZH,K�	i��I� ~q"��r��кk�:��+���R�qo\_kǪ�L`{/��S
y���PCd�%��h��n�d�Jm�����#�]k*��FdB����с0F��h�C=i���P�a�S���R�H� �ƛP
�[䍛_�½�Y�k�x��(V�b6�A�jO'p-���ޢ���������<8�����@�C�Z���;�Ey����R?"N�!��L>�����M_���^����b���ʕ���u�r#N�š�9d�U�A�ݣ����!�uU���٭{�U3f��p��s�:��S�o��F�x�{8c��#�������oq<m���-����04��F $W(���W�}������L��)a���ڍ��Ls\F�RX�#�=K{���;ݓY9C"ڿ���}�Z�M\�ax�J_��4VG`B�inD!��cz�U0��Bd�����4SN'��;�`QO�}?a��s�5S(��-��4�-s�J7�ŗ�d	���vS���e��I�/+���d[�0�z���L]�r�=&��e膆;���K��a5�ln�@Y�5fC	C�nP��;FWw�V$]���U����~RS{!P�ɹ��]A�Nj�|0ę�A�5S,Ȗ�`Lxo�A��t�__%3&�o�x�=����^�����YQ�fN��(�r@{m�JϟO��Tȥ���g7�����I�l-��Zs�=g�GA��������t�@�o=�fZ���*�t]�yY�v��c�� >�(˟o$�p��#t�[�5'`	A�cEg��1��@��8g�ų�^8���:{�%qtR�M���F� #�kQ�6;����tGO�X�E�e�j�0�3�'+���c��	{᳇}�栄��B@)�	��72���<���yB��X��'��v�TJ�Qviӈ�89���~�4ؗ��V����?v�&LC���[ ��_�a�X�^[��%���ԼQ��4��_S�L���6�>\l"O��S��KL{X8���Պq�YT�^òm��kzԟ̩�!x�C�NBv>qu�y���������F�d�G�陵��Ʈʜ���D'�[3�=��$�l��g]
&=�D Uf���A�Q�r�Ƣ�'�(�&�b����kBhk�/;��:��8�f�4:�@3��SU���)0z��%�К}!/{��9��@tw@��V����P�S����䱧�B��@[%�e*��@�[�sJ�2�)g[���)�Y�������gD�;�(�z3�7*"Q>Av탒���N�+P��bǷe�9�ԶW֜�|���0Ǡ��D)E�@I�m&jV���γbZ���kpq�E5�og���ˉA�o	�_J8@rHݣ��c��8�CA����#SA�W������)��e�ѣ���~I�C��-'�EbaN��w_\���%6���^� �٥|P��EX�WLR�dӚ�d��bT�%�Z��%�=��GX?C��M��y}�#��dCE����U�뀔K�Mz��t��ұ6fϐ�&�NE��/� �Y� 7P���Q�#2ʚ�s��:]䅈��;9ݦ���fI��x�ye7z���	N�e��[�(6���̃S�XS��*t�?����c��=s���o�f�v�'*��l���·	vU{�~qЪHMX��>�i�<(��_o��=I��C��z�u!����q=���v�J�?��{���Gx��7��b�=$j�C��we���̍��#���G^Z�=dY;E��b��6�mr%��:��É�ZvJ�.�+���<�>��u�Pa��9�+ۿd#��R֞�(�W�O�E�]�Y�Rx.��d~�U���ܦh�<�1���V�:� w={y�S�hu�) t���BK�S��.B�� s��ڃ1�FO^�mO������噐ss"ĹF�U�=s*"G�[s��%�+G����C�C#�>2�`H�~ez��!A2��D����|n�v@������`����Iy�@��xf3?.-tұ10�w�"�
�2~OF)�F� sI+���L3gm������9��(ׁ��ܐ�s� %�=���Y>��p��Ȟ����}>k���%���Zp�&��� �����<d�Q��{�[k��m^�E�\�T�G=��gc�hP�cm)���f��`"�G"&ӟϞ㿡yq8����"�|�Bo'�Et,���܉�-��=ְ�����Ԉ%M�yp��{`5yaP;�p@�)"�j��E�iZ�
������F�ɳv[�Y\e�RJc|�����u?���9*�;!%Y:�W���@�����u�\L�ֿ�+�����0��D��Q��~�tG問]b����8�Wr��Es�Y3:��`+�4 �?�K�O�պ��V�\���^��~"Qv�<�Њ�M$��n�������(�tfc�$�B�@$Y7��^=��+v�f����?�v�d�F��}��V l;um�)����rGg�_Z����߲Ems���B�φK0fm=ˬ�K�eK�0i34��(�-��R
`(䜼 Z���N�����F�T1Bk�����*��2���eⳅ��*B+DI���s�����c?v�F�U:�.��3t�f�Ţu�M	�Pg�m*�:k(Sk)��W��ʷ�\�W�0���A�u,�����"�-�L>�b�Qͣw�i~6�]�i,��@q��n+�в��j�ѫ<���I�xN����V����cjql�r�l�f>�L�c�3I]���#�
�"��D6p�K�2y�Ǔ8�X��/��UMX���E��]IT	�h��y�<���U9ңJ_�߃�`v��n� �}w3��0��2�,bh�č�9L"8/�)U7��rs������T��k�Ǥ%1�EV��r��_�**iK��e �i�/�n�<H#K>��E{�����~|V(��5�jt����؅�<1��r�>��İ�uF�g��+�5���z��;:���jRG]i�X[WV�X����:(C��䗎���l5�����@�.i���ء�*��"Oe{�,�+4�Wu~~�q��B�� ~n��nK��.��n4����Ǜ�a�X.�֍�уe���ʄ�"9��;���T|wUr�0���(} �_�ibq[��c��^Ө�$B2�GB��?"/��q�{_�i��	���v;e�!�����A�9�lCr�7��|���qW� ��
D/Y�N��D7u��C��lE ��j�3�F���4n���<����gO�����9qp]v%ڴ�XY�}�E�a	�Ve����t�-ga:0j�M�a��-wrв�+���+��b9�ӿ���b/��R�B�gx�B[�Ť��*�ف���4�������/��^_�UaA�B���R��([0��Te�n���/+�{����/^��it�n�����Qt8)�j�\�L�"ef˛ 8�-������}������Լ�;x�/F��M��%Y�����樷�W]�.���o8�O��(�z��?97������n�8~��0c�E��W�xFbG�W֮"敿���N:����L*4�5k�yz'U�G.��N&An�#��Jd�`��Q���Qy]��ٸUrOm�jk��92lW��^Vf�Ԃ�H)$�'����ɔ��Id���ᑪ\�T�<ęv�N�e�����M���a\�.�K�R��b}[$#�&-�K�=t��Z�d�67��ɁSv�m��0K�_-g�Z$JC��n����h%D�����R�~ࣅ�PSL�$���Eǋ�O\�#���ؾ���_�C�����3�&Ⱥx#P|����խc�9�$$N�U�Ra`�����y���%`�k��ۀ�:��H'Ҳ�%0!��k�ݮ��~���İB�\+^:��6��G������x`/��0�v�!�{̣�Zj�J5V�%-"�/��&�M�ͧ�.�m�LA��N:Ssͧ<����1�`�(Rce~���0 �wCI��#^G��SF.����b��"ϖ���N#;��K�Ù�A���0����d�L�|I�f�>Y{¹|��w��JJ��+�f�kf�0�U��n꺺y��G$���z'R��/<��B}X�J��RG�`>ɔ�Lp�;����
QJ IF��X2dCSx��_#��T��ϻu�g�/���Ӥ��W��������m �[TJ���]�������7����_+���_/�NPܼ�&>�͐���h1��p썌����Y?_��뢪�+j�r��9�8� �5M�T%PT\h�c�Q�-�->��i��-�Ǳ?��3]��|�*\����~3_���3'�ڕ��..��;?�?�p9*�Ȫ�����b��cB@���@�t��v��#1�r��]�|��f�r��D�;�\�
�!!�.,�O�̃���t3 Y�R��hj����@�mZ��(�@�:+C� ͮ$6��@����"��a� v~�0��+5�~G��մ�y����n)	��O��|@�uǳm{=^�GLMjU6�m� M�O,RH���}�ʮ.�q2���VL��:sؖ@� �>N^�u����Lj���JR��:���l:6�66?F�r0O=�,Ֆ�5��K���<�-�t02Zgq�m���M����c$�$IYm+��\P~ k��C�f����1�p��	�Q���˰J�p�o��^��8�o���5c2[�f�@�n�����H�h�4�d��'��Ws�����)��VDHi^2u�j)N6_ʑ|"�X����Bu���iFa����������-��8u�Yj:�oH#��5D��я�XB����X�.�®��*��b�Y��v@�p�Q�0 �X�)��y9�-X�+�k؊�kS2�f4�Y��a��9���|d(��|W^���� ��#HDŁ�'EX�xc��YX-f'�A�Q*���6�Qo��d�p��� �+�S!�,��������S���,pɖ�0HC�:�9�S���V�4�Ӝ2%T��meY�
/�^SF�]y����B�����߽<_8	��k���� �W�����u�S�E���sr�D���e=$�Q�$-s�.�(������W�H�UR�ëC9t<?�m�e.|n����}z��=����kbH=vB��g�y��r���D5:��V�S\nԙ9X���r�8�*�ĸjO�Ig'gg������y{�$A�A� b2�ܼ�z�хP�������Y7oF3E��#�&��L�Ϩ�m�uܯ�k<�9�ankkHH#��kX���j;� G$/�/��~�Z{����n��&�Z��u��@E�/ڧ`y;F�M�i�����X[�>�������X@��v�ڥ��'St��g��Zy��g�>��%�n,I%f����{i��٬x�dv��:\���'�>�JaK8B�t*�8�⏰��j,�Ȯ��X2+������$�Q�zU�-�����}nKE`��[��nUpџ�/�j�>%�_��IɄ�\I��Tb���+�� ��a�,�p���w�S?��%=�����ܹo�5�v�s��A���.p�c���M���s��!�N�rI/=O;��)^a���]�>��B��J2.�~�D�������`E���/|/���q�g��;%I�_����S'#E�inh�=�.�)�u�}�'���"1��޹�3���'�n�����LJSH��<7 ʞ2����.rg�)*gb��C1�K`��y*J��>Aq�[��r�א�\w�1=[�n�e�#ќZ�[T��1h����ڥ3+�����d���By�e8�E;�E��R�_k �K6�?�3���#��},����%�u�c�-ʼq.�z�#�ʡLb�2|�U}�"��𮍐�����_��״�u�T{��V��h9�J���Q<�CL����J�j@�{?��Y}�҄=��"4{�ߚ��,����5�:LnM�^��P7Csm"l4�J�(rÚ�_��D�KWyr�R�L|�ï���� Ԯݩ�n�xhc��_�N{����U��fI��l ?���艿�� b4���
���3\4��Z��.Ō8)�<��m0f_4:�M�;mI�FM��?U?�r�3�sFF{s�I��>�!ѐ�[��������iP�c������ռD���1�B�Z��F=�6F���͏5�:�R&`�wC{x"�B� ����2ʩ^7�$q�M}.Dp?���Śh�
$=���s_�}�6�����"�|;e!���^����4@���)z�U��}{���@��s>���h!!����V�%��?~���@�Do�c��*���kt�S<aF��
!�Ϝ'mƋQ&�E�Z�gu	׋C0��jQ�ϖ��\`�.A�e�#�%}R�RA� .N��z�(� A���Z�2�@�;�2s���0߸=���l��ϐ-fr_���^F��0|I���D����"}UR�)Gs�j|�a�l|_�\��e��AG
��!@��e��*2��ґ1���<��M;��n����9�qa�b7&��)o>.kq���=�m�'�i����?����_W�[��b"�qG���0E��C���}� ��G���U-n -��C�ɪi)����u�´*����z�o��4�7W$,�:�m�S#k�ȉX]�w��Z{�mr;�L�a+<�g�c?ӥn���Z$7B�^�-o�9A�)P��)� J��ym�&{���]㤲�(zJPOX/�a7\�����R��;=�_	lv�]*�^%�ʙ/`a~' &m�2��[������%�?Z��{V�����in�����T�E��u*y���Ā>_=����!
�܌{us3q����(:�! \���3���ܵ���V��z�`�<h�3~mڃ�6�i:�h����XP'UF����<�|%���ʰ0���U	q8�����u͒~�r�$d�@
���Ip������h&�_b!%�Hf��O��7mW��k�V�^zF:rg��Kt�8M�����ԅ������NBFc�����fVrV{`�"�x��\vY-�B���'�&`��'I5k�e(��o�	mH(�{���	�F�/7c�v�"��0�K �<��>Z���O�X�rKhx�B���\���q�����*ch�#S�@���`��Ը��ʄ���3�^S�0�y��M�y��|X�sY�d��V��\a��`$�c!�I���f����}���??�v��� ����'�a�$�?;��?[�N��G	�7\l�'��<D��V�Q@�jVp�M&�C?�B��Z0^Qܴ�%S�����i�x?)����eH��z�
|gB�k&��[I![c�����+ȥ��-�EvF�*�f�v<�_h�K%��νBh������	����M�A��%��*+Msq���R������Z��D9%,B�؇Y�ș�
3���s��7E�|i�l_�Y]@e�®��{Yuu�j�#��*����^ze�˂����npA>�E�<��Zr�2�u������--�D,����e�PJ$&V������K�9�����[�(7\@n��g��i�V���6f�(����
>��B��ry�Va�*V��n�ö�~�|����7�'�O��$�������A��CGQ��,�_(��ԟ��@7�������hB�Kci��[f�'<�]6DNwV)��~�Y���]�}%I��S�^�-��b�����)2X���ƋϞ�����?��R~���נ83���K��
 ��lef��K�ߚ�)(�S�k�,%"SN���<,�Ũ��]C�Et͋�n��NϼFUZ`1��(WR=2)�6�z=a^+5	*[�㍺;���BO���A��<�Pc�R�}�m����3�/��2� c�����o�q�n�v6�S���I� ���5�r��G��7� RU�C�!�	�{���ҳus���x4��X�2����У�FǑ��ճ2^�L��i��#�_��x���x&������$���j���"ڼOAT/t���t�eY\ +;�8�ݭ�f��G[���;�c�fc�~�Wk@:�\̜x��}9��9T����m�r���kPɜlV�*�L�Ey��Ї� ��������+��b��^F����b���nۇxsA��ɋ2,��F�����h�&�z軙9�*�R�%)��]�nO��0	� \������ƨ�2���ȝ���������y�Qb��$�Z��c��c�@�x�3N^�}�Tٚ��?nk�܏�mP�_\�$n�����&�X�>����.��K]3�<z�G�z5��o�r��*�Ń�QW@n��r؛�N8cA%Bpw��-t��;D�F|�ӘG�%������c&�P���Yh��&xOU��Ʈ/5Y����ߴ�s��4�����b��=^*OJ�����ۇ՘*'lÂaV���
��t����]�6}j�k���~�.Y�����ht�P3��fJ�׻�w	�Ai� �����]�3�c��������;�_�K����%���Ɇ�&6r��G�H>�eY�Q+�vf[8߮Ⴆ�ά�|���;��z5d�Z����;�4=z��S��㴥IG��p�C�(\��|�K+�=�?f�Y�R��|ۧj4�j)�lBi5����x���ߋ?'�U�{2!/6�