//------------------------------------------------------------
// Project: HYBRID_CONTROL
// Author: Nicola Zaupa
// Date: (2021/01/16) (21:43:22)
// File: trigonometry.v
//------------------------------------------------------------
// Description:
//
// Compuation of sine and cosine of an angle [0,pi]
// angle  x 100
// output x 1000
//------------------------------------------------------------


`timescale 1 ns / 1 ps
//`default_nettype none


module trigonometry (
   o_cos,    // cosine of the input
   o_sin,    // sine of the input
   i_theta   // input angle
);

output  signed [31:0] o_sin;
output  signed [31:0] o_cos;
input   signed [31:0] i_theta;

wire [31:0] o_sin;
wire [31:0] o_cos;
wire [31:0] i_theta;

reg [31:0] r_sin;
reg [31:0] r_cos;

assign o_sin = r_sin;
assign o_cos = r_cos;


always @ ( i_theta )
begin

// computation of sine and cosine using integers
// taking advanatges of look-up-table
// input angle is multiplied by x100
// trigonometric output is multiplied by x1000

case(i_theta)
      32'h00000000: r_sin = 32'h00000000;
      32'h00000001: r_sin = 32'h0000000A;
      32'h00000002: r_sin = 32'h00000014;
      32'h00000003: r_sin = 32'h0000001E;
      32'h00000004: r_sin = 32'h00000028;
      32'h00000005: r_sin = 32'h00000032;
      32'h00000006: r_sin = 32'h0000003C;
      32'h00000007: r_sin = 32'h00000046;
      32'h00000008: r_sin = 32'h00000050;
      32'h00000009: r_sin = 32'h0000005A;
      32'h0000000A: r_sin = 32'h00000064;
      32'h0000000B: r_sin = 32'h0000006E;
      32'h0000000C: r_sin = 32'h00000078;
      32'h0000000D: r_sin = 32'h00000082;
      32'h0000000E: r_sin = 32'h0000008C;
      32'h0000000F: r_sin = 32'h00000095;
      32'h00000010: r_sin = 32'h0000009F;
      32'h00000011: r_sin = 32'h000000A9;
      32'h00000012: r_sin = 32'h000000B3;
      32'h00000013: r_sin = 32'h000000BD;
      32'h00000014: r_sin = 32'h000000C7;
      32'h00000015: r_sin = 32'h000000D0;
      32'h00000016: r_sin = 32'h000000DA;
      32'h00000017: r_sin = 32'h000000E4;
      32'h00000018: r_sin = 32'h000000EE;
      32'h00000019: r_sin = 32'h000000F7;
      32'h0000001A: r_sin = 32'h00000101;
      32'h0000001B: r_sin = 32'h0000010B;
      32'h0000001C: r_sin = 32'h00000114;
      32'h0000001D: r_sin = 32'h0000011E;
      32'h0000001E: r_sin = 32'h00000128;
      32'h0000001F: r_sin = 32'h00000131;
      32'h00000020: r_sin = 32'h0000013B;
      32'h00000021: r_sin = 32'h00000144;
      32'h00000022: r_sin = 32'h0000014D;
      32'h00000023: r_sin = 32'h00000157;
      32'h00000024: r_sin = 32'h00000160;
      32'h00000025: r_sin = 32'h0000016A;
      32'h00000026: r_sin = 32'h00000173;
      32'h00000027: r_sin = 32'h0000017C;
      32'h00000028: r_sin = 32'h00000185;
      32'h00000029: r_sin = 32'h0000018F;
      32'h0000002A: r_sin = 32'h00000198;
      32'h0000002B: r_sin = 32'h000001A1;
      32'h0000002C: r_sin = 32'h000001AA;
      32'h0000002D: r_sin = 32'h000001B3;
      32'h0000002E: r_sin = 32'h000001BC;
      32'h0000002F: r_sin = 32'h000001C5;
      32'h00000030: r_sin = 32'h000001CE;
      32'h00000031: r_sin = 32'h000001D7;
      32'h00000032: r_sin = 32'h000001DF;
      32'h00000033: r_sin = 32'h000001E8;
      32'h00000034: r_sin = 32'h000001F1;
      32'h00000035: r_sin = 32'h000001FA;
      32'h00000036: r_sin = 32'h00000202;
      32'h00000037: r_sin = 32'h0000020B;
      32'h00000038: r_sin = 32'h00000213;
      32'h00000039: r_sin = 32'h0000021C;
      32'h0000003A: r_sin = 32'h00000224;
      32'h0000003B: r_sin = 32'h0000022C;
      32'h0000003C: r_sin = 32'h00000235;
      32'h0000003D: r_sin = 32'h0000023D;
      32'h0000003E: r_sin = 32'h00000245;
      32'h0000003F: r_sin = 32'h0000024D;
      32'h00000040: r_sin = 32'h00000255;
      32'h00000041: r_sin = 32'h0000025D;
      32'h00000042: r_sin = 32'h00000265;
      32'h00000043: r_sin = 32'h0000026D;
      32'h00000044: r_sin = 32'h00000275;
      32'h00000045: r_sin = 32'h0000027D;
      32'h00000046: r_sin = 32'h00000284;
      32'h00000047: r_sin = 32'h0000028C;
      32'h00000048: r_sin = 32'h00000293;
      32'h00000049: r_sin = 32'h0000029B;
      32'h0000004A: r_sin = 32'h000002A2;
      32'h0000004B: r_sin = 32'h000002AA;
      32'h0000004C: r_sin = 32'h000002B1;
      32'h0000004D: r_sin = 32'h000002B8;
      32'h0000004E: r_sin = 32'h000002BF;
      32'h0000004F: r_sin = 32'h000002C6;
      32'h00000050: r_sin = 32'h000002CD;
      32'h00000051: r_sin = 32'h000002D4;
      32'h00000052: r_sin = 32'h000002DB;
      32'h00000053: r_sin = 32'h000002E2;
      32'h00000054: r_sin = 32'h000002E9;
      32'h00000055: r_sin = 32'h000002EF;
      32'h00000056: r_sin = 32'h000002F6;
      32'h00000057: r_sin = 32'h000002FC;
      32'h00000058: r_sin = 32'h00000303;
      32'h00000059: r_sin = 32'h00000309;
      32'h0000005A: r_sin = 32'h0000030F;
      32'h0000005B: r_sin = 32'h00000316;
      32'h0000005C: r_sin = 32'h0000031C;
      32'h0000005D: r_sin = 32'h00000322;
      32'h0000005E: r_sin = 32'h00000328;
      32'h0000005F: r_sin = 32'h0000032D;
      32'h00000060: r_sin = 32'h00000333;
      32'h00000061: r_sin = 32'h00000339;
      32'h00000062: r_sin = 32'h0000033E;
      32'h00000063: r_sin = 32'h00000344;
      32'h00000064: r_sin = 32'h00000349;
      32'h00000065: r_sin = 32'h0000034F;
      32'h00000066: r_sin = 32'h00000354;
      32'h00000067: r_sin = 32'h00000359;
      32'h00000068: r_sin = 32'h0000035E;
      32'h00000069: r_sin = 32'h00000363;
      32'h0000006A: r_sin = 32'h00000368;
      32'h0000006B: r_sin = 32'h0000036D;
      32'h0000006C: r_sin = 32'h00000372;
      32'h0000006D: r_sin = 32'h00000377;
      32'h0000006E: r_sin = 32'h0000037B;
      32'h0000006F: r_sin = 32'h00000380;
      32'h00000070: r_sin = 32'h00000384;
      32'h00000071: r_sin = 32'h00000388;
      32'h00000072: r_sin = 32'h0000038D;
      32'h00000073: r_sin = 32'h00000391;
      32'h00000074: r_sin = 32'h00000395;
      32'h00000075: r_sin = 32'h00000399;
      32'h00000076: r_sin = 32'h0000039D;
      32'h00000077: r_sin = 32'h000003A0;
      32'h00000078: r_sin = 32'h000003A4;
      32'h00000079: r_sin = 32'h000003A8;
      32'h0000007A: r_sin = 32'h000003AB;
      32'h0000007B: r_sin = 32'h000003AE;
      32'h0000007C: r_sin = 32'h000003B2;
      32'h0000007D: r_sin = 32'h000003B5;
      32'h0000007E: r_sin = 32'h000003B8;
      32'h0000007F: r_sin = 32'h000003BB;
      32'h00000080: r_sin = 32'h000003BE;
      32'h00000081: r_sin = 32'h000003C1;
      32'h00000082: r_sin = 32'h000003C4;
      32'h00000083: r_sin = 32'h000003C6;
      32'h00000084: r_sin = 32'h000003C9;
      32'h00000085: r_sin = 32'h000003CB;
      32'h00000086: r_sin = 32'h000003CD;
      32'h00000087: r_sin = 32'h000003D0;
      32'h00000088: r_sin = 32'h000003D2;
      32'h00000089: r_sin = 32'h000003D4;
      32'h0000008A: r_sin = 32'h000003D6;
      32'h0000008B: r_sin = 32'h000003D8;
      32'h0000008C: r_sin = 32'h000003D9;
      32'h0000008D: r_sin = 32'h000003DB;
      32'h0000008E: r_sin = 32'h000003DD;
      32'h0000008F: r_sin = 32'h000003DE;
      32'h00000090: r_sin = 32'h000003DF;
      32'h00000091: r_sin = 32'h000003E1;
      32'h00000092: r_sin = 32'h000003E2;
      32'h00000093: r_sin = 32'h000003E3;
      32'h00000094: r_sin = 32'h000003E4;
      32'h00000095: r_sin = 32'h000003E5;
      32'h00000096: r_sin = 32'h000003E5;
      32'h00000097: r_sin = 32'h000003E6;
      32'h00000098: r_sin = 32'h000003E7;
      32'h00000099: r_sin = 32'h000003E7;
      32'h0000009A: r_sin = 32'h000003E8;
      32'h0000009B: r_sin = 32'h000003E8;
      32'h0000009C: r_sin = 32'h000003E8;
      32'h0000009D: r_sin = 32'h000003E8;
      32'h0000009E: r_sin = 32'h000003E8;
      32'h0000009F: r_sin = 32'h000003E8;
      32'h000000A0: r_sin = 32'h000003E8;
      32'h000000A1: r_sin = 32'h000003E7;
      32'h000000A2: r_sin = 32'h000003E7;
      32'h000000A3: r_sin = 32'h000003E6;
      32'h000000A4: r_sin = 32'h000003E6;
      32'h000000A5: r_sin = 32'h000003E5;
      32'h000000A6: r_sin = 32'h000003E4;
      32'h000000A7: r_sin = 32'h000003E3;
      32'h000000A8: r_sin = 32'h000003E2;
      32'h000000A9: r_sin = 32'h000003E1;
      32'h000000AA: r_sin = 32'h000003E0;
      32'h000000AB: r_sin = 32'h000003DE;
      32'h000000AC: r_sin = 32'h000003DD;
      32'h000000AD: r_sin = 32'h000003DB;
      32'h000000AE: r_sin = 32'h000003DA;
      32'h000000AF: r_sin = 32'h000003D8;
      32'h000000B0: r_sin = 32'h000003D6;
      32'h000000B1: r_sin = 32'h000003D4;
      32'h000000B2: r_sin = 32'h000003D2;
      32'h000000B3: r_sin = 32'h000003D0;
      32'h000000B4: r_sin = 32'h000003CE;
      32'h000000B5: r_sin = 32'h000003CC;
      32'h000000B6: r_sin = 32'h000003C9;
      32'h000000B7: r_sin = 32'h000003C7;
      32'h000000B8: r_sin = 32'h000003C4;
      32'h000000B9: r_sin = 32'h000003C1;
      32'h000000BA: r_sin = 32'h000003BE;
      32'h000000BB: r_sin = 32'h000003BC;
      32'h000000BC: r_sin = 32'h000003B9;
      32'h000000BD: r_sin = 32'h000003B5;
      32'h000000BE: r_sin = 32'h000003B2;
      32'h000000BF: r_sin = 32'h000003AF;
      32'h000000C0: r_sin = 32'h000003AC;
      32'h000000C1: r_sin = 32'h000003A8;
      32'h000000C2: r_sin = 32'h000003A5;
      32'h000000C3: r_sin = 32'h000003A1;
      32'h000000C4: r_sin = 32'h0000039D;
      32'h000000C5: r_sin = 32'h00000399;
      32'h000000C6: r_sin = 32'h00000395;
      32'h000000C7: r_sin = 32'h00000391;
      32'h000000C8: r_sin = 32'h0000038D;
      32'h000000C9: r_sin = 32'h00000389;
      32'h000000CA: r_sin = 32'h00000385;
      32'h000000CB: r_sin = 32'h00000380;
      32'h000000CC: r_sin = 32'h0000037C;
      32'h000000CD: r_sin = 32'h00000377;
      32'h000000CE: r_sin = 32'h00000373;
      32'h000000CF: r_sin = 32'h0000036E;
      32'h000000D0: r_sin = 32'h00000369;
      32'h000000D1: r_sin = 32'h00000364;
      32'h000000D2: r_sin = 32'h0000035F;
      32'h000000D3: r_sin = 32'h0000035A;
      32'h000000D4: r_sin = 32'h00000355;
      32'h000000D5: r_sin = 32'h00000350;
      32'h000000D6: r_sin = 32'h0000034A;
      32'h000000D7: r_sin = 32'h00000345;
      32'h000000D8: r_sin = 32'h0000033F;
      32'h000000D9: r_sin = 32'h0000033A;
      32'h000000DA: r_sin = 32'h00000334;
      32'h000000DB: r_sin = 32'h0000032E;
      32'h000000DC: r_sin = 32'h00000328;
      32'h000000DD: r_sin = 32'h00000323;
      32'h000000DE: r_sin = 32'h0000031D;
      32'h000000DF: r_sin = 32'h00000316;
      32'h000000E0: r_sin = 32'h00000310;
      32'h000000E1: r_sin = 32'h0000030A;
      32'h000000E2: r_sin = 32'h00000304;
      32'h000000E3: r_sin = 32'h000002FD;
      32'h000000E4: r_sin = 32'h000002F7;
      32'h000000E5: r_sin = 32'h000002F0;
      32'h000000E6: r_sin = 32'h000002EA;
      32'h000000E7: r_sin = 32'h000002E3;
      32'h000000E8: r_sin = 32'h000002DC;
      32'h000000E9: r_sin = 32'h000002D5;
      32'h000000EA: r_sin = 32'h000002CE;
      32'h000000EB: r_sin = 32'h000002C7;
      32'h000000EC: r_sin = 32'h000002C0;
      32'h000000ED: r_sin = 32'h000002B9;
      32'h000000EE: r_sin = 32'h000002B2;
      32'h000000EF: r_sin = 32'h000002AB;
      32'h000000F0: r_sin = 32'h000002A3;
      32'h000000F1: r_sin = 32'h0000029C;
      32'h000000F2: r_sin = 32'h00000295;
      32'h000000F3: r_sin = 32'h0000028D;
      32'h000000F4: r_sin = 32'h00000285;
      32'h000000F5: r_sin = 32'h0000027E;
      32'h000000F6: r_sin = 32'h00000276;
      32'h000000F7: r_sin = 32'h0000026E;
      32'h000000F8: r_sin = 32'h00000266;
      32'h000000F9: r_sin = 32'h0000025E;
      32'h000000FA: r_sin = 32'h00000256;
      32'h000000FB: r_sin = 32'h0000024E;
      32'h000000FC: r_sin = 32'h00000246;
      32'h000000FD: r_sin = 32'h0000023E;
      32'h000000FE: r_sin = 32'h00000236;
      32'h000000FF: r_sin = 32'h0000022E;
      32'h00000100: r_sin = 32'h00000225;
      32'h00000101: r_sin = 32'h0000021D;
      32'h00000102: r_sin = 32'h00000215;
      32'h00000103: r_sin = 32'h0000020C;
      32'h00000104: r_sin = 32'h00000204;
      32'h00000105: r_sin = 32'h000001FB;
      32'h00000106: r_sin = 32'h000001F2;
      32'h00000107: r_sin = 32'h000001EA;
      32'h00000108: r_sin = 32'h000001E1;
      32'h00000109: r_sin = 32'h000001D8;
      32'h0000010A: r_sin = 32'h000001CF;
      32'h0000010B: r_sin = 32'h000001C6;
      32'h0000010C: r_sin = 32'h000001BD;
      32'h0000010D: r_sin = 32'h000001B4;
      32'h0000010E: r_sin = 32'h000001AB;
      32'h0000010F: r_sin = 32'h000001A2;
      32'h00000110: r_sin = 32'h00000199;
      32'h00000111: r_sin = 32'h00000190;
      32'h00000112: r_sin = 32'h00000187;
      32'h00000113: r_sin = 32'h0000017E;
      32'h00000114: r_sin = 32'h00000174;
      32'h00000115: r_sin = 32'h0000016B;
      32'h00000116: r_sin = 32'h00000162;
      32'h00000117: r_sin = 32'h00000158;
      32'h00000118: r_sin = 32'h0000014F;
      32'h00000119: r_sin = 32'h00000146;
      32'h0000011A: r_sin = 32'h0000013C;
      32'h0000011B: r_sin = 32'h00000133;
      32'h0000011C: r_sin = 32'h00000129;
      32'h0000011D: r_sin = 32'h0000011F;
      32'h0000011E: r_sin = 32'h00000116;
      32'h0000011F: r_sin = 32'h0000010C;
      32'h00000120: r_sin = 32'h00000103;
      32'h00000121: r_sin = 32'h000000F9;
      32'h00000122: r_sin = 32'h000000EF;
      32'h00000123: r_sin = 32'h000000E6;
      32'h00000124: r_sin = 32'h000000DC;
      32'h00000125: r_sin = 32'h000000D2;
      32'h00000126: r_sin = 32'h000000C8;
      32'h00000127: r_sin = 32'h000000BE;
      32'h00000128: r_sin = 32'h000000B5;
      32'h00000129: r_sin = 32'h000000AB;
      32'h0000012A: r_sin = 32'h000000A1;
      32'h0000012B: r_sin = 32'h00000097;
      32'h0000012C: r_sin = 32'h0000008D;
      32'h0000012D: r_sin = 32'h00000083;
      32'h0000012E: r_sin = 32'h00000079;
      32'h0000012F: r_sin = 32'h0000006F;
      32'h00000130: r_sin = 32'h00000065;
      32'h00000131: r_sin = 32'h0000005B;
      32'h00000132: r_sin = 32'h00000052;
      32'h00000133: r_sin = 32'h00000048;
      32'h00000134: r_sin = 32'h0000003E;
      32'h00000135: r_sin = 32'h00000034;
      32'h00000136: r_sin = 32'h0000002A;
      32'h00000137: r_sin = 32'h00000020;
      32'h00000138: r_sin = 32'h00000016;
      32'h00000139: r_sin = 32'h0000000C;
      32'h0000013A: r_sin = 32'h00000000;
      default: r_sin = 32'h00000000;
endcase

case(i_theta)
      32'h00000000: r_cos = 32'h000003E8;
      32'h00000001: r_cos = 32'h000003E8;
      32'h00000002: r_cos = 32'h000003E8;
      32'h00000003: r_cos = 32'h000003E8;
      32'h00000004: r_cos = 32'h000003E7;
      32'h00000005: r_cos = 32'h000003E7;
      32'h00000006: r_cos = 32'h000003E6;
      32'h00000007: r_cos = 32'h000003E6;
      32'h00000008: r_cos = 32'h000003E5;
      32'h00000009: r_cos = 32'h000003E4;
      32'h0000000A: r_cos = 32'h000003E3;
      32'h0000000B: r_cos = 32'h000003E2;
      32'h0000000C: r_cos = 32'h000003E1;
      32'h0000000D: r_cos = 32'h000003E0;
      32'h0000000E: r_cos = 32'h000003DE;
      32'h0000000F: r_cos = 32'h000003DD;
      32'h00000010: r_cos = 32'h000003DB;
      32'h00000011: r_cos = 32'h000003DA;
      32'h00000012: r_cos = 32'h000003D8;
      32'h00000013: r_cos = 32'h000003D6;
      32'h00000014: r_cos = 32'h000003D4;
      32'h00000015: r_cos = 32'h000003D2;
      32'h00000016: r_cos = 32'h000003D0;
      32'h00000017: r_cos = 32'h000003CE;
      32'h00000018: r_cos = 32'h000003CB;
      32'h00000019: r_cos = 32'h000003C9;
      32'h0000001A: r_cos = 32'h000003C6;
      32'h0000001B: r_cos = 32'h000003C4;
      32'h0000001C: r_cos = 32'h000003C1;
      32'h0000001D: r_cos = 32'h000003BE;
      32'h0000001E: r_cos = 32'h000003BB;
      32'h0000001F: r_cos = 32'h000003B8;
      32'h00000020: r_cos = 32'h000003B5;
      32'h00000021: r_cos = 32'h000003B2;
      32'h00000022: r_cos = 32'h000003AF;
      32'h00000023: r_cos = 32'h000003AB;
      32'h00000024: r_cos = 32'h000003A8;
      32'h00000025: r_cos = 32'h000003A4;
      32'h00000026: r_cos = 32'h000003A1;
      32'h00000027: r_cos = 32'h0000039D;
      32'h00000028: r_cos = 32'h00000399;
      32'h00000029: r_cos = 32'h00000395;
      32'h0000002A: r_cos = 32'h00000391;
      32'h0000002B: r_cos = 32'h0000038D;
      32'h0000002C: r_cos = 32'h00000389;
      32'h0000002D: r_cos = 32'h00000384;
      32'h0000002E: r_cos = 32'h00000380;
      32'h0000002F: r_cos = 32'h0000037C;
      32'h00000030: r_cos = 32'h00000377;
      32'h00000031: r_cos = 32'h00000372;
      32'h00000032: r_cos = 32'h0000036E;
      32'h00000033: r_cos = 32'h00000369;
      32'h00000034: r_cos = 32'h00000364;
      32'h00000035: r_cos = 32'h0000035F;
      32'h00000036: r_cos = 32'h0000035A;
      32'h00000037: r_cos = 32'h00000355;
      32'h00000038: r_cos = 32'h0000034F;
      32'h00000039: r_cos = 32'h0000034A;
      32'h0000003A: r_cos = 32'h00000344;
      32'h0000003B: r_cos = 32'h0000033F;
      32'h0000003C: r_cos = 32'h00000339;
      32'h0000003D: r_cos = 32'h00000334;
      32'h0000003E: r_cos = 32'h0000032E;
      32'h0000003F: r_cos = 32'h00000328;
      32'h00000040: r_cos = 32'h00000322;
      32'h00000041: r_cos = 32'h0000031C;
      32'h00000042: r_cos = 32'h00000316;
      32'h00000043: r_cos = 32'h00000310;
      32'h00000044: r_cos = 32'h0000030A;
      32'h00000045: r_cos = 32'h00000303;
      32'h00000046: r_cos = 32'h000002FD;
      32'h00000047: r_cos = 32'h000002F6;
      32'h00000048: r_cos = 32'h000002F0;
      32'h00000049: r_cos = 32'h000002E9;
      32'h0000004A: r_cos = 32'h000002E2;
      32'h0000004B: r_cos = 32'h000002DC;
      32'h0000004C: r_cos = 32'h000002D5;
      32'h0000004D: r_cos = 32'h000002CE;
      32'h0000004E: r_cos = 32'h000002C7;
      32'h0000004F: r_cos = 32'h000002C0;
      32'h00000050: r_cos = 32'h000002B9;
      32'h00000051: r_cos = 32'h000002B1;
      32'h00000052: r_cos = 32'h000002AA;
      32'h00000053: r_cos = 32'h000002A3;
      32'h00000054: r_cos = 32'h0000029B;
      32'h00000055: r_cos = 32'h00000294;
      32'h00000056: r_cos = 32'h0000028C;
      32'h00000057: r_cos = 32'h00000285;
      32'h00000058: r_cos = 32'h0000027D;
      32'h00000059: r_cos = 32'h00000275;
      32'h0000005A: r_cos = 32'h0000026E;
      32'h0000005B: r_cos = 32'h00000266;
      32'h0000005C: r_cos = 32'h0000025E;
      32'h0000005D: r_cos = 32'h00000256;
      32'h0000005E: r_cos = 32'h0000024E;
      32'h0000005F: r_cos = 32'h00000246;
      32'h00000060: r_cos = 32'h0000023E;
      32'h00000061: r_cos = 32'h00000235;
      32'h00000062: r_cos = 32'h0000022D;
      32'h00000063: r_cos = 32'h00000225;
      32'h00000064: r_cos = 32'h0000021C;
      32'h00000065: r_cos = 32'h00000214;
      32'h00000066: r_cos = 32'h0000020B;
      32'h00000067: r_cos = 32'h00000203;
      32'h00000068: r_cos = 32'h000001FA;
      32'h00000069: r_cos = 32'h000001F2;
      32'h0000006A: r_cos = 32'h000001E9;
      32'h0000006B: r_cos = 32'h000001E0;
      32'h0000006C: r_cos = 32'h000001D7;
      32'h0000006D: r_cos = 32'h000001CE;
      32'h0000006E: r_cos = 32'h000001C6;
      32'h0000006F: r_cos = 32'h000001BD;
      32'h00000070: r_cos = 32'h000001B4;
      32'h00000071: r_cos = 32'h000001AB;
      32'h00000072: r_cos = 32'h000001A2;
      32'h00000073: r_cos = 32'h00000198;
      32'h00000074: r_cos = 32'h0000018F;
      32'h00000075: r_cos = 32'h00000186;
      32'h00000076: r_cos = 32'h0000017D;
      32'h00000077: r_cos = 32'h00000174;
      32'h00000078: r_cos = 32'h0000016A;
      32'h00000079: r_cos = 32'h00000161;
      32'h0000007A: r_cos = 32'h00000158;
      32'h0000007B: r_cos = 32'h0000014E;
      32'h0000007C: r_cos = 32'h00000145;
      32'h0000007D: r_cos = 32'h0000013B;
      32'h0000007E: r_cos = 32'h00000132;
      32'h0000007F: r_cos = 32'h00000128;
      32'h00000080: r_cos = 32'h0000011F;
      32'h00000081: r_cos = 32'h00000115;
      32'h00000082: r_cos = 32'h0000010B;
      32'h00000083: r_cos = 32'h00000102;
      32'h00000084: r_cos = 32'h000000F8;
      32'h00000085: r_cos = 32'h000000EE;
      32'h00000086: r_cos = 32'h000000E5;
      32'h00000087: r_cos = 32'h000000DB;
      32'h00000088: r_cos = 32'h000000D1;
      32'h00000089: r_cos = 32'h000000C7;
      32'h0000008A: r_cos = 32'h000000BE;
      32'h0000008B: r_cos = 32'h000000B4;
      32'h0000008C: r_cos = 32'h000000AA;
      32'h0000008D: r_cos = 32'h000000A0;
      32'h0000008E: r_cos = 32'h00000096;
      32'h0000008F: r_cos = 32'h0000008C;
      32'h00000090: r_cos = 32'h00000082;
      32'h00000091: r_cos = 32'h00000079;
      32'h00000092: r_cos = 32'h0000006F;
      32'h00000093: r_cos = 32'h00000065;
      32'h00000094: r_cos = 32'h0000005B;
      32'h00000095: r_cos = 32'h00000051;
      32'h00000096: r_cos = 32'h00000047;
      32'h00000097: r_cos = 32'h0000003D;
      32'h00000098: r_cos = 32'h00000033;
      32'h00000099: r_cos = 32'h00000029;
      32'h0000009A: r_cos = 32'h0000001F;
      32'h0000009B: r_cos = 32'h00000015;
      32'h0000009C: r_cos = 32'h0000000B;
      32'h0000009D: r_cos = 32'h00000001;
      32'h0000009E: r_cos = 32'hFFFFFFF7;
      32'h0000009F: r_cos = 32'hFFFFFFED;
      32'h000000A0: r_cos = 32'hFFFFFFE3;
      32'h000000A1: r_cos = 32'hFFFFFFD9;
      32'h000000A2: r_cos = 32'hFFFFFFCF;
      32'h000000A3: r_cos = 32'hFFFFFFC5;
      32'h000000A4: r_cos = 32'hFFFFFFBB;
      32'h000000A5: r_cos = 32'hFFFFFFB1;
      32'h000000A6: r_cos = 32'hFFFFFFA7;
      32'h000000A7: r_cos = 32'hFFFFFF9D;
      32'h000000A8: r_cos = 32'hFFFFFF93;
      32'h000000A9: r_cos = 32'hFFFFFF89;
      32'h000000AA: r_cos = 32'hFFFFFF7F;
      32'h000000AB: r_cos = 32'hFFFFFF75;
      32'h000000AC: r_cos = 32'hFFFFFF6B;
      32'h000000AD: r_cos = 32'hFFFFFF61;
      32'h000000AE: r_cos = 32'hFFFFFF58;
      32'h000000AF: r_cos = 32'hFFFFFF4E;
      32'h000000B0: r_cos = 32'hFFFFFF44;
      32'h000000B1: r_cos = 32'hFFFFFF3A;
      32'h000000B2: r_cos = 32'hFFFFFF30;
      32'h000000B3: r_cos = 32'hFFFFFF27;
      32'h000000B4: r_cos = 32'hFFFFFF1D;
      32'h000000B5: r_cos = 32'hFFFFFF13;
      32'h000000B6: r_cos = 32'hFFFFFF09;
      32'h000000B7: r_cos = 32'hFFFFFF00;
      32'h000000B8: r_cos = 32'hFFFFFEF6;
      32'h000000B9: r_cos = 32'hFFFFFEEC;
      32'h000000BA: r_cos = 32'hFFFFFEE3;
      32'h000000BB: r_cos = 32'hFFFFFED9;
      32'h000000BC: r_cos = 32'hFFFFFED0;
      32'h000000BD: r_cos = 32'hFFFFFEC6;
      32'h000000BE: r_cos = 32'hFFFFFEBD;
      32'h000000BF: r_cos = 32'hFFFFFEB3;
      32'h000000C0: r_cos = 32'hFFFFFEAA;
      32'h000000C1: r_cos = 32'hFFFFFEA0;
      32'h000000C2: r_cos = 32'hFFFFFE97;
      32'h000000C3: r_cos = 32'hFFFFFE8E;
      32'h000000C4: r_cos = 32'hFFFFFE85;
      32'h000000C5: r_cos = 32'hFFFFFE7B;
      32'h000000C6: r_cos = 32'hFFFFFE72;
      32'h000000C7: r_cos = 32'hFFFFFE69;
      32'h000000C8: r_cos = 32'hFFFFFE60;
      32'h000000C9: r_cos = 32'hFFFFFE57;
      32'h000000CA: r_cos = 32'hFFFFFE4E;
      32'h000000CB: r_cos = 32'hFFFFFE45;
      32'h000000CC: r_cos = 32'hFFFFFE3C;
      32'h000000CD: r_cos = 32'hFFFFFE33;
      32'h000000CE: r_cos = 32'hFFFFFE2A;
      32'h000000CF: r_cos = 32'hFFFFFE21;
      32'h000000D0: r_cos = 32'hFFFFFE19;
      32'h000000D1: r_cos = 32'hFFFFFE10;
      32'h000000D2: r_cos = 32'hFFFFFE07;
      32'h000000D3: r_cos = 32'hFFFFFDFF;
      32'h000000D4: r_cos = 32'hFFFFFDF6;
      32'h000000D5: r_cos = 32'hFFFFFDED;
      32'h000000D6: r_cos = 32'hFFFFFDE5;
      32'h000000D7: r_cos = 32'hFFFFFDDD;
      32'h000000D8: r_cos = 32'hFFFFFDD4;
      32'h000000D9: r_cos = 32'hFFFFFDCC;
      32'h000000DA: r_cos = 32'hFFFFFDC4;
      32'h000000DB: r_cos = 32'hFFFFFDBC;
      32'h000000DC: r_cos = 32'hFFFFFDB3;
      32'h000000DD: r_cos = 32'hFFFFFDAB;
      32'h000000DE: r_cos = 32'hFFFFFDA3;
      32'h000000DF: r_cos = 32'hFFFFFD9C;
      32'h000000E0: r_cos = 32'hFFFFFD94;
      32'h000000E1: r_cos = 32'hFFFFFD8C;
      32'h000000E2: r_cos = 32'hFFFFFD84;
      32'h000000E3: r_cos = 32'hFFFFFD7C;
      32'h000000E4: r_cos = 32'hFFFFFD75;
      32'h000000E5: r_cos = 32'hFFFFFD6D;
      32'h000000E6: r_cos = 32'hFFFFFD66;
      32'h000000E7: r_cos = 32'hFFFFFD5E;
      32'h000000E8: r_cos = 32'hFFFFFD57;
      32'h000000E9: r_cos = 32'hFFFFFD50;
      32'h000000EA: r_cos = 32'hFFFFFD48;
      32'h000000EB: r_cos = 32'hFFFFFD41;
      32'h000000EC: r_cos = 32'hFFFFFD3A;
      32'h000000ED: r_cos = 32'hFFFFFD33;
      32'h000000EE: r_cos = 32'hFFFFFD2C;
      32'h000000EF: r_cos = 32'hFFFFFD25;
      32'h000000F0: r_cos = 32'hFFFFFD1F;
      32'h000000F1: r_cos = 32'hFFFFFD18;
      32'h000000F2: r_cos = 32'hFFFFFD11;
      32'h000000F3: r_cos = 32'hFFFFFD0B;
      32'h000000F4: r_cos = 32'hFFFFFD04;
      32'h000000F5: r_cos = 32'hFFFFFCFE;
      32'h000000F6: r_cos = 32'hFFFFFCF7;
      32'h000000F7: r_cos = 32'hFFFFFCF1;
      32'h000000F8: r_cos = 32'hFFFFFCEB;
      32'h000000F9: r_cos = 32'hFFFFFCE5;
      32'h000000FA: r_cos = 32'hFFFFFCDF;
      32'h000000FB: r_cos = 32'hFFFFFCD9;
      32'h000000FC: r_cos = 32'hFFFFFCD3;
      32'h000000FD: r_cos = 32'hFFFFFCCD;
      32'h000000FE: r_cos = 32'hFFFFFCC8;
      32'h000000FF: r_cos = 32'hFFFFFCC2;
      32'h00000100: r_cos = 32'hFFFFFCBC;
      32'h00000101: r_cos = 32'hFFFFFCB7;
      32'h00000102: r_cos = 32'hFFFFFCB2;
      32'h00000103: r_cos = 32'hFFFFFCAC;
      32'h00000104: r_cos = 32'hFFFFFCA7;
      32'h00000105: r_cos = 32'hFFFFFCA2;
      32'h00000106: r_cos = 32'hFFFFFC9D;
      32'h00000107: r_cos = 32'hFFFFFC98;
      32'h00000108: r_cos = 32'hFFFFFC93;
      32'h00000109: r_cos = 32'hFFFFFC8E;
      32'h0000010A: r_cos = 32'hFFFFFC8A;
      32'h0000010B: r_cos = 32'hFFFFFC85;
      32'h0000010C: r_cos = 32'hFFFFFC81;
      32'h0000010D: r_cos = 32'hFFFFFC7C;
      32'h0000010E: r_cos = 32'hFFFFFC78;
      32'h0000010F: r_cos = 32'hFFFFFC74;
      32'h00000110: r_cos = 32'hFFFFFC70;
      32'h00000111: r_cos = 32'hFFFFFC6C;
      32'h00000112: r_cos = 32'hFFFFFC68;
      32'h00000113: r_cos = 32'hFFFFFC64;
      32'h00000114: r_cos = 32'hFFFFFC60;
      32'h00000115: r_cos = 32'hFFFFFC5C;
      32'h00000116: r_cos = 32'hFFFFFC59;
      32'h00000117: r_cos = 32'hFFFFFC55;
      32'h00000118: r_cos = 32'hFFFFFC52;
      32'h00000119: r_cos = 32'hFFFFFC4E;
      32'h0000011A: r_cos = 32'hFFFFFC4B;
      32'h0000011B: r_cos = 32'hFFFFFC48;
      32'h0000011C: r_cos = 32'hFFFFFC45;
      32'h0000011D: r_cos = 32'hFFFFFC42;
      32'h0000011E: r_cos = 32'hFFFFFC3F;
      32'h0000011F: r_cos = 32'hFFFFFC3D;
      32'h00000120: r_cos = 32'hFFFFFC3A;
      32'h00000121: r_cos = 32'hFFFFFC37;
      32'h00000122: r_cos = 32'hFFFFFC35;
      32'h00000123: r_cos = 32'hFFFFFC33;
      32'h00000124: r_cos = 32'hFFFFFC30;
      32'h00000125: r_cos = 32'hFFFFFC2E;
      32'h00000126: r_cos = 32'hFFFFFC2C;
      32'h00000127: r_cos = 32'hFFFFFC2A;
      32'h00000128: r_cos = 32'hFFFFFC28;
      32'h00000129: r_cos = 32'hFFFFFC27;
      32'h0000012A: r_cos = 32'hFFFFFC25;
      32'h0000012B: r_cos = 32'hFFFFFC23;
      32'h0000012C: r_cos = 32'hFFFFFC22;
      32'h0000012D: r_cos = 32'hFFFFFC21;
      32'h0000012E: r_cos = 32'hFFFFFC1F;
      32'h0000012F: r_cos = 32'hFFFFFC1E;
      32'h00000130: r_cos = 32'hFFFFFC1D;
      32'h00000131: r_cos = 32'hFFFFFC1C;
      32'h00000132: r_cos = 32'hFFFFFC1B;
      32'h00000133: r_cos = 32'hFFFFFC1B;
      32'h00000134: r_cos = 32'hFFFFFC1A;
      32'h00000135: r_cos = 32'hFFFFFC19;
      32'h00000136: r_cos = 32'hFFFFFC19;
      32'h00000137: r_cos = 32'hFFFFFC18;
      32'h00000138: r_cos = 32'hFFFFFC18;
      32'h00000139: r_cos = 32'hFFFFFC18;
      32'h0000013A: r_cos = 32'hFFFFFC18;
      default: r_cos = 32'hFFFFFC18;
endcase

end


endmodule