//------------------------------------------------------------
// Project: HYBRID_CONTROL
// Author: Nicola Zaupa
// Date: (2021/01/16) (21:43:22)
// File: modelsim.v
//------------------------------------------------------------
// Description:
//
// Compuation of sine and cosine of an angle [0,pi]
// angle  x 100
// output x 1000
//------------------------------------------------------------


`timescale 1 ns / 1 ps
`default_nettype none

module TOP_ResonantConverter_control_loop_tb;

reg          CLK;
reg          CLK_2;
reg          CLK_ADC;
reg          RESET;
reg          main_clk;
reg  [13:0]  SIGNAL_A;
reg  [13:0]  SIGNAL_B;
reg          OCR_A;
reg          OCR_B;

wire Q_POS;
wire Q_NEG;

reg            sigma;
reg    [13:0]  data_control;





TOP_ResonantConverter_control_loop TOP_ResonantConverter_control_loop_inst(
   .OSC        (CLK),
   .CLK_2      (CLK_2),
   .CPU_RESET  (RESET),
   //data + out-of-range
   .ADA_DATA(SIGNAL_A),
   .ADB_DATA(SIGNAL_B),
   .ADA_OR(),
   .ADB_OR(),
   .AD_SCLK(),
   .AD_SDIO(),
   .ADA_OE(),
   .ADA_SPI_CS(),
   .ADB_OE(),
   .ADB_SPI_CS(),
   .FPGA_CLK_A_N(),
   .FPGA_CLK_A_P(),
   .FPGA_CLK_B_N(),
   .FPGA_CLK_B_P(),
   .ADA_DCO(CLK_ADC),
   .ADB_DCO(CLK_ADC),
   // DAC
   .DA(),
   .DB(),
   //output bridge signal
   .OUT(),
   //debugging
   .BUTTON(),  // button on the main board
   .SW(),      // switches on the main board
   .LED(),     // LEDs on the main board
   .SEG0(),    // 7-segments display LSB
   .SEG1()
);





always
   begin
      CLK = 1'b1;
      #1.666;
      CLK = 1'b0;
      #1.666;
end

always
   begin
      CLK_2 = 1'b1;
      #5;
      CLK_2 = 1'b0;
      #5;
end


initial
   begin

RESET = 1'b1;

// samplings of current and voltage



CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110100;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b1111010111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111010111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000101;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010010;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111010110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101100;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111010110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101100;
SIGNAL_B = 14'b1111010110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b1111010110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b1111010100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b1111010011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100011111;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111001;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b1111001111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001010;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b1111001111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b1111001101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b1111001101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b1111001100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111110;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b1111001010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b1111001001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b1111001001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b1111001010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b1111001000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b1111001001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100001111;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100001111;
SIGNAL_B = 14'b1111000110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110110;
SIGNAL_B = 14'b1111000110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b1111000011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100001;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111010;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010100;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1111000001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b1111000001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b1111000000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100101;
SIGNAL_B = 14'b1110111110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010001010;
SIGNAL_B = 14'b1110111111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110001;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b1110111110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b1110111110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110011;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110011;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110011;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101000001;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111000011;
SIGNAL_B = 14'b1110111001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010001;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010000;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b1110111001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b1110110111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111111000;
SIGNAL_B = 14'b1110111000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101010;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011111;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b1110110111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001011111;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b1110110111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b1110110110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b1110110101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001001;
SIGNAL_B = 14'b1110110100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001010;
SIGNAL_B = 14'b1110110011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b1110110011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010110;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111110;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b1110110011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101011000;
SIGNAL_B = 14'b1110110010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110011001;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b1110110001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110011001;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111100111;
SIGNAL_B = 14'b1110110000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b1110101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011011;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001011101;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110101;
SIGNAL_B = 14'b1110101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b1110101111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110110;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010011;
SIGNAL_B = 14'b1110101111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010011;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010011;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111010;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111001;
SIGNAL_B = 14'b1110101011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111010;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111011;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010011;
SIGNAL_B = 14'b1110101011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010100;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010111;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111011000;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111100100;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b1110101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b1110100111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001110;
SIGNAL_B = 14'b1110101000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b1110101000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010011011;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010011011;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011001111;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011110110;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100101010;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101010010;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000101;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000100;
SIGNAL_B = 14'b1110100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b1110100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101011;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000110;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b1110100011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b1110100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001001;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001001;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000110000;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b1110100010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b1110100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001100;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b1110100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b1110100000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001101;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011000;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001111;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110010000;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110001111;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111111001;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111111000;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b1110011101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010010;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010100;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010100;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100011;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100100;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001011;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100011;
SIGNAL_B = 14'b1110011011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100010111;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110010;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101011001;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101011001;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100111;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110110100;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101000;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101001;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000010;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000011101;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101001;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101001;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110111;
SIGNAL_B = 14'b1110011000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000100;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011100000;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011111;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011111;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011111;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100010100;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100010100;
SIGNAL_B = 14'b1110010111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100010;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101010110;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101111100;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110010110;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101110000;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110010111;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b1110010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011001;
SIGNAL_B = 14'b1110010101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b1110010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111111111;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001011010;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001110;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001101;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b1110010100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010110110;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010110101;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100010010;
SIGNAL_B = 14'b1110010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101111010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000110;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111001000;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110111011;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111010101;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111100010;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000001001;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110000;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000100011;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110001;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001010111;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100101;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001101;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001110;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100101000;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100101000;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100101000;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101000010;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110111;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110110111;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010000;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101011;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111010;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000101101;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001001000;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001000111;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100010;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100110;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000000;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110011011;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110011011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b1110010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000010;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000110111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101010;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101010;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001011110;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001011110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010100000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100001;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100110000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100110000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001010;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100110000;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111101;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100100;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011000;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110010;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101001;
SIGNAL_B = 14'b1110001110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110110;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011011110;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010011;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111010;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110000111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b1110001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111101111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000001010;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010000000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110101;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010001100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b1110001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110111;
SIGNAL_B = 14'b1110001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100011100;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101101010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101101011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111000;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110010010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011111;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100010;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001110000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100100;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b1110001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101001101;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101001;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011101;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000011;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000100;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011001000;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101001010;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101010111;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100111101;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110100101;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111110100;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001011100;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010000;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101010;
SIGNAL_B = 14'b1110010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000100;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000110;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100100000;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101000111;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110101111;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010101;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111101;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110101111;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111101;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001010;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000010111;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110100;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100110;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011001;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010000000;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110100;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011011;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100000010;
SIGNAL_B = 14'b1110010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110110;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110101;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100001111;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100011101;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011110;
SIGNAL_B = 14'b1110010011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010100;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000000111;
SIGNAL_B = 14'b1110010100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111011;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b1110010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000101110;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010011000;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100100;
SIGNAL_B = 14'b1110010101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100100111;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000010;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b1110010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b1110010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b1110010111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b1110011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001010011;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111010;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100001;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001000;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111100;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111100;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b1110011010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b1110011001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b1110011010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110011;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b1110011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000001;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b1110011100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111110101;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b1110011100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000001;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000101001;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001110;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001011101;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001011101;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b1110011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100000110;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b1110011111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b1110011111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111011000;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111100100;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110001;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b1110100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000111111;
SIGNAL_B = 14'b1110100000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001001101;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000111111;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011011;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011100;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110110;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011010000;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110111;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b1110100100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b1110100101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b1110100111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b1110101000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110000;
SIGNAL_B = 14'b1110101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b1110101001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b1110101001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000000;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000000;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000000;
SIGNAL_B = 14'b1110101001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001110;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b1110101011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101011;
SIGNAL_B = 14'b1110101101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011111;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010001;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b1110101101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000101;
SIGNAL_B = 14'b1110101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000101;
SIGNAL_B = 14'b1110101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000110;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110110000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010110;
SIGNAL_B = 14'b1110110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010110;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110000;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001011;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001011;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111110;
SIGNAL_B = 14'b1110110100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b1110110011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b1110110101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011011;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011100;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b1110110110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101001;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010000;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b1110111001110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b1110111010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010100000;
SIGNAL_B = 14'b1110111010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010100000;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010100;
SIGNAL_B = 14'b1110111011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111011;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111011;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b1110111101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b1110111101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001000;
SIGNAL_B = 14'b1110111110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b1110111110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1110111111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b1111000001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b1111000001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011001;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b1111000011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111000110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111000110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111000111000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111001000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111001001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101010;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011110;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101011;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b1111010100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010010;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111010111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111010111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b1111011000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111011000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b1111011100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111011110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011101111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b1111100001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111100101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111100110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111100111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111101001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110100;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111101100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110011001101;
SIGNAL_B = 14'b1111110010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111110011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001011;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111110111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b0000000010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b0000000011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000000110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b0000000110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111101;
SIGNAL_B = 14'b0000001010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b0000001010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000001111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101011111;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101011;
SIGNAL_B = 14'b0000010010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000010101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110111;
SIGNAL_B = 14'b0000011000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101010;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011010;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b0000011111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000000;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b0000100001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000100000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000100010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001100;
SIGNAL_B = 14'b0000100011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001100;
SIGNAL_B = 14'b0000100100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b0000100100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100101;
SIGNAL_B = 14'b0000100100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000101000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b0000101000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b0000101011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100000111;
SIGNAL_B = 14'b0000101011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101101;
SIGNAL_B = 14'b0000101101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010000;
SIGNAL_B = 14'b0000101110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000011;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011101;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b0000101110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000110000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010000;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101001;
SIGNAL_B = 14'b0000110000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000001111;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001111;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b0000110010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001111;
SIGNAL_B = 14'b0000110011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b0000110011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b0000110011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110101000;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b0000110100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011000;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000110101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b0000110111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111110;
SIGNAL_B = 14'b0000110111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b0000110110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111110;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000111000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010110000;
SIGNAL_B = 14'b0000111000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010110000;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010110;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100010;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000110;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b0000111101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000110;
SIGNAL_B = 14'b0000111101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b0000111101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101011;
SIGNAL_B = 14'b0000111110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110111000;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010001;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b0000111111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0001000000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b0001000000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100001110;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110101;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011010;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011010;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b0001000001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110011;
SIGNAL_B = 14'b0001000010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110011;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b0001000011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b0001000101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b0001000101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000010110;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b0001000110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101101;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010100;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b0001001000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111011;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001001000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000111;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100111000;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b0001001001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000011;
SIGNAL_B = 14'b0001001010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110110;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010000;
SIGNAL_B = 14'b0001001011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000011;
SIGNAL_B = 14'b0001001011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b0001001100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011011;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b0001001011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100101;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100110;
SIGNAL_B = 14'b0001001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b0001001110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b0001001111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111100101;
SIGNAL_B = 14'b0001001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110111101;
SIGNAL_B = 14'b0001010000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111100;
SIGNAL_B = 14'b0001010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101101;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100111010;
SIGNAL_B = 14'b0001010000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010011;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b0001010010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101101;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b0001010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011110;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110110;
SIGNAL_B = 14'b0001010100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b0001010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000101001;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b0001010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111101000;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111001101;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111101000;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110011;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011010;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b0001010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001100;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b0001010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110011;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b0001010110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100011;
SIGNAL_B = 14'b0001010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b0001010111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010111;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010101;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100010;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010111;
SIGNAL_B = 14'b0001011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001000;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100011;
SIGNAL_B = 14'b0001011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111100;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010000111;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010010101;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111010;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001010011;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001000110;
SIGNAL_B = 14'b0001011011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000101100;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000010010;
SIGNAL_B = 14'b0001011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000010010;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111110111;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110111;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110010000;
SIGNAL_B = 14'b0001011101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000010;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101000;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110011100;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101001;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100100;
SIGNAL_B = 14'b0001011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001100011;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001100011;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b0001011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101101;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110011111;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101100;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111000;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011111;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101000100;
SIGNAL_B = 14'b0001100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010001;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011100;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100011101;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110110;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011001110;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011001110;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010101000;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010000001;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010000000;
SIGNAL_B = 14'b0001100011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000011000;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011010;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001011;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111100101;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111010111;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010110;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b0001100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001010;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010101;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001001;
SIGNAL_B = 14'b0001100101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100100000;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101100001;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100101101;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011111;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100101101;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010110111;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010111000;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010000;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101010;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101011;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101010;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b0001100111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000101000;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b0001100111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000001;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001101;
SIGNAL_B = 14'b0001101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110100101;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111000000;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101111111;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001101;
SIGNAL_B = 14'b0001101000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110110010;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100111101;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111011;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010101;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111011;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001111001;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010100000;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000011;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000100;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000011;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110110110;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101100111;
SIGNAL_B = 14'b0001101011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110101;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101001110;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011100101;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011010111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011100100;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001001;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001110000;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b0001101101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011110;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110010001;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100011100;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100011100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110101;
SIGNAL_B = 14'b0001101110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011101000;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100101;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110010;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110010;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000110001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000001010;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111111101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111110000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110000111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010011;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010011;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101100;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100100000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011011110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110110;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110101;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b0001110000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110100;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110010;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111101;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b0001110010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000111;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111000;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011101;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000010;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001110;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011101;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001110;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101110011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111101;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001100010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000100000;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111000100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111010010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101101010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101101010;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101000010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100000001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001001010;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110000;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101101;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010011;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011110111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111111111;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101100011;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101111101;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100001;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100001000;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001110111;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000100;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001111000;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001000100;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001000011;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001000100;
SIGNAL_B = 14'b0001101011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000011100;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110001100;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b0001101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110001;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100010111;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100011;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011110000;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010100010;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001101110;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b0001101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b0001101001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000011111;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111101011;
SIGNAL_B = 14'b0001100111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011111;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111000100;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001101;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b0001100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100100111;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b0001100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001110;
SIGNAL_B = 14'b0001100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111110;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111101;
SIGNAL_B = 14'b0001100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111100;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101101;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010101;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110101101;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000101;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101010010;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100010000;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100010001;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011101001;
SIGNAL_B = 14'b0001100011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011101;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110011;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001110;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001001100;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100110;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110001;
SIGNAL_B = 14'b0001100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110010;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101111100;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b0001011111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111011;
SIGNAL_B = 14'b0001011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101101;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b0001011110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b0001011111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b0001011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000100;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001011101;
SIGNAL_B = 14'b0001011101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011011;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011100;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110111111;
SIGNAL_B = 14'b0001011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000000;
SIGNAL_B = 14'b0001011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001010;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101011000;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b0001011001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001010;
SIGNAL_B = 14'b0001011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010101;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101100;
SIGNAL_B = 14'b0001011000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b0001010110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011111;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010000;
SIGNAL_B = 14'b0001010101111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011110;
SIGNAL_B = 14'b0001010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010000;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110101;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001101;
SIGNAL_B = 14'b0001010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101000001;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011001;
SIGNAL_B = 14'b0001010011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b0001010011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111111;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110010;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b0001010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100010;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100001;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b0001001111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010011;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010100;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010011;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010100;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110110;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101001;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b0001001000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b0001000111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b0001000111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011000;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b0001000110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b0001000110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b0001000111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b0001000100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b0001000100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b0001000100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b0001000011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100100;
SIGNAL_B = 14'b0001000011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b0001000010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b0001000010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b0001000000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100011111;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100000;
SIGNAL_B = 14'b0001000000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101110;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0000111111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111001;
SIGNAL_B = 14'b0000111110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0000111110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b0000111110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0000111110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b0000111101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b0000111001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110100;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b0000110111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b0000110111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011010;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b0000110110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b0000110110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b0000110110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110011;
SIGNAL_B = 14'b0000110101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100111;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100110;
SIGNAL_B = 14'b0000110100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b0000110011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b0000110010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b0000110001110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010110;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000110000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000110000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000101111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000101111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000101101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000101101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100010;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b0000101011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000101011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000101001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100001;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111010;
SIGNAL_B = 14'b0000100111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b0000100100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b0000100100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101101;
SIGNAL_B = 14'b0000100100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000110111;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b0000011111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b0000011101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000110111;
SIGNAL_B = 14'b0000011101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b0000011001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000011001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000011000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000011000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000011001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011100;
SIGNAL_B = 14'b0000010010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110001110;
SIGNAL_B = 14'b0000010001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000001111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110001110;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110000001;
SIGNAL_B = 14'b0000001011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110001111;
SIGNAL_B = 14'b0000000111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110000001;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110001111;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000000011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110001110;
SIGNAL_B = 14'b0000000010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b0000000000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000000010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b1111111111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b1111111111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b1111111111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b1111111001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111111000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111110111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111110111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101101;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111110010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100001;
SIGNAL_B = 14'b1111101111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101110;
SIGNAL_B = 14'b1111110000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111101110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b1111101111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b1111101110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111011;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b1111101101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100010;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100101111;
SIGNAL_B = 14'b1111101010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100101111;
SIGNAL_B = 14'b1111101010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111101010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001000;
SIGNAL_B = 14'b1111101001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111101000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100010;
SIGNAL_B = 14'b1111100111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111000000;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111100001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111100000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b1111011111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011010;
SIGNAL_B = 14'b1111011110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b1111011100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b1111011001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b1111011000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111011000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111010111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111010111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101011;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101100;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101100;
SIGNAL_B = 14'b1111010100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101100;
SIGNAL_B = 14'b1111010100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100000;
SIGNAL_B = 14'b1111010100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000110;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100010;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110110000;
SIGNAL_B = 14'b1111001111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010111;
SIGNAL_B = 14'b1111001111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001010;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111001110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b1111001110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100100;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b1111001101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b1111001100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100101;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001111;
SIGNAL_B = 14'b1111001010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b1111001011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110101;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011100;
SIGNAL_B = 14'b1111001010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101001;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011100;
SIGNAL_B = 14'b1111000111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b1111000101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110110;
SIGNAL_B = 14'b1111000110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b1111000100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b1111000011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010011;
SIGNAL_B = 14'b1111000010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b1111000010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000000111;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b1111000010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100001;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000000111;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010001010;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111111;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110010;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001100;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100000000;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b1110111100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110011;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101011011;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110101;
SIGNAL_B = 14'b1110111011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b1110111010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b1110111001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000101;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000101;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101100;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b1110110110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b1110110110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010110;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010111;
SIGNAL_B = 14'b1110110011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001001;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111110;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b1110110010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111110;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110011001;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110011001;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b1110110001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000001;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b1110110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000000;
SIGNAL_B = 14'b1110110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000001;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110101;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b1110101111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001011101;
SIGNAL_B = 14'b1110101110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110111;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000100;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101010;
SIGNAL_B = 14'b1110101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010010;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111001;
SIGNAL_B = 14'b1110101100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111011;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100001;
SIGNAL_B = 14'b1110101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110001001;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b1110101010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110001001;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110010;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110010;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011000;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b1110101000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010101000;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001110;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010101000;
SIGNAL_B = 14'b1110100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011101001;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011101001;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011110110;
SIGNAL_B = 14'b1110100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b1110100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000101;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000101;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101010010;
SIGNAL_B = 14'b1110100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011110;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111001;
SIGNAL_B = 14'b1110100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b1110100011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111011;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100010;
SIGNAL_B = 14'b1110100011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b1110100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010110;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000101111;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001001010;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010110;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011001;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011001;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001101;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101000010;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101000010;
SIGNAL_B = 14'b1110011111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b1110011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b1110011110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110011101;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000011111;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010011;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001010100;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100000;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111011;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010000111;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010001000;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011110000;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011110000;
SIGNAL_B = 14'b1110011100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b1110011100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110001;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b1110011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000011101;
SIGNAL_B = 14'b1110011001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b1110011010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000011100;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110110;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001000011;
SIGNAL_B = 14'b1110011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001000011;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000011100;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001111000;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001111000;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011111;
SIGNAL_B = 14'b1110011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011111;
SIGNAL_B = 14'b1110011000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b1110011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011100000;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100111011;
SIGNAL_B = 14'b1110010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100001;
SIGNAL_B = 14'b1110010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101001000;
SIGNAL_B = 14'b1110010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101101111;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101110000;
SIGNAL_B = 14'b1110010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b1110010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101111100;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110100100;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110100011;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111111111;
SIGNAL_B = 14'b1110010101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b1110010110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b1110010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001101;
SIGNAL_B = 14'b1110010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010000010;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010110110;
SIGNAL_B = 14'b1110010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011011101;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011110111;
SIGNAL_B = 14'b1110010011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101111001;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111001000;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101110;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000001001;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110111011;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110111010;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111100010;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110000;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000111101;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110010;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000111101;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110010;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011000;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001110;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011110100;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101000011;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101001111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110110;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110000011;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110110;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110000100;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111000101;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000111;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000100000;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000100000;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000101101;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001001000;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001000111;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001111100;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100010;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100101;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101011001;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101011001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100110;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110011010;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110001110;
SIGNAL_B = 14'b1110001110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000001;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110100;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011101;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000110111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011101;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010100000;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010010011;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010010011;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011010100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100001;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011010100;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011010100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111101;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001001;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100100;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111101;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001011;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110100;
SIGNAL_B = 14'b1110001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110010101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111010110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110111100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111111101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000110001;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001111111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100000010;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101101010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b1110001101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111000101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000010100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001010101;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100011;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010010110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010010110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100011;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011100101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101001101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000010;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000010;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110110110;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110110110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000100;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000111000;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000111000;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000110;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010100000;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011101111;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101100100;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101011000;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111000000;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001000010;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001011100;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001110110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101011;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010011110;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000101;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000110;
SIGNAL_B = 14'b1110010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000101;
SIGNAL_B = 14'b1110010001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100011;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111101;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010101;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111100;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001011;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110010;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011010;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011001;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011001;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010000000;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010000000;
SIGNAL_B = 14'b1110010010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b1110010010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100011110;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101000100;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011110;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101100;
SIGNAL_B = 14'b1110010011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000101;
SIGNAL_B = 14'b1110010100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110011111;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111000111;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000001000;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000001000;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b1110010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001100011;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100100;
SIGNAL_B = 14'b1110010101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b1110010110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110010;
SIGNAL_B = 14'b1110010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b1110010101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b1110010111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101001;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110011100;
SIGNAL_B = 14'b1110011000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110011100;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000101;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000101101;
SIGNAL_B = 14'b1110011000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000100;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011111;
SIGNAL_B = 14'b1110011000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010000111;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100001;
SIGNAL_B = 14'b1110011000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010101;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010111;
SIGNAL_B = 14'b1110011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110010;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101111111;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b1110011010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111110100;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b1110011101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011011111;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100000111;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111101;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110111110;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110010111;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100100;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111100100;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111111;
SIGNAL_B = 14'b1110100000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b1110100000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b1110100001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001001101;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b1110100001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b1110100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011010000;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110101;
SIGNAL_B = 14'b1110100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010000;
SIGNAL_B = 14'b1110100011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011101;
SIGNAL_B = 14'b1110100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010011;
SIGNAL_B = 14'b1110100101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111011;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000010101;
SIGNAL_B = 14'b1110100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b1110100111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b1110101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011001;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b1110101001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001100;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000000;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b1110101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b1110101010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b1110101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b1110101011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b1110101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b1110101100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b1110101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010001;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111000;
SIGNAL_B = 14'b1110101100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101100;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b1110101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b1110101110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111010;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b1110101110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b1110101111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100011;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110110000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111101;
SIGNAL_B = 14'b1110110001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111101;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111110;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001010;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001011;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100010111;
SIGNAL_B = 14'b1110110010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b1110110010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001011;
SIGNAL_B = 14'b1110110010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b1110110101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b1110110101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b1110110110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b1110110110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001111;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101001;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b1110111001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b1110111001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000011;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b1110111001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b1110111011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010100000;
SIGNAL_B = 14'b1110111011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000111;
SIGNAL_B = 14'b1110111011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b1110111101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100001;
SIGNAL_B = 14'b1110111101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b1110111110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1110111111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b1111000000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111101;
SIGNAL_B = 14'b1111000010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b1111000011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b1111000010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b1111000011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b1111000011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b1111000100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111001000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000100;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110111;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011111000;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b1111001111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b1111010010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010010;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101110;
SIGNAL_B = 14'b1111010101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010110110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b1111011000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111011000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b1111011001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b1111011011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111101;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111100001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b1111100001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b1111100011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111100101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100110;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111101000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111101011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111101010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101101111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111101101111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111110000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011010;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111110000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110100;
SIGNAL_B = 14'b1111110001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011010;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110011;
SIGNAL_B = 14'b1111110011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111110101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111111010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b1111111111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b0000000001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b0000000100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000000101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111101;
SIGNAL_B = 14'b0000000110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111100;
SIGNAL_B = 14'b0000001000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000001001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000001110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000010000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000001111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101011111;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b0000010001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b0000010011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b0000010100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000101;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011110;
SIGNAL_B = 14'b0000010111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101011;
SIGNAL_B = 14'b0000010111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001100111;
SIGNAL_B = 14'b0000011110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000000;
SIGNAL_B = 14'b0000011111000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000011111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001100;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111111;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b0000100100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001100;
SIGNAL_B = 14'b0000100100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100101;
SIGNAL_B = 14'b0000100100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100101;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010101;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b0000101000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b0000101000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100001;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b0000101001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b0000101010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100000111;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b0000101100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b0000101011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010010;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000101;
SIGNAL_B = 14'b0000101101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b0000101110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b0000101110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111010;
SIGNAL_B = 14'b0000101111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010000;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b0000110001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b0000110010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110101;
SIGNAL_B = 14'b0000110101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110101;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b0000110110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110001;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001011;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111101;
SIGNAL_B = 14'b0000110111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000110111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111110;
SIGNAL_B = 14'b0000111000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000111000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010111;
SIGNAL_B = 14'b0000111000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b0000111001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001010;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100011;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b0000111011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b0000111011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000110;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000110;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010010;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010001;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010010;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b0000111111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b0000111111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b0001000000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b0001000000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011011;
SIGNAL_B = 14'b0001000000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110110;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011011;
SIGNAL_B = 14'b0001000001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100001101;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000000;
SIGNAL_B = 14'b0001000010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011011;
SIGNAL_B = 14'b0001000001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001100;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001001;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000010110;
SIGNAL_B = 14'b0001000101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b0001000110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b0001000111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b0001001000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100111000;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011101;
SIGNAL_B = 14'b0001001011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b0001001010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101001;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110111;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b0001001100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b0001001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b0001001101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100110;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000111111;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110011;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011000;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110011;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111111;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111110;
SIGNAL_B = 14'b0001001111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111011000;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001010;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110010110;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b0001010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111100;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b0001010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100111011;
SIGNAL_B = 14'b0001010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b0001010000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b0001010010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011110;
SIGNAL_B = 14'b0001010010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010010;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000110;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011111;
SIGNAL_B = 14'b0001010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001111000;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110101;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001110;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111101000;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111100111;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b0001010101111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101111111;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101111111;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b0001011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010110;
SIGNAL_B = 14'b0001011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001000;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010101110;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100011;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100011;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100010;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010000111;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b0001011011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000101;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110011100;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101000;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101001;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101001;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100100110;
SIGNAL_B = 14'b0001011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100001100;
SIGNAL_B = 14'b0001011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100101;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110001;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110010;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111110;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110001;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000111100;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100001;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111010;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111011;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111010;
SIGNAL_B = 14'b0001100001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111000110;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101101;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110011111;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000101;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000101;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011111;
SIGNAL_B = 14'b0001100001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010001;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100011100;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100000011;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011100;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100001111;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110100;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110100;
SIGNAL_B = 14'b0001100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100111;
SIGNAL_B = 14'b0001100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000111111;
SIGNAL_B = 14'b0001100011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000011000;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b0001100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111110;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001001;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111010111;
SIGNAL_B = 14'b0001100101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001001;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001010;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001010;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101111;
SIGNAL_B = 14'b0001100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010101;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100100000;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101000111;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101110;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010011;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011101100;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010111000;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010011101;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101010;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010000;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010000;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001000010;
SIGNAL_B = 14'b0001100111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000101000;
SIGNAL_B = 14'b0001100111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001101;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000001;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b0001101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001101;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110110011;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110100101;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101111111;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101100101;
SIGNAL_B = 14'b0001101001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011100010;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111011;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011001000;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010100;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011101;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011101;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111010000;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000010;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101100111;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100100110;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011111110;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100100110;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011011000;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010111110;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001001000;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001010;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001001000;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101101;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010011;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111000110;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101101010;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101001;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100000010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100000010;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100000010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100011100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010001100;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010001100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010000000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100101;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000001010;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000001010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010100;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111010;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011100;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011011;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011011;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011011;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100101;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100101;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100110000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010100000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010010011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101011;
SIGNAL_B = 14'b0001110000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011101;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110100;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101011001;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111101;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001100001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101101010;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110111;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010111111;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110010;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000111110;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101101;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000110;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101111010;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000101;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010001111;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110100;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001011011;
SIGNAL_B = 14'b0001101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001110;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110111110;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101001001;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101010110;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100111011;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100010100;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011111;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010010001;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001111000;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101001;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101010;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000010;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110001101;
SIGNAL_B = 14'b0001101011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b0001101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110001;
SIGNAL_B = 14'b0001101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101011001;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011110000;
SIGNAL_B = 14'b0001101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001010;
SIGNAL_B = 14'b0001101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010001000;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001101110;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001010100;
SIGNAL_B = 14'b0001101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000011111;
SIGNAL_B = 14'b0001101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111111001;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b0001101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011011;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100100111;
SIGNAL_B = 14'b0001100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001110001;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111110;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001001010;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100010;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111100;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111011;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110101101;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011110110;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000100;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000100;
SIGNAL_B = 14'b0001100011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011101001;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b0001100011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011001111;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100110;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110001;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101111100;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111010;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b0001011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111001;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101101;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110111;
SIGNAL_B = 14'b0001011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101010;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b0001011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110110;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111100111;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000000;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111101;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001001;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b0001011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b0001010111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101100;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101100;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010010;
SIGNAL_B = 14'b0001010101111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101010;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110101;
SIGNAL_B = 14'b0001010011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101100111;
SIGNAL_B = 14'b0001010100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101000001;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100111;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100111;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011001;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011001;
SIGNAL_B = 14'b0001010011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001100;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b0001010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110010;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b0001010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b0001010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100001;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000000111;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010100;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000111;
SIGNAL_B = 14'b0001001101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111010;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101010;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010000;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b0001001011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b0001001011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b0001001010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b0001000111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b0001001000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010101000;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001011;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111110;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111110;
SIGNAL_B = 14'b0001000110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000010111;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001010;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b0001000011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b0001000011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b0001000100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010111;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110110000;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100000;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b0001000001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100011111;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010011;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b0000111111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0000111111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0000111110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011111;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b0000111110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b0000111101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b0000111100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011011;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011011;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000111010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000111000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000100111;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110100;
SIGNAL_B = 14'b0000111000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b0000111000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b0000110110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001010;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b0000110011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b0000110000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100101111;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000101111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b0000101101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000101010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000100111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000100111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000100110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b0000100101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000111;
SIGNAL_B = 14'b0000100011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000101;
SIGNAL_B = 14'b0000100011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b0000100011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000100010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b0000100000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000011110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000011011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000011010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000010111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000010110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000010101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000010001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000001110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000001101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000001100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000001100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110001110;
SIGNAL_B = 14'b0000001010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000001010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000000110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000000100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000000001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b1111111111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b1111111110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b1111111011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b1111111001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b1111111000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b1111110111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b1111110111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111111000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b1111110101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111110000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111101111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101110;
SIGNAL_B = 14'b1111110000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b1111101110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111101110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001000;
SIGNAL_B = 14'b1111101110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101110;
SIGNAL_B = 14'b1111101101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b1111101101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b1111101101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010101;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111101010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110001;
SIGNAL_B = 14'b1111101010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b1111101010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111110;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111100;
SIGNAL_B = 14'b1111101000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010110;
SIGNAL_B = 14'b1111101000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111100110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010110;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111100110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001001;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011001;
SIGNAL_B = 14'b1111100011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b1111011110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011010;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011011;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011110;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111011000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000101;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111010110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011111;
SIGNAL_B = 14'b1111010111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010010;
SIGNAL_B = 14'b1111010100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101100;
SIGNAL_B = 14'b1111010100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111001;
SIGNAL_B = 14'b1111010001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b1111010011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110110000;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100010;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111101;
SIGNAL_B = 14'b1111001111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111001110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100100;
SIGNAL_B = 14'b1111001110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000010111;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100111;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b1111001010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b1111001010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b1111001001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b1111001001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b1111001000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b1111001000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b1111000111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b1111000111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100001111;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b1111000110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000011;
SIGNAL_B = 14'b1111000110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010011;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010011;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111010;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b1111000000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b1111000000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b1111000000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b1111000000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100010;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100010;
SIGNAL_B = 14'b1110111111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110001;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110001;
SIGNAL_B = 14'b1110111110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b1110111110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b1110111101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100110;
SIGNAL_B = 14'b1110111101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b1110111100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011001;
SIGNAL_B = 14'b1110111100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101000001;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110100;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111111000;
SIGNAL_B = 14'b1110111010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101010;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110111;
SIGNAL_B = 14'b1110111000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011110;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b1110111000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011111;
SIGNAL_B = 14'b1110110110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010010;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b1110110111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001011111;
SIGNAL_B = 14'b1110110111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b1110110110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b1110110101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b1110110100011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001001;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101011000;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111101;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110001;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001101;
SIGNAL_B = 14'b1110110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001101;
SIGNAL_B = 14'b1110110001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111100111;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101000;
SIGNAL_B = 14'b1110110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000001;
SIGNAL_B = 14'b1110101111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110111;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000011;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101010;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b1110101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b1110101101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011100000;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100000;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b1110101100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101111100;
SIGNAL_B = 14'b1110101100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b1110101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101111011;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101111100;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110001001;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111100100;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111100101;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011001;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110010;
SIGNAL_B = 14'b1110101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011000;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001001101;
SIGNAL_B = 14'b1110101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b1110100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001110;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010000001;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010011011;
SIGNAL_B = 14'b1110100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011110110;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b1110100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b1110100110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100101010;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101011;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000110;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000110;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111000111;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111011;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b1110100011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111011;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000101111;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000101111;
SIGNAL_B = 14'b1110100010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010110;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001100100;
SIGNAL_B = 14'b1110100010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001110001;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111101;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110100000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100100111;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011011;
SIGNAL_B = 14'b1110100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001110;
SIGNAL_B = 14'b1110011111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110010000;
SIGNAL_B = 14'b1110011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111101100;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b1110011101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000011111;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010010;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000110;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b1110011100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010100;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111011;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010100010;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010101111;
SIGNAL_B = 14'b1110011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010101111;
SIGNAL_B = 14'b1110011100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001010;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001011;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001010;
SIGNAL_B = 14'b1110011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b1110011011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110001101;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110110100;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111110101;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110110;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000010000;
SIGNAL_B = 14'b1110011001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011110;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000001111;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110110;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010010010;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101010;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010010010;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011110;
SIGNAL_B = 14'b1110011000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011010011;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101110;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100010100;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101110;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101100011;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101010110;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101110000;
SIGNAL_B = 14'b1110010110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100111011;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110010110;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b1110010110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011010;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001011010;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010001111;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011000;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b1110010101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010000010;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b1110010101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011011101;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101000101;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110100001;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101110;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111100010;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110111011;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111001000;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000111110;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001011000;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000100011;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110010;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111110;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101000010;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001111;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101000010;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110111;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011100;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011100;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011101;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101011;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011101;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111010001;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000010011;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000101110;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000101101;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000011111;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111011;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100011;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111100;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111101;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100101;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100111111;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000001;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110011011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110011010;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011011;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101011;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101011;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010100000;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111000;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010010011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111001;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110000;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110010111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100101;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000101000;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110101;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110110;
SIGNAL_B = 14'b1110001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011011110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111010;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110111100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b1110001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010001100;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011001110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011001110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011001110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000011;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110101;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000100;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101101010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000101;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010011;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000010100;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100011;
SIGNAL_B = 14'b1110001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010111110;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010111110;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100100110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101001101;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110110101;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111110111;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000111000;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011001000;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010100;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100111101;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001101;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101111110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101111110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111110100;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010000;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000110101;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000101;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010001;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011111;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011101100;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011111001;
SIGNAL_B = 14'b1110010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010011;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111100;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110101111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110101111;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111010111;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111010111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001011;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100110;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011010;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000001;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101001;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100011100;
SIGNAL_B = 14'b1110010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101000;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100011101;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101000100;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111001;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111000111;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101100;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100000;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000001000;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101110;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111011;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001100011;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110001;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100100;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100001100;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b1110010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101110101;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000010;
SIGNAL_B = 14'b1110010110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101110100;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000010010;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000100;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011111;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011111;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001000110;
SIGNAL_B = 14'b1110011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010000111;
SIGNAL_B = 14'b1110011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010010101;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100010;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100010;
SIGNAL_B = 14'b1110011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001000;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b1110011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100011;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100100;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100001010;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010111;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011010;
SIGNAL_B = 14'b1110011001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101111111;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111001101;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110011;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111101000;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111110100;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000100;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001111000;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010010;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111001;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111001;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100111010;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b1110011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b1110011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110001;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110010110;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110010111;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001010;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001010;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111111;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111100100;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b1110100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100110;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100110;
SIGNAL_B = 14'b1110100000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001001101;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011011;
SIGNAL_B = 14'b1110100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011011;
SIGNAL_B = 14'b1110100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110101;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b1110100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011101;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011100;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011100;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b1110100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b1110100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110110;
SIGNAL_B = 14'b1110100100011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b1110100011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101101;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b1110100110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000010101;
SIGNAL_B = 14'b1110100111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001001;
SIGNAL_B = 14'b1110100110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b1110100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100010;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000101111;
SIGNAL_B = 14'b1110100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b1110101000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b1110100111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b1110101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011010;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b1110101010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001100;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100001110;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011010;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100101000;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b1110101011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011110;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110111000;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000110;
SIGNAL_B = 14'b1110101101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010010;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b1110101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000110;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100011;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b1110110001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b1110110001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110001;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110000;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b1110110011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110101;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110101;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b1110110110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110110;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b1110111010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011101;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b1110111011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b1110111011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b1110111011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101110;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111011;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b1110111100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b1110111110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001000;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010100;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111101;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1110111110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100010;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100010;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001011;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b1111000001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100101;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100101;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b1111000010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011001;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b1111000100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000000000;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b1111000100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111001000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001100111;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111001000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110111;
SIGNAL_B = 14'b1111001010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b1111001011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101011;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011111000;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011111000;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011111000;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010001;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010001;
SIGNAL_B = 14'b1111001110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111001111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b1111010000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000101;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111010111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111010111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b1111011001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b1111011001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b1111011010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111011011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111011111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b1111100000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b1111100001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111100110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111100110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111110001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b0000000010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b0000000100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b0000000101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000001000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b0000000111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b0000000111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000001010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b0000001100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b0000001111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000001111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111100;
SIGNAL_B = 14'b0000010000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000010000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000010001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010001;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011110;
SIGNAL_B = 14'b0000010111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000011001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011110;
SIGNAL_B = 14'b0000011000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000100;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110111;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011101;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001100111;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011111000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b0000011111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000100000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000100000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000100001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000100001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001100;
SIGNAL_B = 14'b0000100001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100110;
SIGNAL_B = 14'b0000100011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100110;
SIGNAL_B = 14'b0000100010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110010;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001100;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b0000100100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b0000100111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010101;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001000;
SIGNAL_B = 14'b0000100111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b0000101010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100001;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010100;
SIGNAL_B = 14'b0000101001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101110;
SIGNAL_B = 14'b0000101011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010100;
SIGNAL_B = 14'b0000101011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010100000;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b0000101111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110110;
SIGNAL_B = 14'b0000101111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011101;
SIGNAL_B = 14'b0000101111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b0000101111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101001;
SIGNAL_B = 14'b0000110011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b0000110011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001011;
SIGNAL_B = 14'b0000110101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110001;
SIGNAL_B = 14'b0000110110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001011;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b0000110110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b0000111000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000111000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b0000111001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000111001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100011;
SIGNAL_B = 14'b0000111010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010110;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b0000111011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b0000111011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111001;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111010;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111010;
SIGNAL_B = 14'b0000111101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010010;
SIGNAL_B = 14'b0000111101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011111;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000101;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b0000111111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b0000111111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b0001000000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110101;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100001101;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001100;
SIGNAL_B = 14'b0001000010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b0001000010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001101;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001100;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b0001000101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b0001000011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001000;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b0001000110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b0001000111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010101;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010101;
SIGNAL_B = 14'b0001000111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010011;
SIGNAL_B = 14'b0001000111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b0001000111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b0001001001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011101;
SIGNAL_B = 14'b0001001010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b0001001010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b0001001011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b0001001011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b0001001100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001001101;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100110;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b0001001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110011;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001010;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001011;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001011;
SIGNAL_B = 14'b0001010000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b0001010001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b0001010000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001010;
SIGNAL_B = 14'b0001010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100111011;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100000;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101101;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b0001010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111010;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010011;
SIGNAL_B = 14'b0001010011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111001;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011101;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001011101;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110110;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000010;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000001;
SIGNAL_B = 14'b0001010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111100111;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111001101;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001100;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110100;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110011;
SIGNAL_B = 14'b0001010110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110011;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110011;
SIGNAL_B = 14'b0001011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b0001011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100011;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111100;
SIGNAL_B = 14'b0001010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010101111;
SIGNAL_B = 14'b0001011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100011;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001000;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010101110;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111010;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010000111;
SIGNAL_B = 14'b0001011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000100;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001010011;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000101;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111000011;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b0001011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000010;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000010;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101110101;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101000;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011111111;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b0001011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110010;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b0001011110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100100;
SIGNAL_B = 14'b0001011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b0001011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b0001011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000101111;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000000111;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111011;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b0001100001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101100;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111010;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000110;
SIGNAL_B = 14'b0001100001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000101;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000101;
SIGNAL_B = 14'b0001100010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b0001100011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010001;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b0001100011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101000100;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110101;
SIGNAL_B = 14'b0001100011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110110;
SIGNAL_B = 14'b0001100010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110100;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110100;
SIGNAL_B = 14'b0001100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011010;
SIGNAL_B = 14'b0001100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100110;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110001;
SIGNAL_B = 14'b0001100011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110000;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111101;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111100100;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111100011;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111101;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010101;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110101111;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101100001;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100101101;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010010;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010011;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011111001;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011101011;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000100;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011101100;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010110111;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b0001100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010011101;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000110101;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b0001100111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000110101;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011001;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110100101;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101010111;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101010111;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101001010;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011101110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111011;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b0001101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000110;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001011111;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001011111;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001011111;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000111000;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010001;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010001;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101001;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000011;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110110101;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101101000;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101100111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100100110;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011100101;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100100;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100100;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001010101;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000101111;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111000;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110010010;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000011;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101010000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100000010;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011101000;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011001101;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100101;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001111111;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100101;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100101;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001011;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000110001;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111010110;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111110000;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101110;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110001000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100100000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011011110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011011101;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011100;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000010;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011100;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011011;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001111;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110001;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100101;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110001;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001010;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110000;
SIGNAL_B = 14'b0001110001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110001;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101100;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111000;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001000100;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000100;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000010;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011110;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010001;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000110;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101010;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011101;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110110;
SIGNAL_B = 14'b0001101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011110100;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001101;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100100;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110010;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001010111;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000001001;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111101111;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110100001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101011111;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101000101;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100010001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100010001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011011101;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010000010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011011;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010001110;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010000010;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001101000;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111111111;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110111110;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110100100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101100010;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100010100;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011100000;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011010011;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011111;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011110;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110111;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000001111;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000010;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101111111;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110001;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100011000;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111101;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001010;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010110;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010001000;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010000111;
SIGNAL_B = 14'b0001101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001101101;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000110;
SIGNAL_B = 14'b0001101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101101;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111000100;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111000100;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110011101;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b0001100111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101000010;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001110;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001110;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100101000;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011010;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010011000;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001110001;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111101;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001100011;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101111;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100010;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b0001100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010100;
SIGNAL_B = 14'b0001100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000101;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101010001;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101010010;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011110110;
SIGNAL_B = 14'b0001100011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010101000;
SIGNAL_B = 14'b0001100010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010011011;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010000001;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b0001100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011000;
SIGNAL_B = 14'b0001100000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111100100;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111001010;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b0001100001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b0001011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111010;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010010;
SIGNAL_B = 14'b0001011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111001;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110111;
SIGNAL_B = 14'b0001011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011011111;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000100;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110111;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000010;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101010;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110101;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000001;
SIGNAL_B = 14'b0001011100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000001;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111100111;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111100111;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b0001011011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000000;
SIGNAL_B = 14'b0001011010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b0001011010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b0001011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111101;
SIGNAL_B = 14'b0001011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110000;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b0001010110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b0001010110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011111;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b0001010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b0001010101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b0001010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110101;
SIGNAL_B = 14'b0001010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101011010;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101100111;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100111;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b0001010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100000000;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110001;
SIGNAL_B = 14'b0001010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100110;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b0001010001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010001010;
SIGNAL_B = 14'b0001010000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b0001001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101110;
SIGNAL_B = 14'b0001001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101110;
SIGNAL_B = 14'b0001001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b0001001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000111;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b0001001010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b0001001010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101001;
SIGNAL_B = 14'b0001001001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b0001001010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110101;
SIGNAL_B = 14'b0001001000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010101000;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001111;
SIGNAL_B = 14'b0001001000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011000;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b0001000111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b0001000110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b0001000101111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000010111;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100100;
SIGNAL_B = 14'b0001000011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b0001000010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100010;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b0001000010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110000111;
SIGNAL_B = 14'b0001000011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010011;
SIGNAL_B = 14'b0001000000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b0000111110110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011111;
SIGNAL_B = 14'b0000111110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011110;
SIGNAL_B = 14'b0000111101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000111001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b0000110111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b0000111000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001101;
SIGNAL_B = 14'b0000111000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000111000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b0000110110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011010;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000000;
SIGNAL_B = 14'b0000110101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001101;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000110000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b0000101111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001001;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101110110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000101110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000101110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010110;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001001;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b0000101101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b0000101100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000101010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b0000101010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000100111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111000;
SIGNAL_B = 14'b0000100100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100001;
SIGNAL_B = 14'b0000100100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000110111;
SIGNAL_B = 14'b0000100011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111010;
SIGNAL_B = 14'b0000100001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b0000100000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000011111000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000110111;
SIGNAL_B = 14'b0000011100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000011100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000010101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000010101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000001011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011100;
SIGNAL_B = 14'b0000001011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000001010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000001000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000000001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000000000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b1111111101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b1111111100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111111010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000110111;
SIGNAL_B = 14'b1111111011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b1111111000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111110111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111110110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b1111110001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001000;
SIGNAL_B = 14'b1111101010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001000;
SIGNAL_B = 14'b1111101010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001001;
SIGNAL_B = 14'b1111101000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111101000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100101111;
SIGNAL_B = 14'b1111101000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111100110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111000000;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111100010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111100000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111000000;
SIGNAL_B = 14'b1111100000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110100;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000000;
SIGNAL_B = 14'b1111011110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100111;
SIGNAL_B = 14'b1111011110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b1111011110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b1111011101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011010;
SIGNAL_B = 14'b1111011101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b1111011101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111011001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010010;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010111000;
SIGNAL_B = 14'b1111011000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101011;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000101;
SIGNAL_B = 14'b1111010110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b1111010110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b1111010101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000101;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b1111010011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000110;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101100;
SIGNAL_B = 14'b1111010010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111001;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111001111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110001;
SIGNAL_B = 14'b1111001101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110001;
SIGNAL_B = 14'b1111001101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110001;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001011;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100100;
SIGNAL_B = 14'b1111001100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001011;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110101;
SIGNAL_B = 14'b1111001001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110101;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110101;
SIGNAL_B = 14'b1111001001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b1111001001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110110;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001111;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b1111001000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b1111000111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101001;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011100;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100001111;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b1111000101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b1111000100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000111;
SIGNAL_B = 14'b1111000011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1111000001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111010;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001000;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b1111000001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1110111111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b1111000000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100010;
SIGNAL_B = 14'b1110111111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b1110111111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110010;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b1110111110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100111;
SIGNAL_B = 14'b1110111101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110011;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011001;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101000001;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100110;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110101;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110100;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111000011;
SIGNAL_B = 14'b1110111001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101010;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111111000;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b1110111000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101100;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b1110110111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101011;
SIGNAL_B = 14'b1110110110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b1110110110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b1110110101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b1110110011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b1110110011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b1110110011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110011001;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000001;
SIGNAL_B = 14'b1110110000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011011;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011100;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011100;
SIGNAL_B = 14'b1110101111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b1110101110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101001;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110101;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b1110101101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000110;
SIGNAL_B = 14'b1110101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010011;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010010;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010011;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b1110101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000111;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100000;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b1110101100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011001;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110001;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b1110101010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b1110101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000111111;
SIGNAL_B = 14'b1110101001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b1110101000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001110;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010011011;
SIGNAL_B = 14'b1110100111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001101;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011001111;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000100;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100010001;
SIGNAL_B = 14'b1110100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011110;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000101;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111000;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111000111;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101111;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100010;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111100;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100011;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111101;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001001010;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b1110100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011100110;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b1110100000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011001;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110100;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100100111;
SIGNAL_B = 14'b1110011111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110100;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101000010;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001110;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b1110011111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110011101;
SIGNAL_B = 14'b1110011111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010010;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111101011;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111111000;
SIGNAL_B = 14'b1110011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100000;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111010;
SIGNAL_B = 14'b1110011100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010001000;
SIGNAL_B = 14'b1110011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010000111;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010100010;
SIGNAL_B = 14'b1110011100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010100010;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001010;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b1110011100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110010;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100111;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101000;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101000;
SIGNAL_B = 14'b1110011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101001;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000011100;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101000;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101001;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011101;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b1110011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011101;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011110;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010101011;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011010011;
SIGNAL_B = 14'b1110010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011100000;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b1110010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100001000;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101110;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100111011;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101010110;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101101111;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110111110;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110100011;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110100011;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b1110010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010000010;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001100111;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010101001;
SIGNAL_B = 14'b1110010100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011011;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000010;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b1110010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100010001;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100010010;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000101;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101000101;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000110;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110111010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110111011;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000001001;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001001011;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000100011;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000111101;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110000;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001001011;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001010111;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110110;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110000100;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101010;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000101101;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000100001;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001000111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000101110;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111101;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101011001;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101110100;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101110100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110100;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011101;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010001;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000110111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101010;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010001;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001011110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001011111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010100000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001001;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100100;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b1110001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110010;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011011;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100100000;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b1110001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010011;
SIGNAL_B = 14'b1110001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110000111;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110111100;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111010110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111110000;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100110;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011001101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000100;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111000110;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110010001;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101101;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011001011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011100101;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101000001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101001101;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101001;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000011;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011101;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001111010;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011001000;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010100;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010101;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101111110;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000001;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001000010;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001000010;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010011110;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010000;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010011101;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011110;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010010;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011111;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100101101;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101100001;
SIGNAL_B = 14'b1110010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101100001;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101100010;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111010110;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111101;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001011;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010000000;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110100;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110100;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110100;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011011;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101000100;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011110;
SIGNAL_B = 14'b1110010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000101;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111000;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110100000;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111011;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010100;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000001000;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000101111;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001100011;
SIGNAL_B = 14'b1110010101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b1110010101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110010;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b1110010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100100111;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b1110010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101000;
SIGNAL_B = 14'b1110010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011100;
SIGNAL_B = 14'b1110010111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110011101;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111000100;
SIGNAL_B = 14'b1110010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000101;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001010011;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b1110011000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001000;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111010;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010101;
SIGNAL_B = 14'b1110011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100100;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010111;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b1110011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110010;
SIGNAL_B = 14'b1110011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110011;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111110100;
SIGNAL_B = 14'b1110011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111110101;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b1110011100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110110;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001011101;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011110;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b1110011101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b1110011110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110000;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111100;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b1110100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110001;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110011;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b1110100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011011;
SIGNAL_B = 14'b1110100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011100;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b1110100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b1110100010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110110;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100111000;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010011;
SIGNAL_B = 14'b1110100101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100010;
SIGNAL_B = 14'b1110100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b1110100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b1110100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b1110101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100101000;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110101;
SIGNAL_B = 14'b1110101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011110;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110110111;
SIGNAL_B = 14'b1110101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011111;
SIGNAL_B = 14'b1110101100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010010;
SIGNAL_B = 14'b1110101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010001;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010010;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110101101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000011111;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b1110101111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010110;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b1110110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001011;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b1110110010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100010111;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001011;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b1110110100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001011;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001111;
SIGNAL_B = 14'b1110110110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b1110110110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001111;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000001111;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b1110110111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b1110111000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010000;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000011;
SIGNAL_B = 14'b1110111001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011101;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b1110111001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b1110111100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100000111;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b1110111100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b1110111101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100000111;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100010;
SIGNAL_B = 14'b1110111101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b1110111101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111011;
SIGNAL_B = 14'b1110111101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1110111101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1110111111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b1111000000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b1111000000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b1111000000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b1111000001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011001;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001100;
SIGNAL_B = 14'b1111000011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b1111000011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b1111000100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011001;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b1111000110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001101;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111001000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111001000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110011;
SIGNAL_B = 14'b1111001000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101010;
SIGNAL_B = 14'b1111001011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011110;
SIGNAL_B = 14'b1111001011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011110;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101011;
SIGNAL_B = 14'b1111001111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b1111010000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000101;
SIGNAL_B = 14'b1111010001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000101;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b1111010011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101011111;
SIGNAL_B = 14'b1111010101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111011000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111011001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010100;
SIGNAL_B = 14'b1111011000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b1111011010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111011101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111100000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111100000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111100001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111100111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111100111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111101000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111101000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111101011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111101100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111101110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110011000000;
SIGNAL_B = 14'b1111110010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111110111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111110111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111110111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b0000000010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000000111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000001010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b0000001101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000001110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000010000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b0000010011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b0000010100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b0000010110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011111000;
SIGNAL_B = 14'b0000010111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000011000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000010101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000010111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000010111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101010;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000011110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000100000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000100000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b0000100000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b0000100010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100110;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b0000100101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001000;
SIGNAL_B = 14'b0000101000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010100;
SIGNAL_B = 14'b0000101010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000101001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b0000101001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101101;
SIGNAL_B = 14'b0000101011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101101;
SIGNAL_B = 14'b0000101100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b0000101100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000101110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b0000101111000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010000;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b0000101111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110110;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000110001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b0000110010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000110011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001111;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001111;
SIGNAL_B = 14'b0000110100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b0000110100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b0000110101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b0000110101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001011;
SIGNAL_B = 14'b0000110101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000110110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b0000110111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110001;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000111000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001010;
SIGNAL_B = 14'b0000111001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b0000111001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b0000111001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b0000111001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b0000111011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b0000111010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b0000111100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b0000111011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111001;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b0000111101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111000;
SIGNAL_B = 14'b0000111100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101011;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110110111;
SIGNAL_B = 14'b0000111101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101011;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b0000111111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110110111;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b0001000000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100101000;
SIGNAL_B = 14'b0001000000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011011;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110101;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100001110;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b0001000010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011010;
SIGNAL_B = 14'b0001000010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b0001000010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b0001000011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b0001000011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b0001000100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b0001000101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b0001000110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000010110;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000101111;
SIGNAL_B = 14'b0001000110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b0001000110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100010;
SIGNAL_B = 14'b0001000111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101101;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b0001001000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100001;
SIGNAL_B = 14'b0001001000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010100;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b0001001001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100110111;
SIGNAL_B = 14'b0001001001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011100;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b0001001011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110110;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110101;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101001;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110011;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110001;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111111;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100110;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111011000;
SIGNAL_B = 14'b0001001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001010;
SIGNAL_B = 14'b0001001110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001011;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110111110;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b0001010000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b0001010000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b0001010010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b0001010010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010010;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011111;
SIGNAL_B = 14'b0001010011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010101011;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001110111;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001011101;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000101;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b0001010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001110;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000010;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001110;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111110101;
SIGNAL_B = 14'b0001010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111001101;
SIGNAL_B = 14'b0001010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110100;
SIGNAL_B = 14'b0001010101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001100;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b0001010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b0001010110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101111111;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001101;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011010;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b0001010111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100100;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b0001011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010101110;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001000;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111010;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001000110;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001000110;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000101011;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101010;
SIGNAL_B = 14'b0001011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000010001;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111000011;
SIGNAL_B = 14'b0001011100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101110101;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000010;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b0001011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b0001011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011001;
SIGNAL_B = 14'b0001011101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110001;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100101;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110001;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011011001;
SIGNAL_B = 14'b0001011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111110;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000111100;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101110;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101101;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101110;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111000110;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101100;
SIGNAL_B = 14'b0001100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110011111;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011110;
SIGNAL_B = 14'b0001100001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010001;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100011101;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b0001100010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100011101;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101000;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011100;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011010;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100111;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000010111;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110001;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111100011;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111010111;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001010;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010110;
SIGNAL_B = 14'b0001100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101100001;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101110;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100101101;
SIGNAL_B = 14'b0001100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101000111;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011111001;
SIGNAL_B = 14'b0001100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011110;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000110;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000101;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010001;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010010;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101011;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010110111;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001110110;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b0001100111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000110101;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000110101;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011001;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b0001100111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001100;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110110011;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001100;
SIGNAL_B = 14'b0001101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101100100;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101100101;
SIGNAL_B = 14'b0001101001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b0001101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001000;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111011;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111010;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010101;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001111010;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001111010;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011101;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101001;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000101;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111110111;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000011;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001111;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101000000;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101000000;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101000000;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010111110;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010010111;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010010110;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100010;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100010;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000010100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001001000;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000010100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010011;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111000;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110010001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101010000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101001;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101010000;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110100;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100000010;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100101;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011001;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000110001;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000110001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111111101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111010101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000110;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011011110;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010111000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101000;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011010;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110100;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110010111;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001011;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110000;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001010;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100001;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010100000;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010000110;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001011110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000110111;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110001110;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001100;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001100010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000101101;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000010100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111000101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101010;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101001111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110001;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001010111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000111101;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000001001;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110111011;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101000110;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011011101;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010001111;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110011;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111111111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110010111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101110000;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101100011;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100010100;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010010010;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011111;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011111;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011110;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011110;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110110;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101000;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111110101;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110001101;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101111111;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011011;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011001;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001011;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111110;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010101111;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b0001101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b0001101000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100000;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001010100;
SIGNAL_B = 14'b0001101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000011111;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b0001101000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b0001100111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101000010;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001110;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100100111;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110100;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011010;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011011;
SIGNAL_B = 14'b0001100110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111110;
SIGNAL_B = 14'b0001100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001110001;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001001010;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001001010;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000110000;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000101111;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010101;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100010;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111000111;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110101101;
SIGNAL_B = 14'b0001100101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000110;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111000;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100110111;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100010000;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011110110;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011110110;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011010000;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001110;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100110;
SIGNAL_B = 14'b0001100010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110010;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011000;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110010;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110001000;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b0001011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100000;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100000;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000111;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010011;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000100;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010011110;
SIGNAL_B = 14'b0001011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011100;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001001111;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011100;
SIGNAL_B = 14'b0001011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011011;
SIGNAL_B = 14'b0001011100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001110;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001101;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000000;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b0001011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111101;
SIGNAL_B = 14'b0001011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b0001011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b0001011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010110;
SIGNAL_B = 14'b0001011001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b0001011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b0001011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b0001010110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b0001010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111000011;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111000011;
SIGNAL_B = 14'b0001010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110111;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110101;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b0001010100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101000001;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b0001010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b0001010010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b0001010011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b0001010010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b0001010001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010001010;
SIGNAL_B = 14'b0001010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010101;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111011;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001000;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b0001001110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b0001001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010010;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b0001001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000011;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b0001001011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b0001001010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b0001001001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b0001001000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110001;
SIGNAL_B = 14'b0001000110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b0001000100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100010;
SIGNAL_B = 14'b0001000010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b0001000001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010011;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010010;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101100;
SIGNAL_B = 14'b0001000000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010010;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0000111111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011111;
SIGNAL_B = 14'b0000111110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011110;
SIGNAL_B = 14'b0000111011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001110;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101001;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b0000111000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000111000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011010;
SIGNAL_B = 14'b0000111001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b0000110111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001101;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001101;
SIGNAL_B = 14'b0000110111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111000000;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b0000110110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011010;
SIGNAL_B = 14'b0000110101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100110;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000110011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000101111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100010;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111100;
SIGNAL_B = 14'b0000101111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100010;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011001000;
SIGNAL_B = 14'b0000101100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111011;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011001000;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000101001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000101000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101110;
SIGNAL_B = 14'b0000100111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000100001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b0000100001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000011111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b0000011111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000100000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000011110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000011101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b0000011110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000011100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000011001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000011001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000010100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000001101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000001100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000001001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000000100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000000010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b1111111110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b1111111100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b1111111100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b1111111100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b1111111010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111111001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b1111111001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b1111110110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b1111110101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111110010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111110000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111101111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b1111101101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b1111101011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111101011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111101010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111101000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111101000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111101000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001001;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111100;
SIGNAL_B = 14'b1111100110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011001;
SIGNAL_B = 14'b1111100011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011001;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011001;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110011;
SIGNAL_B = 14'b1111100001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111100001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111100000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100110;
SIGNAL_B = 14'b1111100001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111100001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011010;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110100;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000100111;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111011111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011101111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011010;
SIGNAL_B = 14'b1111011100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000100111;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001110;
SIGNAL_B = 14'b1111011100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001110;
SIGNAL_B = 14'b1111011010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011110;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111011001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b1111010110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011111;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b1111010110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111010110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b1111010101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111010100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b1111010100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010011;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b1111010100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111001;
SIGNAL_B = 14'b1111010011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001001;
SIGNAL_B = 14'b1111010010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111010;
SIGNAL_B = 14'b1111001111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001010;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b1111001111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b1111001101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b1111001110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111001101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b1111001101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000010111;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001010;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001011;
SIGNAL_B = 14'b1111001100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001011;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100101;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111110;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b1111001011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100101;
SIGNAL_B = 14'b1111001010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b1111001001110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b1111001001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b1111001001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b1111001000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110110;
SIGNAL_B = 14'b1111001000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b1111000111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b1111000110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100001111;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101001;
SIGNAL_B = 14'b1111000101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111010;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010011;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b1111000010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b1111000010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b1111000001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b1111000000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001000;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100010;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110010;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111101;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b1110111101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110011;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101000001;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b1110111011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b1110111011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b1110111010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111000011;
SIGNAL_B = 14'b1110111010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b1110111001110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010000;
SIGNAL_B = 14'b1110111000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b1110111001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010001;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101100;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b1110110111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b1110110111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011110000;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001010;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010110;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101011000;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b1110110010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101011000;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b1110110010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b1110110010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110100;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000000;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111100111;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011011;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111100111;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110110;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101000;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101000;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101001;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001011101;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000100;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010010;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011011111;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010011;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111001;
SIGNAL_B = 14'b1110101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b1110101100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010100;
SIGNAL_B = 14'b1110101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111010;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b1110101011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110001001;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b1110101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111100101;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011001;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110011;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b1110100111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010000001;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b1110100111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010011011;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010101000;
SIGNAL_B = 14'b1110100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010101000;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011001111;
SIGNAL_B = 14'b1110100110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011110110;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100101010;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011110;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100101010;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011110;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111001;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111001;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110101101;
SIGNAL_B = 14'b1110100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100100011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111000111;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b1110100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100010;
SIGNAL_B = 14'b1110100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111100;
SIGNAL_B = 14'b1110100010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001100011;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001110001;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111101;
SIGNAL_B = 14'b1110100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010010111;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100100;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011100110;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001101;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001110;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b1110100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001110;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101000;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b1110011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111000100;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111101011;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010011;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000110;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111111000;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010010;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111011;
SIGNAL_B = 14'b1110011100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111010;
SIGNAL_B = 14'b1110011101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010001000;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100011;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111110;
SIGNAL_B = 14'b1110011100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b1110011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100010111;
SIGNAL_B = 14'b1110011011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b1110011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001011;
SIGNAL_B = 14'b1110011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100111;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110001101;
SIGNAL_B = 14'b1110011001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100111;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101001;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000011;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000001111;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110111;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b1110010111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b1110011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010010010;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011010011;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100001;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101001000;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101110;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100111011;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110111110;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111111111;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110100;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001101;
SIGNAL_B = 14'b1110010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110100;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010000001;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011011101;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101000110;
SIGNAL_B = 14'b1110010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100010001;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010011;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010011;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101110;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101110;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111001000;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111001000;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110001;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010111;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001010111;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001001010;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100100;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001101;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001101;
SIGNAL_B = 14'b1110010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100000001;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001110;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011101;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010000;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101101010;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101011;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110111;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110111;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b1110010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111010;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001000111;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001010101;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001111100;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100011;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010101;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111101;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001001;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100101;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001011;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100111111;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101110100;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000001;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110011010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011101;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101011;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101010;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101011;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010000110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010001;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111101;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111110;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110001;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111010;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b1110001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110111100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111010110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100101;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010000000;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100000010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000011;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011111;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110010001;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011110;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000101110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010111110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011001011;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010111110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011111111;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101001;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111110111;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001111001;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000111;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001111001;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011100001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011101110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011100001;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101100100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100111101;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001100;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110100110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101111110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101111110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b1110010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001110111;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010110111;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010001;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101011;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000110;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011111001;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100101101;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101110;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010011;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010101;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101110;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111100;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111100;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111010110;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110001;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000111111;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011001;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011010;
SIGNAL_B = 14'b1110010010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011001;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110101;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100000011;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100000011;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110110;
SIGNAL_B = 14'b1110010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101001;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101100;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111000;
SIGNAL_B = 14'b1110010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101100;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101110;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000001000;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b1110010100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000101111;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001100011;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b1110010100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b1110010101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b1110010110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b1110010101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011001;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110111;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b1110010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000101;
SIGNAL_B = 14'b1110010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011101;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001000110;
SIGNAL_B = 14'b1110010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000010010;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010001000;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111010;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001000110;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111010;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010101;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100011;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010111;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100100;
SIGNAL_B = 14'b1110011011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110010;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001100;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001100;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110011;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111101000;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111001101;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111001110;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110110;
SIGNAL_B = 14'b1110011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001011101;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b1110011100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010101011;
SIGNAL_B = 14'b1110011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010010;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010011;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100000;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100111011;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b1110011111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111101;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110000;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110001;
SIGNAL_B = 14'b1110011111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001010;
SIGNAL_B = 14'b1110100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001011;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001011;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110011;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110011;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001111;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011101;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110101;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110111;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101110;
SIGNAL_B = 14'b1110100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111001000;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100010;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b1110100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b1110100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001100;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011010;
SIGNAL_B = 14'b1110101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b1110101011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010001;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b1110101011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b1110101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010001;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b1110101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b1110101101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b1110101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010010;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101100;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111101;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b1110110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111110;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110000;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b1110110100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b1110110011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011100;
SIGNAL_B = 14'b1110110110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b1110110110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000010;
SIGNAL_B = 14'b1110110111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b1110111000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b1110111001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010100000;
SIGNAL_B = 14'b1110111001110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b1110111011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b1110111011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b1110111100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111011;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b1110111101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100000111;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101110;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b1110111101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b1110111110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1111000000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100010;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b1111000000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000000000;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000000000;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111000100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011001;
SIGNAL_B = 14'b1111000110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111000110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111000111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111001000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101010;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010001;
SIGNAL_B = 14'b1111001010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010001;
SIGNAL_B = 14'b1111001011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010001;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101011111;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101011111;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111101;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b1111011111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b1111100011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111100100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b1111101000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111110000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111110100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111110111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111111001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111111010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111111010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111111110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111100;
SIGNAL_B = 14'b0000000101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b0000001000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b0000000111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b0000001100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000001111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111100;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000010000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b0000010001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101011;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b0000010100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011111000;
SIGNAL_B = 14'b0000010110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000011000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110111;
SIGNAL_B = 14'b0000011011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000011110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000011111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000100001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110011;
SIGNAL_B = 14'b0000100001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b0000100010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001100;
SIGNAL_B = 14'b0000100010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100110;
SIGNAL_B = 14'b0000100011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110010;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b0000100100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110000;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000101000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b0000101000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100001;
SIGNAL_B = 14'b0000101001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b0000101001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b0000101001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100000111;
SIGNAL_B = 14'b0000101001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101110;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b0000101011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b0000101011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b0000101110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011111;
SIGNAL_B = 14'b0000101111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101001;
SIGNAL_B = 14'b0000101110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b0000110000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b0000110000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000110001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b0000110010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b0000110100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b0000110101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b0000110101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b0000110111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110001;
SIGNAL_B = 14'b0000110110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001011;
SIGNAL_B = 14'b0000110111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b0000111000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010111;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100011;
SIGNAL_B = 14'b0000111000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000111000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100100;
SIGNAL_B = 14'b0000111001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010110000;
SIGNAL_B = 14'b0000111010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010110;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111010;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b0000111100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111001;
SIGNAL_B = 14'b0000111010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b0000111100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111000;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010001;
SIGNAL_B = 14'b0000111110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110110111;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000001;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b0001000000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100101000;
SIGNAL_B = 14'b0001000010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100001110;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110011;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110011;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001101;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100110;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b0001000100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b0001000100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b0001000110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101110;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b0001000110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010100;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000111;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b0001001001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100111000;
SIGNAL_B = 14'b0001001001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100111000;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b0001001011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b0001001011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000011;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001001101;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111100101;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b0001001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111100101;
SIGNAL_B = 14'b0001001110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001010;
SIGNAL_B = 14'b0001001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b0001001111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001011;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111100;
SIGNAL_B = 14'b0001010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b0001010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100111011;
SIGNAL_B = 14'b0001010001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100000;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010010;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011110;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000101000;
SIGNAL_B = 14'b0001010011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001110111;
SIGNAL_B = 14'b0001010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110101;
SIGNAL_B = 14'b0001010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b0001010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111101000;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001110;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b0001010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b0001010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111101000;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110011;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111101000;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100111;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b0001010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110000;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010111;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b0001011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010110;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100011;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100010;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010101;
SIGNAL_B = 14'b0001011001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011101111;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001000;
SIGNAL_B = 14'b0001011001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111100;
SIGNAL_B = 14'b0001011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001000110;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001000110;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000101100;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001000110;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000101;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000101;
SIGNAL_B = 14'b0001011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000010001;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010000;
SIGNAL_B = 14'b0001011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110111;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101110101;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000000;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011010;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100001101;
SIGNAL_B = 14'b0001011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100001101;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011010;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111111;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100100;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b0001011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110001;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100101;
SIGNAL_B = 14'b0001011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000111100;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111011;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111000111;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101100;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110100000;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b0001100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111000;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101000100;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111000;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010001;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100000011;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110110;
SIGNAL_B = 14'b0001100010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011001111;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011100;
SIGNAL_B = 14'b0001100011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110100;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001110;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011011;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010000001;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010000000;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000111111;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000111111;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b0001100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000111111;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b0001100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111101;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110001;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001011;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001001;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010110;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b0001100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110101111;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101100001;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101110;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101100001;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000101;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101000111;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010011;
SIGNAL_B = 14'b0001100111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100100000;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011111001;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010011;
SIGNAL_B = 14'b0001100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010010;
SIGNAL_B = 14'b0001100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101010;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010011101;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010110111;
SIGNAL_B = 14'b0001100111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001000010;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000001;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001000010;
SIGNAL_B = 14'b0001101000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b0001101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111110011;
SIGNAL_B = 14'b0001100111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111110101;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001101;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110110011;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001101;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101010111;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101001010;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100111101;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101001010;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011101111;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100111101;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011101111;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011100001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010101;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111011;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011000111;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111011;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001111001;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010100;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000110;
SIGNAL_B = 14'b0001101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010001;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010001;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111110111;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000010;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000100;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111010000;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101000;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101001110;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100100110;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011111111;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011111111;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011100101;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011111110;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011111111;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110000;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100011;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001010101;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001001001;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000010100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111000110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111000;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000101;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011110;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011101000;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000000;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110010;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110010;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100011;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111010110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110010100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110111011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100001;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100100000;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101100;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101000;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101001;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100110;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100101;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110001;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111101;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111101;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001010;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010100000;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b0001110000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010100000;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010010011;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110100;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000110111;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110001110;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001100;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010101111;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001001;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001100001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001010100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000110;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101001111;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001101;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110000;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111010101;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101111010;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101011111;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010101001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010101001;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000001;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001101;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110010111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110010111;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101110000;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101010110;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100001000;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101111;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101110;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011010011;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011110;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010010010;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110111;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110111;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010000;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110001101;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110010;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b0001101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111110;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001010;
SIGNAL_B = 14'b0001101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011110001;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010101111;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010100;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010101111;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000011111;
SIGNAL_B = 14'b0001101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011101;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110011101;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010000;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101000;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101000;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011001;
SIGNAL_B = 14'b0001100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001100100;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b0001100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111011;
SIGNAL_B = 14'b0001100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100010;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100010;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101111;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b0001100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101111;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000110;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111001;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000101;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100101010;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100010001;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100010000;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011001111;
SIGNAL_B = 14'b0001100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010101000;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110011;
SIGNAL_B = 14'b0001100010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b0001100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011000;
SIGNAL_B = 14'b0001100001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110001;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110001;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110001001;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101111011;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101110;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b0001011111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111011;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010011;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010011;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111001;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010011110;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101010;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101001;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110110;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b0001011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011011;
SIGNAL_B = 14'b0001011100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b0001011100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111100111;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000001;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111110;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b0001011001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110001;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100011;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001001;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010110;
SIGNAL_B = 14'b0001011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010110;
SIGNAL_B = 14'b0001011001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001001;
SIGNAL_B = 14'b0001011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b0001011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001001;
SIGNAL_B = 14'b0001011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b0001010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000101;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010010;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b0001010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101010;
SIGNAL_B = 14'b0001010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101010;
SIGNAL_B = 14'b0001010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b0001010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101010;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b0001010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101011011;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101100111;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101000001;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100111;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100110;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110001;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110001;
SIGNAL_B = 14'b0001010010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010001010;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b0001010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001000;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b0001001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b0001001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000000111;
SIGNAL_B = 14'b0001001110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b0001001101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b0001001101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b0001001100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b0001001011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b0001001011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000010;
SIGNAL_B = 14'b0001001010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000010;
SIGNAL_B = 14'b0001000111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010101000;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b0001000111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100101;
SIGNAL_B = 14'b0001000110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110001;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b0001000100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100100;
SIGNAL_B = 14'b0001000101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111101;
SIGNAL_B = 14'b0001000011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100100;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100011;
SIGNAL_B = 14'b0001000011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100010;
SIGNAL_B = 14'b0001000100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100011111;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b0000111111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010111000;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011110;
SIGNAL_B = 14'b0000111011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b0000111010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000001;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b0000111000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b0000111001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110100;
SIGNAL_B = 14'b0000111000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000111000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000110110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001101;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010110;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000101111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000101111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000101110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111100;
SIGNAL_B = 14'b0000101110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010101;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111011;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000101101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111011;
SIGNAL_B = 14'b0000101011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b0000101010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111011;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000101000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011001000;
SIGNAL_B = 14'b0000100111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011001000;
SIGNAL_B = 14'b0000101000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100001;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000100000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b0000011111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000011111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000011101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000011110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000011011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000011001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000010111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000010111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000010011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000010001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110000001;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000001111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000001101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000001011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000001011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000000111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000000101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000000011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000000001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000000001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000110111;
SIGNAL_B = 14'b1111111101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b1111111010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000110111;
SIGNAL_B = 14'b1111111010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b1111111001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b1111111010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b1111111000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111110001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111011;
SIGNAL_B = 14'b1111110000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111110000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b1111101111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011001000;
SIGNAL_B = 14'b1111101101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b1111101101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b1111101110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b1111101101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001000;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111011;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b1111101010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111101001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010101;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001000;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100101111;
SIGNAL_B = 14'b1111100111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111100111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111100101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011001;
SIGNAL_B = 14'b1111100011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011001;
SIGNAL_B = 14'b1111100011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b1111100001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100110;
SIGNAL_B = 14'b1111100001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111000000;
SIGNAL_B = 14'b1111100001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110100;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b1111011110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100111;
SIGNAL_B = 14'b1111011110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000000;
SIGNAL_B = 14'b1111011101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110100;
SIGNAL_B = 14'b1111011101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000101;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000101;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b1111010110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101100;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b1111010101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b1111010100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000110;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b1111001111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b1111001111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110001;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111110;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b1111001101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b1111001100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b1111001001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b1111001000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011100;
SIGNAL_B = 14'b1111000111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b1111000111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000011;
SIGNAL_B = 14'b1111000111000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b1111000110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b1111000101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000001000;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010100;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000000111;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b1111000000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b1110111111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010001010;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011001;
SIGNAL_B = 14'b1110111100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b1110111101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001101;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001101;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110100;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111000011;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111000100;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011111;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101100;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b1110110111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b1110110111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101100;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b1110110110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b1110110110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b1110110100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100011;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011110000;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b1110110100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010110;
SIGNAL_B = 14'b1110110011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110001;
SIGNAL_B = 14'b1110110011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101011000;
SIGNAL_B = 14'b1110110010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101011000;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b1110110010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001011;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110011001;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000000;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111101000;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101010;
SIGNAL_B = 14'b1110101110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101010;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001011101;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101001;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000100;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010011110;
SIGNAL_B = 14'b1110101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000100;
SIGNAL_B = 14'b1110101100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b1110101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101101;
SIGNAL_B = 14'b1110101101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010010;
SIGNAL_B = 14'b1110101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010011;
SIGNAL_B = 14'b1110101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111001;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b1110101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010011;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100001;
SIGNAL_B = 14'b1110101100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101110;
SIGNAL_B = 14'b1110101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b1110101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b1110101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b1110101001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111100100;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b1110101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011001;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010101000;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010000001;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011001111;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011110111;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000100;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100110111;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111001;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011110;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000110;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111000;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111000111;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b1110100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111011;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111101;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000101111;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010011000;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010010111;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001110001;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b1110100001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011001;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011100110;
SIGNAL_B = 14'b1110100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001101;
SIGNAL_B = 14'b1110011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001111;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b1110100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110010000;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b1110011111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111111000;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010011;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100000;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100000;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010101111;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010001000;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011110000;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111101;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011110000;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100101;
SIGNAL_B = 14'b1110011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111101;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110001101;
SIGNAL_B = 14'b1110011001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011001;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100110;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b1110011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b1110011001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000011100;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110111;
SIGNAL_B = 14'b1110011001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000010;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101010;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000010;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b1110011001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001000011;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000110;
SIGNAL_B = 14'b1110011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011110;
SIGNAL_B = 14'b1110011000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010010001;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011100000;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011010011;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011010011;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101110;
SIGNAL_B = 14'b1110010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101100010;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101111101;
SIGNAL_B = 14'b1110010111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101111101;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001101;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011010;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110100;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001110;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000001;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110100;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001101000;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010101000;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010101001;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011011101;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011111000;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101000101;
SIGNAL_B = 14'b1110010101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110100001;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110100001;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000001001;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111010101;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111101111;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110001;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000100011;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110000;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001011;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001001011;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010111111;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001101;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001110;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100000001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101000011;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101000010;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011100;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011100;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110000100;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101011;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000100000;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000100000;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001010101;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000100001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111011;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001001;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001011;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110001;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001100;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001100;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110011011;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001100;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110011011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110100111;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011101;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001000100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101010;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001011110;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010000110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010010011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111100;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111101;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011000;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100110;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011100;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000010;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000011;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010000;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010011;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010100;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100001;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110010101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001100;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001011;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110011;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101010000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000101111;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010010110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011011000;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b1110001110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100100110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110110101;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b1110001111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000111;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010100;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111011;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010101;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011101111;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101001010;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111000000;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001100;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000110101;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000100;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001110110;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010001;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010001;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011101011;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000110;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011111001;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100100000;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100100000;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010101;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b1110010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101110;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111010110;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111010111;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000010111;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010000000;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110100;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110110;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011110;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100001111;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011110;
SIGNAL_B = 14'b1110010011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110011111;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000001000;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100000;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101110;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010100;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000101111;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b1110010110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011010;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101110110;
SIGNAL_B = 14'b1110010110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101001;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110111;
SIGNAL_B = 14'b1110010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111000011;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011101;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011101;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101110;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010010100;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100010;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100001010;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100100;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b1110011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001100;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110000000;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001101;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011010;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110100;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000001;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111110101;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b1110011100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010010;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010101011;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b1110011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110010110;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110000;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111110;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111110;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110001;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100110;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100101;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b1110100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b1110100000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101001;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011100;
SIGNAL_B = 14'b1110100010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011100;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b1110100100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010011;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b1110100101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100010;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000010110;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b1110100111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b1110100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b1110100111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001001;
SIGNAL_B = 14'b1110100111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b1110101000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001100;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110011;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b1110101001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011010;
SIGNAL_B = 14'b1110101001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000001;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100101000;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110101;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b1110101010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000101;
SIGNAL_B = 14'b1110101100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b1110101100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010010;
SIGNAL_B = 14'b1110101100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000101;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011111;
SIGNAL_B = 14'b1110101100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000110;
SIGNAL_B = 14'b1110101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011111;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b1110101110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000011111;
SIGNAL_B = 14'b1110101111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010110000;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001010;
SIGNAL_B = 14'b1110110000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010111;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110001;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111110;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110001;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b1110110011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b1110110011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b1110110101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b1110110110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101001;
SIGNAL_B = 14'b1110110111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b1110111000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110110;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b1110111001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b1110111001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b1110111010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101110;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b1110111101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101110;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b1110111101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b1110111110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1110111111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110010;
SIGNAL_B = 14'b1111000000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110011;
SIGNAL_B = 14'b1111000010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110011;
SIGNAL_B = 14'b1111000010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b1111000011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b1111000011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111000101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110011;
SIGNAL_B = 14'b1111000110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111000110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011010;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b1111001011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110111;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110111;
SIGNAL_B = 14'b1111001100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000101;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b1111001110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b1111001111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101011;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111011000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111011001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111101;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b1111011100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111100000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111100100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111100110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111101000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111101000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111101010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111110010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111110;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111111110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111111101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b0000000010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b0000000100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b0000000110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b0000001000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000001000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b0000001001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000001001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000010000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000010001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101011;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b0000010011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101011;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b0000010101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000010101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b0000010101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000010110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000000;
SIGNAL_B = 14'b0000011101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b0000011111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b0000011111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000000000;
SIGNAL_B = 14'b0000100001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001100;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001100;
SIGNAL_B = 14'b0000100101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b0000100100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b0000101000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101110;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b0000101001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b0000101001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b0000101001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b0000101011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111011;
SIGNAL_B = 14'b0000101010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010100;
SIGNAL_B = 14'b0000101011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111010;
SIGNAL_B = 14'b0000101100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b0000101011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000111;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b0000101100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000101111000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010100000;
SIGNAL_B = 14'b0000101110110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b0000101110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b0000101111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b0000101111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000011;
SIGNAL_B = 14'b0000101111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b0000101111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b0000110000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101001;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000110000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101001;
SIGNAL_B = 14'b0000110010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b0000110011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b0000110101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b0000110101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000110110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001011;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111110;
SIGNAL_B = 14'b0000110110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001010;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110000;
SIGNAL_B = 14'b0000110111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010111;
SIGNAL_B = 14'b0000111000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b0000111000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b0000111000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b0000111001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b0000111100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010011;
SIGNAL_B = 14'b0000111011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000110;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111010;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111010;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b0000111101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101100;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110111000;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010010;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011110;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0000111111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000001;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b0001000001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100100111;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b0001000000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110100;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001100;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011010;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001100;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b0001000010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001100;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b0001000110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b0001000110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b0001000110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b0001000111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101110;
SIGNAL_B = 14'b0001000110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010011;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b0001000111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b0001001000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001001001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100111000;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000100;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110111;
SIGNAL_B = 14'b0001001010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011010000;
SIGNAL_B = 14'b0001001011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b0001001100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b0001001011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b0001001100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001001101;
SIGNAL_B = 14'b0001001101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000111111;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b0001001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b0001001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001011;
SIGNAL_B = 14'b0001001110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111111;
SIGNAL_B = 14'b0001001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110000;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110111101;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b0001010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111100;
SIGNAL_B = 14'b0001010000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110010110;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111101;
SIGNAL_B = 14'b0001001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b0001010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101101;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010011;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101101;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000110;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011110;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010010;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110110;
SIGNAL_B = 14'b0001010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b0001010100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111001110;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110101;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b0001010101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111001101;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110010;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111101;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010111;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110010;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100100;
SIGNAL_B = 14'b0001010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100001010;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100011;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010000111;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010000111;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100001;
SIGNAL_B = 14'b0001011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111010;
SIGNAL_B = 14'b0001011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010010101;
SIGNAL_B = 14'b0001011010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010000111;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000010010;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111110111;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111000011;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010000;
SIGNAL_B = 14'b0001011101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000010;
SIGNAL_B = 14'b0001011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000010;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101000;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011010;
SIGNAL_B = 14'b0001011101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b0001011101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100001100;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b0001011111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011111111;
SIGNAL_B = 14'b0001011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110001;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001100011;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100100;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100001;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000101111;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000111100;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111011;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010110;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000001000;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101101;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101100;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111000111;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000110;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000101;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010001;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010001;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101000100;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110110;
SIGNAL_B = 14'b0001100010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101001;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011100;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011100;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011011;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011001111;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100110;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011010;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100110;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111101;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111110;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000010111;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111100011;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110001;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111101;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110101111;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010101;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b0001100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010101;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100100000;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000101;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010111000;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010011110;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101010;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010001;
SIGNAL_B = 14'b0001100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010111000;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010110111;
SIGNAL_B = 14'b0001100111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101010;
SIGNAL_B = 14'b0001100111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000101000;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000110101;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b0001100111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111110100;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100110;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100110;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110110010;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011001;
SIGNAL_B = 14'b0001101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110000;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100111101;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b0001101001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010100000;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010101;
SIGNAL_B = 14'b0001101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010100;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101101;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101101;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010100000;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010011;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001011111;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010000;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111110110;
SIGNAL_B = 14'b0001101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111010000;
SIGNAL_B = 14'b0001101011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101001;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000010;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101101000;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011111110;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011111111;
SIGNAL_B = 14'b0001101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011100101;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001001;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010010110;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001110000;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111101;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001010101;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010011;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111000101;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011110;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111000101;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100000010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100011100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011001;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001111111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100101;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000110001;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111111101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111111101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110111011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110000111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110010100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010000;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101001;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000010;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010001111;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011011;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011001;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110010;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110010111;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001001;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100110000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100010;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101100;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010000101;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001011110;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010000110;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000111000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110001101;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b0001110000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001000;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000100000;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111000101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111010010;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110110;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101101010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100101000;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100000001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001100;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100101;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110010;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001001010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000100011;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111010101;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101111010;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101010;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011011;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001011011;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111111111;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001001;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110010111;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101001000;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100010;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011100000;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010010010;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010010010;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011110;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110110;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111110110;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101001;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100110;
SIGNAL_B = 14'b0001101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110001101;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100101;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101011001;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100011;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111101;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010101111;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010000111;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001101110;
SIGNAL_B = 14'b0001101001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010000111;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111010;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010010;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000011111;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111111000;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111101100;
SIGNAL_B = 14'b0001101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110001111;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101000001;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001110;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001101;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b0001100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b0001100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010011000;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001110001;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111101;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001001010;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100010;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111100;
SIGNAL_B = 14'b0001100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100010;
SIGNAL_B = 14'b0001100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010011;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111000;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100110111;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100101010;
SIGNAL_B = 14'b0001100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011101010;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b0001100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001110;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011001;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110011;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b0001100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110001;
SIGNAL_B = 14'b0001100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111100100;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111100100;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110001;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101111011;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111011;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b0001011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010011;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111001;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b0001011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011100000;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b0001011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010011110;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110110;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001011101;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000100;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b0001011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110101;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011011;
SIGNAL_B = 14'b0001011100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b0001011100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001101;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b0001011011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101011000;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111101;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011110000;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111100;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001011111;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111000;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101011;
SIGNAL_B = 14'b0001010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111000;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011111;
SIGNAL_B = 14'b0001010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011110;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110111;
SIGNAL_B = 14'b0001010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010000;
SIGNAL_B = 14'b0001010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110011;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100111;
SIGNAL_B = 14'b0001010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100110;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100110;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010001010;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b0001010001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b0001010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001000;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101110;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111010;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000000111;
SIGNAL_B = 14'b0001001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000000111;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101110;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111010;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010100;
SIGNAL_B = 14'b0001001101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101101;
SIGNAL_B = 14'b0001001101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101101;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b0001001100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b0001001100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b0001001011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101001;
SIGNAL_B = 14'b0001001001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000011;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100001111;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000010;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b0001001001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b0001000111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b0001000110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b0001000110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b0001000100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100100;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110110000;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100010;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b0001000010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b0001000000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111001;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101100;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b0001000000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101100;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0000111111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101100;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b0000111101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b0000111101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011011;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110100;
SIGNAL_B = 14'b0000111001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110100;
SIGNAL_B = 14'b0000111000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110100;
SIGNAL_B = 14'b0000111000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000111000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000001;
SIGNAL_B = 14'b0000111000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000111000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000111000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000110110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111000000;
SIGNAL_B = 14'b0000110110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b0000110101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001101;
SIGNAL_B = 14'b0000110011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b0000110010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110000;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000101111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000101110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000101111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010101;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111100;
SIGNAL_B = 14'b0000101110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b0000101101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010101;
SIGNAL_B = 14'b0000101100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000101010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000101001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000101001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011001000;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b0000101000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000100110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000100010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000011100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000011010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000011001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000011000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b0000010111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000010101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000010011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110001110;
SIGNAL_B = 14'b0000001011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000001010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000001010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b1111111111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b1111111111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b1111111011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111111010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001100000;
SIGNAL_B = 14'b1111111001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b1111110111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111110111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111110110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b1111110100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111110100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111011;
SIGNAL_B = 14'b1111110001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011001000;
SIGNAL_B = 14'b1111110000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101110;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101110;
SIGNAL_B = 14'b1111110001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111110000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111110000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111011;
SIGNAL_B = 14'b1111101110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b1111101110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b1111101101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b1111101101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001000;
SIGNAL_B = 14'b1111101011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b1111101100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b1111101001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b1111101010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111101001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111101001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100101111;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111100111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110011;
SIGNAL_B = 14'b1111100011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100110;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111100001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111100001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011010;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100111;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011010;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111011101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001110;
SIGNAL_B = 14'b1111011100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b1111011010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111011000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011110;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010010;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111010111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b1111010110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111010110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b1111010110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111001;
SIGNAL_B = 14'b1111010101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100011111;
SIGNAL_B = 14'b1111010100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b1111010100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b1111010100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010011;
SIGNAL_B = 14'b1111010100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100000;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b1111010001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111101;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111001111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111101;
SIGNAL_B = 14'b1111001111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001010;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001010;
SIGNAL_B = 14'b1111001110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b1111001110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100100;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111110;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b1111001010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b1111000111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b1111001000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b1111000111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011101;
SIGNAL_B = 14'b1111000110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b1111000110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101010;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b1111000110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101101;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100001;
SIGNAL_B = 14'b1111000011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111010;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101110;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b1111000001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001000;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001101111;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100110;
SIGNAL_B = 14'b1110111110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100110;
SIGNAL_B = 14'b1110111101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b1110111100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b1110111101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100111;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b1110111100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101011011;
SIGNAL_B = 14'b1110111100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110101;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110111;
SIGNAL_B = 14'b1110111010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010000;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011110;
SIGNAL_B = 14'b1110111000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b1110111000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010010;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101100;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010010;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111000;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b1110110111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b1110110101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b1110110110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001011111;
SIGNAL_B = 14'b1110110110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111101;
SIGNAL_B = 14'b1110110101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b1110110101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b1110110011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b1110110100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001001;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b1110110100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111101;
SIGNAL_B = 14'b1110110011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b1110110010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b1110110001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110101;
SIGNAL_B = 14'b1110110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000001;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011011;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110101;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001011101;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001011101;
SIGNAL_B = 14'b1110101110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b1110101110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010011110;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000011;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010010;
SIGNAL_B = 14'b1110101101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100001;
SIGNAL_B = 14'b1110101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111010;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111010;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101000111;
SIGNAL_B = 14'b1110101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b1110101100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b1110101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101111100;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110001001;
SIGNAL_B = 14'b1110101010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b1110101001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111001010;
SIGNAL_B = 14'b1110101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011000;
SIGNAL_B = 14'b1110101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000111111;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111111;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001101;
SIGNAL_B = 14'b1110101000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b1110100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001001101;
SIGNAL_B = 14'b1110100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100110;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b1110100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b1110100110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011010000;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011101010;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100101010;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011110;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111000;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b1110100101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111000;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110101101;
SIGNAL_B = 14'b1110100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b1110100010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b1110100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101111;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111100;
SIGNAL_B = 14'b1110100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111101;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001010;
SIGNAL_B = 14'b1110100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111101;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111101;
SIGNAL_B = 14'b1110100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001010;
SIGNAL_B = 14'b1110100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011100110;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101000010;
SIGNAL_B = 14'b1110100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100100111;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101000010;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111011;
SIGNAL_B = 14'b1110011101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111011;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001101110;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010001000;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010100;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b1110011101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001010;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b1110011011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b1110011011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001011;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b1110011011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100111;
SIGNAL_B = 14'b1110011011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000010;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b1110011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111110100;
SIGNAL_B = 14'b1110011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000011;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000011100;
SIGNAL_B = 14'b1110011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000001111;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b1110011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101010;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001110111;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b1110011000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010101100;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b1110011000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011010011;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011100000;
SIGNAL_B = 14'b1110011000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100001000;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100111100;
SIGNAL_B = 14'b1110010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101101111;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101010110;
SIGNAL_B = 14'b1110010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101001000;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110010111;
SIGNAL_B = 14'b1110010110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110100100;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b1110010101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111111111;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110100;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001101;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010000010;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001101000;
SIGNAL_B = 14'b1110010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011011101;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b1110010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101111010;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111010101;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101110;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101110;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111101111;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000001001;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110000;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011000;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000111101;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001011;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011110100;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001110;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100000010;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001110;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101101010;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101001111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011100;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110000100;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101001111;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101011;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000010100;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000010100;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111010;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111011;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100011;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100010;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100011;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100011;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010101111;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111101;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010110;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101011001;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101110100;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001100;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110001110;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110001110;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110001110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000110111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001000100;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010000110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100110000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010111;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110010111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011001;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011011;
SIGNAL_B = 14'b1110001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110110;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011011110;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101100;
SIGNAL_B = 14'b1110001100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111011;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111011;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110010101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111110000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100101;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111111101;
SIGNAL_B = 14'b1110001101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110010;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010000000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011101000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101101010;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000010;
SIGNAL_B = 14'b1110001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110010001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000010100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000101110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001010101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010010110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011011000;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101001;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110110101;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000100;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000111000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001111010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000110;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111011;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010101;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011101111;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101001010;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101010111;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101010111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111000000;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001110110;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010011110;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101010;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010111000;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000101;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010010;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010011;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100100000;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111101;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001010;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001010;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001011;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000111111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100110;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100111;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011010;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101001;
SIGNAL_B = 14'b1110010001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110110;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b1110010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b1110010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101000100;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000110;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111000;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110011111;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111010;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000101111;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000111100;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b1110010100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110001;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011011001;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011011001;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100100111;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b1110010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011101;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b1110011000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000100;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011110;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b1110011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100001;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010101;
SIGNAL_B = 14'b1110011001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010110;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b1110011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100011;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110010;
SIGNAL_B = 14'b1110011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b1110011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b1110011011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110011;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111100111;
SIGNAL_B = 14'b1110011011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000010;
SIGNAL_B = 14'b1110011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b1110011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001011101;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011110;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001110111;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111010;
SIGNAL_B = 14'b1110011101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100111011;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b1110011101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100111010;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111100;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110111101;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110001;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111011000;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111100101;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110001;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000111111;
SIGNAL_B = 14'b1110100001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100110;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110101;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110101;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011010000;
SIGNAL_B = 14'b1110100010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110111;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110111;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b1110100100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010011;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111001000;
SIGNAL_B = 14'b1110100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b1110100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b1110100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b1110100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b1110101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011010;
SIGNAL_B = 14'b1110101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100001110;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011010;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100101000;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100100111;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001110;
SIGNAL_B = 14'b1110101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b1110101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110110111;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110111000;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111010;
SIGNAL_B = 14'b1110101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111010;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b1110110000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010111;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111110;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010110000;
SIGNAL_B = 14'b1110110001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110000;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110000;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011000;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b1110110011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b1110110100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011100;
SIGNAL_B = 14'b1110110110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b1110110110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b1110110111000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b1110111000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b1110111001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110110;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b1110111001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011101;
SIGNAL_B = 14'b1110111010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b1110111001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101101;
SIGNAL_B = 14'b1110111010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010100000;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010100000;
SIGNAL_B = 14'b1110111011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111010;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101110;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b1110111101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b1110111101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111011;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100010;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111111;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011001;
SIGNAL_B = 14'b1111000100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111111;
SIGNAL_B = 14'b1111000010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100110;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011010;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111001000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b1111001001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110111;
SIGNAL_B = 14'b1111001001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000100;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010001;
SIGNAL_B = 14'b1111001110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b1111001110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111001111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101011;
SIGNAL_B = 14'b1111010001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b1111010111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b1111011110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111100010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111100101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111100111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111100111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111101000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b1111101000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111101001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111101100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111101111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110011001100;
SIGNAL_B = 14'b1111110000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011000;
SIGNAL_B = 14'b1111110000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110100;
SIGNAL_B = 14'b1111110100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111111000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111111011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111111111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b0000000000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b0000000001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b0000000100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000000101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000000111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000001000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b0000001010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000010000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101011111;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b0000010011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b0000010100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b0000010101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b0000010100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101011;
SIGNAL_B = 14'b0000010110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b0000010111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101011;
SIGNAL_B = 14'b0000010111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011110;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010001;
SIGNAL_B = 14'b0000011001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101010;
SIGNAL_B = 14'b0000011100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b0000011101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b0000011110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011010;
SIGNAL_B = 14'b0000011110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b0000011110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b0000011111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000011111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001101;
SIGNAL_B = 14'b0000011111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000100001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100001110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011001;
SIGNAL_B = 14'b0000100011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100110;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110010;
SIGNAL_B = 14'b0000100011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110010;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b0000100101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b0000100100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000100101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010110;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000100111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000100111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b0000101010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b0000101001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100001;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b0000101011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b0000101011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111011;
SIGNAL_B = 14'b0000101011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b0000101011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b0000101101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b0000101110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000101110110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000101111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b0000101111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b0000101110110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b0000110000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b0000110001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011100;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b0000110010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b0000110011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011011;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b0000110110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100010111;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100100;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001011;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000110111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001010;
SIGNAL_B = 14'b0000111000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b0000111000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b0000111000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b0000111010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111010;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b0000111101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000110;
SIGNAL_B = 14'b0000111110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101100;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b0000111110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011111;
SIGNAL_B = 14'b0000111110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000101;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b0000111111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110110111;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110101;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110100;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011011;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100101000;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100001101;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011011;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110011;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b0001000010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011000000;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b0001000010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011000000;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001010;
SIGNAL_B = 14'b0001000101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b0001000110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000010101;
SIGNAL_B = 14'b0001000110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b0001000110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000010110;
SIGNAL_B = 14'b0001000110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b0001001000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b0001001000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b0001001001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100001;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100111000;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000011;
SIGNAL_B = 14'b0001001010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011010000;
SIGNAL_B = 14'b0001001100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110110;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011011;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b0001001100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b0001001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001001101;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011000;
SIGNAL_B = 14'b0001001110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b0001001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b0001001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110111101;
SIGNAL_B = 14'b0001010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110001;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001010;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b0001010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110010110;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111101;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b0001010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101101;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010011;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100000111;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b0001010010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111001;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b0001010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111010;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010010;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011110;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001011101;
SIGNAL_B = 14'b0001010011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010101011;
SIGNAL_B = 14'b0001010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000010;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000010;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100111;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000001;
SIGNAL_B = 14'b0001010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101111111;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110010;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101111111;
SIGNAL_B = 14'b0001010110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100001010;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111100;
SIGNAL_B = 14'b0001011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100010111;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100011;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001000;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010101111;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101110;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000101100;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000010010;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011111;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011110;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000101100;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011111;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110111;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b0001011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b0001011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100001101;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011010;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100001101;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111111;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100101;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001100011;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000101111;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101110;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101110;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111000111;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101100;
SIGNAL_B = 14'b0001100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101100;
SIGNAL_B = 14'b0001100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b0001100011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011111;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b0001100010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100001111;
SIGNAL_B = 14'b0001100011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101001;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011011;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011011;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011010;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011001;
SIGNAL_B = 14'b0001100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b0001100101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b0001100011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001010;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001011;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110001;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000011000;
SIGNAL_B = 14'b0001100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111100011;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111101;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001010;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111100;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111100;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101000111;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101000111;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000101;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000110;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011111;
SIGNAL_B = 14'b0001100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010010;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010001;
SIGNAL_B = 14'b0001100110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000100;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101010;
SIGNAL_B = 14'b0001100111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010000;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001011100;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001110110;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111110100;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b0001100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000000;
SIGNAL_B = 14'b0001101000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000001;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110110011;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111000000;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111000000;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011001;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101100100;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101100100;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100111101;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011101111;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101001010;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011100001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000110;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001111010;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000111;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001100000;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010001;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000111000;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000100;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011101;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111110111;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111010000;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000010;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011100;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101001101;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101000000;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011011000;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110000;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011011000;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011010111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100100;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001001;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100100;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001001000;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100010;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000010100;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000000111;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111000110;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011111;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101111000;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101101010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101010000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100011100;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110100;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b0001101110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010001100;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110010;
SIGNAL_B = 14'b0001101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001011;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000110001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000001010;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110001000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110000111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110000111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100001;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000011;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000010;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110101;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001111;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011010;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100101;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110010;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110010;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110001;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111101;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100000;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011010011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010000101;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111001;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011011;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110011011;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101011001;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000101101;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111000101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101011;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110111;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110000100;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100000001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010111;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111101;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100010001;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011011101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010110110;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010001111;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110100;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110000;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110100100;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101110000;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101110000;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101111;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100010100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011110;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010101100;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000100;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000100;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000010;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110111;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101000;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100101;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101011001;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100010111;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111110;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111110;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001101110;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111011;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010101111;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001101110;
SIGNAL_B = 14'b0001101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b0001101000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000100000;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b0001101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110011101;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110010000;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000010;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100101000;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110100;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b0001100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011100111;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111110;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111110;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111101;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111101;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111010;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001001;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010101;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111000111;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010010;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000110;
SIGNAL_B = 14'b0001100011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000110;
SIGNAL_B = 14'b0001100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111001;
SIGNAL_B = 14'b0001100011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000100;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100110111;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011101001;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010000001;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001001101;
SIGNAL_B = 14'b0001100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011001;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b0001100010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000111111;
SIGNAL_B = 14'b0001100010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111001010;
SIGNAL_B = 14'b0001100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110001;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101111100;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100000;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111011;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011011111;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000110;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b0001011111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000110;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110111;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001011101;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b0001011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011011;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000010;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000001;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b0001011011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001101;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111110;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b0001011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001001;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b0001011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111011;
SIGNAL_B = 14'b0001011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b0001011000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001011111;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b0001010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101011;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011111;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101010;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011111;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b0001010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b0001010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110100;
SIGNAL_B = 14'b0001010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101011011;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101011010;
SIGNAL_B = 14'b0001010011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001101;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001101;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b0001010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100110;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011001;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b0001010001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100010;
SIGNAL_B = 14'b0001010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111010;
SIGNAL_B = 14'b0001001111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010010;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111011;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101010;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b0001001100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000011;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b0001001010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101001;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b0001000111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111110;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100100;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b0001000101111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b0001000100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b0001000100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110001;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b0001000011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111011;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b0001000010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b0001000010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110000111;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010011;
SIGNAL_B = 14'b0001000000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100011111;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010010;
SIGNAL_B = 14'b0000111111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b0000111111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b0000111101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011110;
SIGNAL_B = 14'b0000111101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010001111;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b0000111011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011011;
SIGNAL_B = 14'b0000111001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b0000111001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000111000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110100;
SIGNAL_B = 14'b0000110111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b0000110111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110100;
SIGNAL_B = 14'b0000110110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110011;
SIGNAL_B = 14'b0000110111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b0000110101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111000000;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100110;
SIGNAL_B = 14'b0000110011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011001;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010110;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010110;
SIGNAL_B = 14'b0000110000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001001;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b0000110000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000101111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000101110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111100;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b0000101110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111011;
SIGNAL_B = 14'b0000101011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101110;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000100110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000100110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000011010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110000001;
SIGNAL_B = 14'b0000010001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000001010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000001011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011100;
SIGNAL_B = 14'b0000001000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000000110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000000101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000000110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000000100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000000100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000000001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b1111111111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b1111111100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111111100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b1111111010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b1111111001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b1111111001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111110111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b1111110110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111110101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b1111110011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100001;
SIGNAL_B = 14'b1111110010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b1111110010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b1111101111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b1111101111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111110000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111011;
SIGNAL_B = 14'b1111101110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b1111101101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b1111101101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b1111101011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111101010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100101111;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111101001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b1111100111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100101111;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001001;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011010;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111100000101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000000;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011010;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011010;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b1111011101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011011;
SIGNAL_B = 14'b1111011011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011110;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101011;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111011000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b1111011000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111011000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b1111010101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100011111;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b1111010100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000110;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b1111010100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b1111010011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b1111010001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b1111010000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100100;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110001;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b1111001111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001010;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b1111001110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b1111001100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b1111001011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100101;
SIGNAL_B = 14'b1111001010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000010;
SIGNAL_B = 14'b1111001001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011100;
SIGNAL_B = 14'b1111000110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b1111000110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000110110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101110111;
SIGNAL_B = 14'b1111000011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101101;
SIGNAL_B = 14'b1111000011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b1111000010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010100;
SIGNAL_B = 14'b1111000001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b1111000000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001101111;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b1111000000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110010;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001100;
SIGNAL_B = 14'b1110111110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100000000;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110100;
SIGNAL_B = 14'b1110111011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111000011;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010000;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010001;
SIGNAL_B = 14'b1110111001110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011111;
SIGNAL_B = 14'b1110111000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b1110111001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111000;
SIGNAL_B = 14'b1110110110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101100;
SIGNAL_B = 14'b1110110111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101100;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b1110110111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111001;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b1110110101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101100;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b1110110110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b1110110101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011110000;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b1110110100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111101;
SIGNAL_B = 14'b1110110100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111110;
SIGNAL_B = 14'b1110110100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010110;
SIGNAL_B = 14'b1110110011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001010;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110001;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110011001;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101011000;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b1110110010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001110;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001101;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b1110110000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011011;
SIGNAL_B = 14'b1110110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b1110110000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110110;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110110;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000100;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110111;
SIGNAL_B = 14'b1110101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110111;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010010;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010011;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100000;
SIGNAL_B = 14'b1110101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111011;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b1110101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111011;
SIGNAL_B = 14'b1110101011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b1110101010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011000;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000111111;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001001101;
SIGNAL_B = 14'b1110101000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b1110101000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b1110101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010000001;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010000001;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001101;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011110110;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011010000;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011001111;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100010000;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100110111;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100101010;
SIGNAL_B = 14'b1110100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101010010;
SIGNAL_B = 14'b1110100100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b1110100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110101101;
SIGNAL_B = 14'b1110100100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110101101;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b1110100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100010;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b1110100011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000101111;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100011;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001100100;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111110;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b1110100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b1110100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011010;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011100111;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011100110;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001111;
SIGNAL_B = 14'b1110011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001111;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011011;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001111;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110011100;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110101010;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111101011;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111111000;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111101100;
SIGNAL_B = 14'b1110011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010010;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000100000;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001101110;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111011;
SIGNAL_B = 14'b1110011100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010000111;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010100010;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100100;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100100;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111110;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100010111;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100101;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110001;
SIGNAL_B = 14'b1110011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101011001;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100101;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101000;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100111;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b1110011010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000010;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101001;
SIGNAL_B = 14'b1110011001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000001111;
SIGNAL_B = 14'b1110011001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110110;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b1110011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011110;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010101011;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010101011;
SIGNAL_B = 14'b1110011000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010101100;
SIGNAL_B = 14'b1110010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111011;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100001;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101001000;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101110;
SIGNAL_B = 14'b1110010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100111011;
SIGNAL_B = 14'b1110010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101110000;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b1110010111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001001;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101101111;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110100100;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b1110010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011001;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001101000;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b1110010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010001111;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010110110;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000101;
SIGNAL_B = 14'b1110010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100010001;
SIGNAL_B = 14'b1110010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011110111;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101100000;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b1110010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000110;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110100000;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000110;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111001000;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000110;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111101111;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111001000;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000001001;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000111110;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000111110;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100100;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110001;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001010111;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010001011;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001101;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100101000;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101001111;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101010000;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011100;
SIGNAL_B = 14'b1110010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110111;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110111;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000010100;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000100000;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000110;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111010;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001000111;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001000111;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001000;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001000;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111100;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001011;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100111111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101110100;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001101;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000001;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011101;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001000100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001000100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001000101;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010000110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010011111;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010010011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011010100;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b1110001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111100;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101111110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011000;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011011;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110101;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b1110001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111010;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111011;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110001000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110111100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111101111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111110000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111110000;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111111;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010001101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010000000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011101000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101010001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000101110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100010;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001100011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001010101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110000;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011001011;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011010111;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100100110;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101001101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011101;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111110111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111110111;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000100;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001011111;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010100001;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011001000;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101100100;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110100110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001101;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111110100;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000110101;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001011100;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001011100;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001011101;
SIGNAL_B = 14'b1110010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010010;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011110;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011111;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011101100;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010011;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101000111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001001;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110001;
SIGNAL_B = 14'b1110010010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111110;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000011000;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011001;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100111;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b1110010010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110100;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010101000;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101001;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b1110010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100011100;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b1110010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101110;
SIGNAL_B = 14'b1110010100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000000111;
SIGNAL_B = 14'b1110010100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000111100;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b1110010101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011011001;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100110100;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101000;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110010000;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b1110010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110011101;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b1110010111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011111;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000101;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010001000;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010001000;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100001;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010010100;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010101110;
SIGNAL_B = 14'b1110011001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110000;
SIGNAL_B = 14'b1110011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110000;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101111111;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b1110011011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100111;
SIGNAL_B = 14'b1110011010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b1110011011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b1110011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111110100;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110110;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001011101;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000110;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100000111;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b1110011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111010;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111100;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001010;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100011;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011001;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111111;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b1110100001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001001101;
SIGNAL_B = 14'b1110100010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111110;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b1110100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b1110100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b1110100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000011;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b1110100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000011;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110111;
SIGNAL_B = 14'b1110100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011100;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b1110100011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100001;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100001;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101101;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000010110;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b1110100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b1110100111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b1110101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b1110101001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000000;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100101000;
SIGNAL_B = 14'b1110101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b1110101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100100111;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000001;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110101;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011110;
SIGNAL_B = 14'b1110101011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011111;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b1110101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b1110101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000011111;
SIGNAL_B = 14'b1110101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000110;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010011;
SIGNAL_B = 14'b1110110000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110101111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001010;
SIGNAL_B = 14'b1110110001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001010;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111110;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110001;
SIGNAL_B = 14'b1110110011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b1110110010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001011;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b1110110011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b1110110100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000001;
SIGNAL_B = 14'b1110110011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011011;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b1110110101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110101000;
SIGNAL_B = 14'b1110110110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b1110110111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000010;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b1110111001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010100000;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b1110111100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010100;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100001;
SIGNAL_B = 14'b1110111101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111011;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1110111110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1111000000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b1111000000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b1111000011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000000000;
SIGNAL_B = 14'b1111000011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111000110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011010;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111000110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b1111000111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011101;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b1111001010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010001;
SIGNAL_B = 14'b1111001011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010001;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b1111001111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111001111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111011000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111011001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b1111011010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111011100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111101;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b1111100000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111100011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111100110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111101000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111101000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111101011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111101100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111110000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111110101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111110111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110011;
SIGNAL_B = 14'b1111110111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111111000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b0000000000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b0000000010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000001000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000001010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b0000001010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b0000001100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000010001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000010010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101011;
SIGNAL_B = 14'b0000010011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101011;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011111000;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010001;
SIGNAL_B = 14'b0000010100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000010111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000010110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000011000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000010111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000100;
SIGNAL_B = 14'b0000011010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000011010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000011111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000100000000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110011;
SIGNAL_B = 14'b0000011111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000100001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110011;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b0000100010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111111;
SIGNAL_B = 14'b0000100001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001100;
SIGNAL_B = 14'b0000100011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b0000100100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110010;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b0000100101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100010;
SIGNAL_B = 14'b0000100111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000100111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001000;
SIGNAL_B = 14'b0000101001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111011;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b0000101001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100000111;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b0000101010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b0000101011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b0000101100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111010;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b0000101101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b0000101101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b0000101110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000011;
SIGNAL_B = 14'b0000101111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010000;
SIGNAL_B = 14'b0000110000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010010;
SIGNAL_B = 14'b0000110000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b0000110001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110110;
SIGNAL_B = 14'b0000110010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110110;
SIGNAL_B = 14'b0000110011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000010;
SIGNAL_B = 14'b0000110011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110100101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110101000;
SIGNAL_B = 14'b0000110100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b0000110110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b0000110110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110010;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110000;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111110;
SIGNAL_B = 14'b0000111000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000111000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110000;
SIGNAL_B = 14'b0000111000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111011;
SIGNAL_B = 14'b0000111000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001010;
SIGNAL_B = 14'b0000111010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b0000111001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001001;
SIGNAL_B = 14'b0000111011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b0000111100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001010100;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111101000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000110;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010001;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110110111;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110100;
SIGNAL_B = 14'b0001000010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011010;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b0001000010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001101;
SIGNAL_B = 14'b0001000011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b0001000100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100010;
SIGNAL_B = 14'b0001000101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000101111;
SIGNAL_B = 14'b0001000110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b0001000110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b0001000110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101110;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010011;
SIGNAL_B = 14'b0001000110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111011;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101101;
SIGNAL_B = 14'b0001000111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010011;
SIGNAL_B = 14'b0001000111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b0001001001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100111000;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b0001001010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000011;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b0001001100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b0001001100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011100;
SIGNAL_B = 14'b0001001011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011101;
SIGNAL_B = 14'b0001001100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110101;
SIGNAL_B = 14'b0001001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011011;
SIGNAL_B = 14'b0001001100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001110;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011011;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110010;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110010;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100110;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111111;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001010;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110000;
SIGNAL_B = 14'b0001010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110000;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101101111;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111100;
SIGNAL_B = 14'b0001010000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100111011;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100000110;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100000110;
SIGNAL_B = 14'b0001010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111010;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b0001010011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101100;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010010;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b0001010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000100;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b0001010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000101001;
SIGNAL_B = 14'b0001010100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b0001010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000101001;
SIGNAL_B = 14'b0001010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b0001010100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b0001010100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000010;
SIGNAL_B = 14'b0001010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111101000;
SIGNAL_B = 14'b0001010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110011;
SIGNAL_B = 14'b0001010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110011;
SIGNAL_B = 14'b0001010110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110011;
SIGNAL_B = 14'b0001010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110010;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101111111;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b0001011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100100;
SIGNAL_B = 14'b0001010111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100100;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b0001010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100001010;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011100010;
SIGNAL_B = 14'b0001011001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100001;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001000;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111010;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100010;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001010011;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b0001011010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000101100;
SIGNAL_B = 14'b0001011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000010001;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000110;
SIGNAL_B = 14'b0001011011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000100;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110011100;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101110101;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101000;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100101;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100100;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111111;
SIGNAL_B = 14'b0001011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110001;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111011;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000110000;
SIGNAL_B = 14'b0001100000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111010;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101110;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101100;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110100000;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111001;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111001;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100001111;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101000;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100000011;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011100;
SIGNAL_B = 14'b0001100011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101001;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101000;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101001;
SIGNAL_B = 14'b0001100010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011010;
SIGNAL_B = 14'b0001100011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011001;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100110;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000111111;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111110;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111110;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000011000;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110001;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110111100;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100011;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110101111;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010101;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010101;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101000111;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101110;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010010;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010010;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010010;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011111001;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000101;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010010;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011111;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b0001100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001110110;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001000010;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001110110;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001000010;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100110;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000001;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110110011;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101001010;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101010111;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111011;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011100010;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011001000;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011101111;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101101;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011001000;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010010011;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010100001;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010001;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010001;
SIGNAL_B = 14'b0001101011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010001;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110110110;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000010;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101100111;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010111110;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011111110;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010010110;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111101;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001010110;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001010110;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000010100;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000010100;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000101110;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101100;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010011;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111000110;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101011;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101101010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000011;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100011100;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110100;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011101000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011001101;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001111111;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111111;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001111111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111111;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110010101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110000111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111011;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000110;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000010;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001010;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100101;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100100;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110000;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100110000;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001110001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010101;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b0001110000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001011110;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000010;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000001;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101011001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111101;
SIGNAL_B = 14'b0001110000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010110;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010101111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001000111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000100001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111010001;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111000100;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110110111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101101001;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011110100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100000001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110001;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111001000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111100010;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110100001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110100001;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111001000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101011111;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100000100;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011011101;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010101001;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010001110;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001011011;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011001;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110111110;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101110000;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101101111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100001;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010101100;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001011110;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101001;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110110;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101000;
SIGNAL_B = 14'b0001101011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110010;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110001;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100100100;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100011;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100011;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b0001101001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b0001101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001010011;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000110;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001010100;
SIGNAL_B = 14'b0001101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101101;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111101100;
SIGNAL_B = 14'b0001101001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111000100;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111000100;
SIGNAL_B = 14'b0001101000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000010;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110011101;
SIGNAL_B = 14'b0001101000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101000;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001110;
SIGNAL_B = 14'b0001100110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b0001100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001100100;
SIGNAL_B = 14'b0001100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001100100;
SIGNAL_B = 14'b0001100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100011;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000110000;
SIGNAL_B = 14'b0001100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001001010;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111011;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111011;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100010;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110101101;
SIGNAL_B = 14'b0001100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101011;
SIGNAL_B = 14'b0001100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100101010;
SIGNAL_B = 14'b0001100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100010000;
SIGNAL_B = 14'b0001100011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100010000;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011101;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011001111;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010101000;
SIGNAL_B = 14'b0001100010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001001101;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011001;
SIGNAL_B = 14'b0001100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001001101;
SIGNAL_B = 14'b0001100010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001001101;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110001;
SIGNAL_B = 14'b0001100001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110001;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111110010;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111001010;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101100010;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111011;
SIGNAL_B = 14'b0001100000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010100;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010010;
SIGNAL_B = 14'b0001011110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b0001011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011011111;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110110;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000011;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110111;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000010;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001110;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b0001011101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111101000;
SIGNAL_B = 14'b0001011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b0001011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000000;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000001;
SIGNAL_B = 14'b0001011011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001101;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b0001011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111101;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010110;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b0001011001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111100;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b0001010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101100;
SIGNAL_B = 14'b0001010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011110;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b0001010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101011;
SIGNAL_B = 14'b0001010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111110111;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010000;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b0001010011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100111;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b0001010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100110;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110001;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110001;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001101111;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010101;
SIGNAL_B = 14'b0001010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101110;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000001000;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000000111;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010011;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111100000;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b0001001011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b0001001001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b0001001011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011100;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000011;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b0001001001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b0001001000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b0001001000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001111;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b0001000111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011000;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110001;
SIGNAL_B = 14'b0001000110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011010;
SIGNAL_B = 14'b0001000110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b0001000110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b0001000101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b0001000101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010111;
SIGNAL_B = 14'b0001000011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111101;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b0001000010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b0001000010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b0001000000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010010;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b0000111111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b0000111111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b0000111101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b0000111101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b0000111100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b0000111001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b0000111000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110100;
SIGNAL_B = 14'b0000111001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b0000111000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b0000111001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000000;
SIGNAL_B = 14'b0000110111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b0000110110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110111001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110011;
SIGNAL_B = 14'b0000110011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b0000110011000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001101;
SIGNAL_B = 14'b0000110011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110001110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110010;
SIGNAL_B = 14'b0000101111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000110000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b0000110000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111100;
SIGNAL_B = 14'b0000110000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000101111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000101110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b0000101110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000101101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111011;
SIGNAL_B = 14'b0000101100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001000;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b0000101010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000101001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100001;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000101000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b0000100101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111000;
SIGNAL_B = 14'b0000100011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b0000100010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100001110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000110111;
SIGNAL_B = 14'b0000011110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000011110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000011000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b0000011000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000010110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000010101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000010110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110100111;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000010011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000010010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000010000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000010000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000001110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110000001;
SIGNAL_B = 14'b0000001101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110110;
SIGNAL_B = 14'b0000001100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001101100111;
SIGNAL_B = 14'b0000001011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000000111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000000100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110001110;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b1111111110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b1111111101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b1111111001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011101;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111111000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010001;
SIGNAL_B = 14'b1111110111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111110100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100001;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b1111110000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111101111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111101110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b1111101110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b1111101011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b1111101100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101111;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111101010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111101010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111100;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b1111101001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111101000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111100111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111100111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b1111100111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110011;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110111111;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b1111100001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001101;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001101;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011010;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111011111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b1111011110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b1111011110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000101000;
SIGNAL_B = 14'b1111011100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b1111011100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110100;
SIGNAL_B = 14'b1111011101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b1111011010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010010;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101001;
SIGNAL_B = 14'b1111011001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b1111011001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111010111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b1111010111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111001;
SIGNAL_B = 14'b1111010110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111010110110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010110110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b1111010101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010010;
SIGNAL_B = 14'b1111010011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100000;
SIGNAL_B = 14'b1111010011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000110;
SIGNAL_B = 14'b1111010010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000110;
SIGNAL_B = 14'b1111010001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b1111010001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110110000;
SIGNAL_B = 14'b1111001111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b1111001111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b1111001110011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100011;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011000;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b1111001011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001001110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b1111001001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b1111001001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001111;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101001;
SIGNAL_B = 14'b1111001001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011100;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b1111000101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101011110;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b1111000011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110011111;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b1111000011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010100;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010100;
SIGNAL_B = 14'b1111000010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b1111000001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010100;
SIGNAL_B = 14'b1111000001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001000;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010001010;
SIGNAL_B = 14'b1111000000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b1110111111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110010;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011001011;
SIGNAL_B = 14'b1110111111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100111;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110011;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101011011;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101000001;
SIGNAL_B = 14'b1110111011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110101;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b1110111010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b1110111001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101100;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b1110110111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b1110110111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111011;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000110;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b1110110111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b1110110110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011001000;
SIGNAL_B = 14'b1110110100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100011;
SIGNAL_B = 14'b1110110100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100011;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010111;
SIGNAL_B = 14'b1110110011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010110;
SIGNAL_B = 14'b1110110011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110000;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100101;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001110;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111101000;
SIGNAL_B = 14'b1110101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000001111;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b1110101111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011100;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101000;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000011;
SIGNAL_B = 14'b1110101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101010;
SIGNAL_B = 14'b1110101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001010000;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b1110101110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011010011;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000110;
SIGNAL_B = 14'b1110101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010011110;
SIGNAL_B = 14'b1110101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011011111;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011011111;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100000;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010011;
SIGNAL_B = 14'b1110101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110001001;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110001001;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110100011;
SIGNAL_B = 14'b1110101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111001010;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111100100;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011001;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b1110101010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011001;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001110;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000111111;
SIGNAL_B = 14'b1110101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010000001;
SIGNAL_B = 14'b1110100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010101000;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010000001;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010011011;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000100;
SIGNAL_B = 14'b1110100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100000011;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011101010;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100110111;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000101;
SIGNAL_B = 14'b1110100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b1110100101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010011;
SIGNAL_B = 14'b1110100011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b1110100100011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110010010;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b1110100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111011;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100011;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000110000;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000110000;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000101111;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001110000;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001100100;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010001011;
SIGNAL_B = 14'b1110100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011010;
SIGNAL_B = 14'b1110100001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010111111;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000001;
SIGNAL_B = 14'b1110100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011111111;
SIGNAL_B = 14'b1110100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011100110;
SIGNAL_B = 14'b1110011110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100101000;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001110;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b1110011111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b1110011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101011100;
SIGNAL_B = 14'b1110011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110011101;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110010000;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111000100;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010010;
SIGNAL_B = 14'b1110011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b1110011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101101;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b1110011100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101101;
SIGNAL_B = 14'b1110011100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b1110011100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111011;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010101111;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100011;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100100;
SIGNAL_B = 14'b1110011100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110010;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100010111;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100011000;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110001;
SIGNAL_B = 14'b1110011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b1110011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b1110011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110110100;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110101000;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101000;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000010;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111101000;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000010;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000000011;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000001111;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101001;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110110;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101010;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001111000;
SIGNAL_B = 14'b1110011000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100010;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101110;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100001;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101001000;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110010111;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101001000;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110100100;
SIGNAL_B = 14'b1110010111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001010;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110100100;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110011;
SIGNAL_B = 14'b1110010100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000011001;
SIGNAL_B = 14'b1110010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001101;
SIGNAL_B = 14'b1110010110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001110;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001110;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001011011;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010000010;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010110110;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011110111;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b1110010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101000110;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111001;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101110;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110111011;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111100010;
SIGNAL_B = 14'b1110010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111010101;
SIGNAL_B = 14'b1110010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000100011;
SIGNAL_B = 14'b1110010010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000001001;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000100011;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001010111;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001010111;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001011000;
SIGNAL_B = 14'b1110010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011110100;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b1110010010001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001110;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100011011;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011110100;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101001111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101000010;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101001111;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111000101;
SIGNAL_B = 14'b1110010001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110000100;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111000100;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111010010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000110;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000010011;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111010;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000010011;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000111010;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001100001;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001001;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100101;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100100101;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110011;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101110100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110000001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110001101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000111000;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001011110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001000100;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010101101;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111001;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010010010;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100001;
SIGNAL_B = 14'b1110001111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011010100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011010011;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111101;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010111;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100101;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001011;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011001;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001111;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000011;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100000101;
SIGNAL_B = 14'b1110001101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000111;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111010;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101100;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110010101;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b1110001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000001010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111111101;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011001;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001111111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010000000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b1110001100110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011001110;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011101000;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100011100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101010;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101010000;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101111000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110101100;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010011;
SIGNAL_B = 14'b1110001101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101101;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111100;
SIGNAL_B = 14'b1110001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001001000;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010111110;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011100101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011111111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101100111;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101101000;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101001;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111010000;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011101;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000101011;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000111000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001011111;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010100000;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011100010;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b1110001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101010111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101010111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001101;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110100101;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001101;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111110100;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000001;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000101000;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001001111;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001110110;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010000;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000110;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101000111;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101000111;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100101101;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101110;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b1110010010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001010;
SIGNAL_B = 14'b1110010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001011;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001011001;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110100;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100110;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b1110010010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011010;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110100;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011001111;
SIGNAL_B = 14'b1110010010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101000;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010001;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010001;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011110;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111001;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111000111;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000000111;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b1110010011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000111100;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010100100;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111110;
SIGNAL_B = 14'b1110010101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b1110010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011011001;
SIGNAL_B = 14'b1110010101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011100110;
SIGNAL_B = 14'b1110010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b1110010101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011001;
SIGNAL_B = 14'b1110010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101110101;
SIGNAL_B = 14'b1110010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000010;
SIGNAL_B = 14'b1110010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101000;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110001111;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101010;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011101;
SIGNAL_B = 14'b1110011000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011111;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000101100;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b1110011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010010100;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b1110011000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010000111;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100001;
SIGNAL_B = 14'b1110011001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b1110011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100100;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011101111;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100100;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011001;
SIGNAL_B = 14'b1110011011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b1110011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b1110011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111110101;
SIGNAL_B = 14'b1110011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000011100;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b1110011100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010000101;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011111;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011011111;
SIGNAL_B = 14'b1110011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000110;
SIGNAL_B = 14'b1110011100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111001;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010010;
SIGNAL_B = 14'b1110011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b1110011110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100000;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b1110011101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110000;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111101;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001010;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111001010;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111100101;
SIGNAL_B = 14'b1110100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011000;
SIGNAL_B = 14'b1110100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110011;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b1110100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001100111;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011011;
SIGNAL_B = 14'b1110100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b1110100011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110101;
SIGNAL_B = 14'b1110100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000100;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b1110100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b1110100101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110011111;
SIGNAL_B = 14'b1110100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101101;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101110;
SIGNAL_B = 14'b1110100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111010;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b1110100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111011;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b1110100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b1110100110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b1110100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100101;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100110;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010111111;
SIGNAL_B = 14'b1110101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001101;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b1110101001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110101;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b1110101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110101;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b1110101010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110111000;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b1110101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b1110101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b1110101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000110;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000011111;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b1110101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b1110101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b1110110000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111101;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100001011;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b1110110011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b1110110011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b1110110010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b1110110101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b1110110100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011100;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000010;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b1110111000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011100;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000001111;
SIGNAL_B = 14'b1110111001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b1110111001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011110;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b1110111011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010101;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101110;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100000111;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100001;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100000111;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010101;
SIGNAL_B = 14'b1110111110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b1110111111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100010;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1111000000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b1111000000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110010;
SIGNAL_B = 14'b1111000001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001011;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011001;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011001;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b1111000101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111000111110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011010;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111001001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b1111001010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000100;
SIGNAL_B = 14'b1111001001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101010;
SIGNAL_B = 14'b1111001001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000101;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000101;
SIGNAL_B = 14'b1111001100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101011;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111001111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111001111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011110;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000101;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b1111010010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000101;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111010110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b1111011000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111011000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111011000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111011001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111100;
SIGNAL_B = 14'b1111011010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111000111;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111011011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111101;
SIGNAL_B = 14'b1111011011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b1111011011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111011110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b1111011111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b1111100010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111100001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100001101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111100011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111100110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b1111100110010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111100111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110011000001;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110100;
SIGNAL_B = 14'b1111110010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110011000000;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110011000000;
SIGNAL_B = 14'b1111110110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b0000000000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b0000000001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b0000000010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b0000000001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b0000000011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001010;
SIGNAL_B = 14'b0000000101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000000110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000001000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000001000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111101;
SIGNAL_B = 14'b0000000110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001000;
SIGNAL_B = 14'b0000001010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000001101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111100;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000001110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000001111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000010001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010010;
SIGNAL_B = 14'b0000010010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000101;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010001;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000010101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000010101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101011;
SIGNAL_B = 14'b0000010111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000010111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b0000010111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010001;
SIGNAL_B = 14'b0000011001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110111;
SIGNAL_B = 14'b0000011001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011110;
SIGNAL_B = 14'b0000011010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011100011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010011100;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b0000011101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000011110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001000001;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b0000100001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100010000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100010100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000100001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111001100;
SIGNAL_B = 14'b0000100011100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111111;
SIGNAL_B = 14'b0000100100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110010111;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110010;
SIGNAL_B = 14'b0000100101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b0000100101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000100110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100110111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000100111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b0000101000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b0000101000111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100010100;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001000;
SIGNAL_B = 14'b0000101000111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b0000101001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101110;
SIGNAL_B = 14'b0000101010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b0000101010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b0000101010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b0000101011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010100;
SIGNAL_B = 14'b0000101100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b0000101101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b0000101100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b0000101110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101101;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010100000;
SIGNAL_B = 14'b0000101110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010000;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b0000101110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b0000101111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b0000110000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b0000101111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b0000110000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000101010;
SIGNAL_B = 14'b0000110000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000000011;
SIGNAL_B = 14'b0000110010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001111;
SIGNAL_B = 14'b0000110001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000001;
SIGNAL_B = 14'b0000110011011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110101000;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011011;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000001;
SIGNAL_B = 14'b0000110101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b0000110101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100010111;
SIGNAL_B = 14'b0000110110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001011;
SIGNAL_B = 14'b0000110110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010111;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110000;
SIGNAL_B = 14'b0000111000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b0000111010001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110001;
SIGNAL_B = 14'b0000111001001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b0000111001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010110000;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b0000111010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111100;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b0000111011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000101;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000110;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010010;
SIGNAL_B = 14'b0000111101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101100;
SIGNAL_B = 14'b0000111101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111111001;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111011110;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000101;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010001;
SIGNAL_B = 14'b0000111110110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b0000111111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000100;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0001000000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101110110;
SIGNAL_B = 14'b0001000000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b0001000000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011011;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100001110;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b0001000001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011100110;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b0001000010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011000000;
SIGNAL_B = 14'b0001000010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b0001000100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001110001;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001001010;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b0001000110011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b0001000110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101101;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101101;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101101;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b0001001010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b0001001001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b0001001001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100010001;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011101010;
SIGNAL_B = 14'b0001001010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011100;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011010000;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011011;
SIGNAL_B = 14'b0001001011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010011100;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000010;
SIGNAL_B = 14'b0001001011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000000;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000011000;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b0001001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111111;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110100100;
SIGNAL_B = 14'b0001001111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110111101;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001001;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110001010;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b0001010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b0001010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b0001010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b0001010001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111001;
SIGNAL_B = 14'b0001010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010011;
SIGNAL_B = 14'b0001010001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b0001010011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010011;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001110111;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010101011;
SIGNAL_B = 14'b0001010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001011101;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110101;
SIGNAL_B = 14'b0001010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110110;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111110101;
SIGNAL_B = 14'b0001010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000101000;
SIGNAL_B = 14'b0001010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000000;
SIGNAL_B = 14'b0001010110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110110011;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b0001010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001100;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001100;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101110010;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001011;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100100011;
SIGNAL_B = 14'b0001011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111100;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b0001011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011110000;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111100;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100001;
SIGNAL_B = 14'b0001011001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100001;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010010100;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101101;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001100000;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001000110;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b0001011011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111011110;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000010010;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111101011;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111000100;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111000100;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b0001011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000011;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110000010;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100100110;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101001110;
SIGNAL_B = 14'b0001011101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100100111;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001011;
SIGNAL_B = 14'b0001011111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011001100;
SIGNAL_B = 14'b0001011110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110001;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001001001;
SIGNAL_B = 14'b0001011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001111101;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111110;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b0001011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001100011;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000101111;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000010101;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111011;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101100;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110101101;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111000;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011111;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101000100;
SIGNAL_B = 14'b0001100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010010;
SIGNAL_B = 14'b0001100010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b0001100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100011100;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b0001100001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011001111;
SIGNAL_B = 14'b0001100011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011001111;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101001;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010110101;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011010;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010011010;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000111111;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000100101;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000011000;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000010111;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111110;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111110;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001010;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111010110;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010101;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b0001100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101100001;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b0001100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010010;
SIGNAL_B = 14'b0001100110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011101100;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011111001;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011111001;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010011;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010111000;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010010;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010010;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000101;
SIGNAL_B = 14'b0001100111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010001;
SIGNAL_B = 14'b0001100110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001110110;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001000010;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000100;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001011100;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000101000;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001011100;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000011011;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100110;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011001;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111110100;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110001011;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001100;
SIGNAL_B = 14'b0001101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101011000;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101011000;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100100011;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101001010;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b0001101011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011010100;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011001000;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010100001;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010000110;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111011;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b0001101011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001111001;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001011111;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000011;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b0001101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000011;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000100;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111010000;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000011;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111011101;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110110110;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101000000;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101000000;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011001011;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110001;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011110010;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011001010;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010111110;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001001000;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001001001;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000111011;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001001000;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000101111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101101;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110111001;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010011;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110010001;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101110111;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101001;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110101;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011101000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100011100;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100000010;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010011010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010100111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001100101;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010000000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001011;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000110001;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111100011;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110111011;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111001001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110000111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110001000;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101111011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010011;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101110;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100100000;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b0001110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011010001;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011111000;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000011;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010110111;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010011101;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000011;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011011;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110101;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000101000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011001;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111011001;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110010;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110011000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001011;
SIGNAL_B = 14'b0001110000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101001010;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100101111;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100010110;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011010100;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011010011;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010011111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010010011;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010000110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001110000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010000;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111110110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000010;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111011011;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100110;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100001100;
SIGNAL_B = 14'b0001101111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011100100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011010111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010101;
SIGNAL_B = 14'b0001110000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010100011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001111100;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001100001;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001010101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000101101;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111011111;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000110;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110101011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011101;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101110111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101000010;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011110100;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111111;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010111111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001111110;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110000;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110111011;
SIGNAL_B = 14'b0001101101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110100001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101111001;
SIGNAL_B = 14'b0001101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101111010;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010010;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101000110;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010011;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101111001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011011101;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010001111;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001101;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001001101;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001101;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111110010;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111001011;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110111110;
SIGNAL_B = 14'b0001101100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101111101;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101100011;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101101111;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100010;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011000110;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010101100;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010001;
SIGNAL_B = 14'b0001101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001000011;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000001111;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000010000;
SIGNAL_B = 14'b0001101011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111110101;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110001101;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110010;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101011001;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111111;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011100011;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100001011;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011110000;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010101111;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111010;
SIGNAL_B = 14'b0001101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111001;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101101;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000111010;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110010000;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110001111;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101001111;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000010;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b0001101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101000010;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001101;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110010;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011011001;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b0001100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b0001100110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001001001;
SIGNAL_B = 14'b0001100101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001001010;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000101111;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111111100;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b0001100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110101101;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111000111;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110101101;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101011111;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000101;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100101010;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000100;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100010000;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b0001100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b0001100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000011000;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b0001100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b0001100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111001010;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111001010;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111001010;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101111100;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101110000;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101001000;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101101;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111001;
SIGNAL_B = 14'b0001011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101101;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011111001;
SIGNAL_B = 14'b0001011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b0001011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000100;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010011110;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010011110;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101001;
SIGNAL_B = 14'b0001011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110110;
SIGNAL_B = 14'b0001011110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101000;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011011;
SIGNAL_B = 14'b0001011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000001;
SIGNAL_B = 14'b0001011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111101000;
SIGNAL_B = 14'b0001011100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111001100;
SIGNAL_B = 14'b0001011100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110100110;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111110;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111110;
SIGNAL_B = 14'b0001011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111110;
SIGNAL_B = 14'b0001011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b0001011010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b0001011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b0001010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b0001010111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b0001010111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001100000;
SIGNAL_B = 14'b0001010110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b0001010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000000100;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101011;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110111;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b0001010110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b0001010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101011011;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110100;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100111;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011010;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101000001;
SIGNAL_B = 14'b0001010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b0001010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b0001010010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011100101;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b0001010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b0001010010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110001;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010101;
SIGNAL_B = 14'b0001010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b0001010000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111011;
SIGNAL_B = 14'b0001001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001100011;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111011;
SIGNAL_B = 14'b0001010000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111011;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000010101;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111010;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111001;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101010;
SIGNAL_B = 14'b0001001100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b0001001011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b0001001100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b0001001011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110110;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100011101;
SIGNAL_B = 14'b0001001011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b0001001010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011001110;
SIGNAL_B = 14'b0001001001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b0001001001001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b0001000111111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b0001000111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001011001;
SIGNAL_B = 14'b0001000111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b0001000110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b0001000111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b0001000110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111110;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b0001000101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110001;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100100;
SIGNAL_B = 14'b0001000100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b0001000011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111100100;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110111100;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100011;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001010;
SIGNAL_B = 14'b0001000011101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100010;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000110;
SIGNAL_B = 14'b0001000000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101100001;
SIGNAL_B = 14'b0001000001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0001000000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111001;
SIGNAL_B = 14'b0000111111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100011111;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101011;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011101100;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b0000111110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010010;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000101;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b0000111101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b0000111100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011110;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000111001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000110101;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b0000111001001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b0000111000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000000;
SIGNAL_B = 14'b0000111000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b0000110110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110100;
SIGNAL_B = 14'b0000110110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b0000110101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b0000110100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b0000110011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000110011111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110001;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011001;
SIGNAL_B = 14'b0000110001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000110001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b0000110000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000110000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010110;
SIGNAL_B = 14'b0000101111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b0000101111110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b0000101110110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b0000101110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100001001;
SIGNAL_B = 14'b0000101101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111011;
SIGNAL_B = 14'b0000101101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b0000101101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111011;
SIGNAL_B = 14'b0000101011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b0000101011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b0000101010111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101001011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010101;
SIGNAL_B = 14'b0000101001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011101110;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b0000101001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000100111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b0000101000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000100111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111010;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b0000100111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100110001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b0000100100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b0000100101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000100011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b0000100010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000100001000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b0000100001100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b0000100000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000100000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000110111;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101010;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b0000011110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011101010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000011010111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b0000011010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b0000011010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000011001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000011000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000011000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000011000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000011001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000011001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000011;
SIGNAL_B = 14'b0000010111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000010100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000010011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b0000010010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000010001010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011100;
SIGNAL_B = 14'b0000010000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000010000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000010000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000001110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000001101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001100101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000001010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000001010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110011011;
SIGNAL_B = 14'b0000001001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000001000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000001000111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101000;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110101001;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000000100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b0000000011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111010000;
SIGNAL_B = 14'b0000000010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111001111;
SIGNAL_B = 14'b0000000001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001110110101;
SIGNAL_B = 14'b0000000010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011101;
SIGNAL_B = 14'b0000000001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b0000000001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b0000000001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000011;
SIGNAL_B = 14'b0000000000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b0000000000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b0000000000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111000010;
SIGNAL_B = 14'b1111111110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110110;
SIGNAL_B = 14'b1111111110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111011100;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111101001;
SIGNAL_B = 14'b1111111100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101010;
SIGNAL_B = 14'b1111111010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110001111110111;
SIGNAL_B = 14'b1111111011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010000;
SIGNAL_B = 14'b1111111001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000010001;
SIGNAL_B = 14'b1111111010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000101011;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111111010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111111000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000000100;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111111000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000110111;
SIGNAL_B = 14'b1111111000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000011110;
SIGNAL_B = 14'b1111110111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111110110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001010010;
SIGNAL_B = 14'b1111110101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010000111000;
SIGNAL_B = 14'b1111110110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001011111;
SIGNAL_B = 14'b1111110101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000101;
SIGNAL_B = 14'b1111110100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001000100;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001111001;
SIGNAL_B = 14'b1111110011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111110011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111110010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010000110;
SIGNAL_B = 14'b1111110010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010001101100;
SIGNAL_B = 14'b1111110001100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111110001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111110001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111110001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111100;
SIGNAL_B = 14'b1111110001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010100;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011001000;
SIGNAL_B = 14'b1111110000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010100000;
SIGNAL_B = 14'b1111101110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011010100;
SIGNAL_B = 14'b1111101111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010111011;
SIGNAL_B = 14'b1111101110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100001;
SIGNAL_B = 14'b1111101110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b1111101110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111101100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010010011;
SIGNAL_B = 14'b1111101100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011000111;
SIGNAL_B = 14'b1111101101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010010101101;
SIGNAL_B = 14'b1111101101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100010110;
SIGNAL_B = 14'b1111101100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111101011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011100010;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111101011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111101001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010011111011;
SIGNAL_B = 14'b1111101001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001001;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111101000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101001010;
SIGNAL_B = 14'b1111101001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111101001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101110000;
SIGNAL_B = 14'b1111101000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111101000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100100011;
SIGNAL_B = 14'b1111100111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100111101;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010100110000;
SIGNAL_B = 14'b1111100110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101010111;
SIGNAL_B = 14'b1111100110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100101110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101100100;
SIGNAL_B = 14'b1111100101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100100100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110001011;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100011110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110011000;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010101111110;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001100;
SIGNAL_B = 14'b1111100001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100110;
SIGNAL_B = 14'b1111100010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110110010;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111001101;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010110100101;
SIGNAL_B = 14'b1111100000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111000000;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111011001;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000001110;
SIGNAL_B = 14'b1111011110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111110011;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011101111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110010111100110;
SIGNAL_B = 14'b1111011110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000001;
SIGNAL_B = 14'b1111011110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000000000;
SIGNAL_B = 14'b1111011110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b1111011101001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011000011011;
SIGNAL_B = 14'b1111011101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000001;
SIGNAL_B = 14'b1111011011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b1111011100011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001001111;
SIGNAL_B = 14'b1111011011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010000;
SIGNAL_B = 14'b1111011010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001101001;
SIGNAL_B = 14'b1111011010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b1111011001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111011001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111011001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111011000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b1111011000100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111010111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b1111010111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011111;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b1111010110100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b1111010110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100000110;
SIGNAL_B = 14'b1111010101100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b1111010110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010011;
SIGNAL_B = 14'b1111010100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b1111010011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101101;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b1111010100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b1111010001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110001000;
SIGNAL_B = 14'b1111010011000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b1111010001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100010;
SIGNAL_B = 14'b1111010001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111010001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100011;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111001111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b1111001111001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b1111001111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110100011;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001111011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b1111001110111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111111101;
SIGNAL_B = 14'b1111001110101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000010111;
SIGNAL_B = 14'b1111001101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000011000;
SIGNAL_B = 14'b1111001101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b1111001100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b1111001100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b1111001100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000100101;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000111111;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010001101;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010000000;
SIGNAL_B = 14'b1111001011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001100;
SIGNAL_B = 14'b1111001011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110100;
SIGNAL_B = 14'b1111001010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b1111001010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b1111001001110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b1111001001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010100111;
SIGNAL_B = 14'b1111001010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011011;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b1111001000100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b1111001000010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b1111001000000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011110101;
SIGNAL_B = 14'b1111000110100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b1111000111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b1111000110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100000010;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101010;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000101000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101000100;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100101001;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101010001;
SIGNAL_B = 14'b1111000100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110010010;
SIGNAL_B = 14'b1111000101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b1111000011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b1111000100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b1111000100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101111000;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000111;
SIGNAL_B = 14'b1111000010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111010;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111111010;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000001000;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101110;
SIGNAL_B = 14'b1111000000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010011;
SIGNAL_B = 14'b1111000001111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000100010;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b1111000000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b1111000000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001110000;
SIGNAL_B = 14'b1111000000011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001001;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110001;
SIGNAL_B = 14'b1110111111101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010010111;
SIGNAL_B = 14'b1110111111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010001010;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b1110111110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b1110111101111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100001100;
SIGNAL_B = 14'b1110111101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011111111;
SIGNAL_B = 14'b1110111101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100011001;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111100000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b1110111011100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101110101;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110000010;
SIGNAL_B = 14'b1110111011010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110111;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110001111;
SIGNAL_B = 14'b1110111010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111010000;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111000011;
SIGNAL_B = 14'b1110111010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111111000;
SIGNAL_B = 14'b1110111001010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101010;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000010001;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111011101;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111001;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011110;
SIGNAL_B = 14'b1110111000100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011110;
SIGNAL_B = 14'b1110110110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b1110110110110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b1110110110010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b1110110110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010000111;
SIGNAL_B = 14'b1110110111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010101;
SIGNAL_B = 14'b1110110101011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010111100;
SIGNAL_B = 14'b1110110100101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011111100;
SIGNAL_B = 14'b1110110101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100011;
SIGNAL_B = 14'b1110110101001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b1110110110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100111110;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b1110110011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101100100;
SIGNAL_B = 14'b1110110011001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b1110110001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110010;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110001100;
SIGNAL_B = 14'b1110110011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111110;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000000;
SIGNAL_B = 14'b1110110001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110011001;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b1110110010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111000000;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000001;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011010;
SIGNAL_B = 14'b1110110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000000001;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110110;
SIGNAL_B = 14'b1110110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000110101;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b1110101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010000100;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110110;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010010001;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b1110101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100000110;
SIGNAL_B = 14'b1110101100010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010111000;
SIGNAL_B = 14'b1110101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011000101;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100010011;
SIGNAL_B = 14'b1110101101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101110;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101010101;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100001;
SIGNAL_B = 14'b1110101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101101;
SIGNAL_B = 14'b1110101010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b1110101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110110000;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111001010;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110111101;
SIGNAL_B = 14'b1110101001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001100;
SIGNAL_B = 14'b1110101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100101;
SIGNAL_B = 14'b1110101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001001101;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000110011;
SIGNAL_B = 14'b1110101001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b1110100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001001101;
SIGNAL_B = 14'b1110101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001110;
SIGNAL_B = 14'b1110100111100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010001110;
SIGNAL_B = 14'b1110100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b1110101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011100;
SIGNAL_B = 14'b1110100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011101;
SIGNAL_B = 14'b1110100111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011001111;
SIGNAL_B = 14'b1110100111110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011011011;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011101001;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b1110100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011101;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100110111;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101000100;
SIGNAL_B = 14'b1110100101101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000101;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111001;
SIGNAL_B = 14'b1110100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101010010;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b1110100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110111010;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111101110;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001000;
SIGNAL_B = 14'b1110100010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111010100;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b1110100010101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b1110100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000111101;
SIGNAL_B = 14'b1110100010011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010111;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001110001;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010110;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100110;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b1110100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010011001;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011001100;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100001110;
SIGNAL_B = 14'b1110100000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110100;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100011010;
SIGNAL_B = 14'b1110011111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110100;
SIGNAL_B = 14'b1110100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101001;
SIGNAL_B = 14'b1110100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101101000;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b1110011111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110010000;
SIGNAL_B = 14'b1110011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111101011;
SIGNAL_B = 14'b1110011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111111000;
SIGNAL_B = 14'b1110011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010010;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000110;
SIGNAL_B = 14'b1110011101110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000101100;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001010100;
SIGNAL_B = 14'b1110011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001101110;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b1110011101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111010;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111011;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001111011;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011010110;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010100011;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011111101;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010111100;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110001;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101001100;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110000000;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101011001;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101011001;
SIGNAL_B = 14'b1110011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101110011;
SIGNAL_B = 14'b1110011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100110;
SIGNAL_B = 14'b1110011011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100110;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110100111;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011011;
SIGNAL_B = 14'b1110011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b1110011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000011100;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110110;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110111;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000110111;
SIGNAL_B = 14'b1110011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001000011;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001101011;
SIGNAL_B = 14'b1110011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010000101;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b1110011001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011010011;
SIGNAL_B = 14'b1110011000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011101101;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100000111;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100001;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101110;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100001;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100111011;
SIGNAL_B = 14'b1110010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100010;
SIGNAL_B = 14'b1110010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101010110;
SIGNAL_B = 14'b1110010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101101111;
SIGNAL_B = 14'b1110010110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101111101;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110001;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110111110;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111011000;
SIGNAL_B = 14'b1110010110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111111111;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b1110010101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b1110010110111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110100;
SIGNAL_B = 14'b1110010101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000001100;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100111;
SIGNAL_B = 14'b1110010101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b1110010101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001011011;
SIGNAL_B = 14'b1110010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001110101;
SIGNAL_B = 14'b1110010101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010001111;
SIGNAL_B = 14'b1110010110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010101001;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010101001;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010110110;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011111;
SIGNAL_B = 14'b1110010100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011111000;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b1110010011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100111000;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b1110010100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101000101;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101111010;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101110;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110101101;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111100010;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111101111;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110111010;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111111100;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001001010;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001001010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110001;
SIGNAL_B = 14'b1110010010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000110000;
SIGNAL_B = 14'b1110010010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110010;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110010;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011011010;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011000000;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011100111;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001111;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100000010;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100101000;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101000010;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100101000;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100110101;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011100;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101101011100;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110011110;
SIGNAL_B = 14'b1110010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110000100;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111010010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111010001;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111000101;
SIGNAL_B = 14'b1110010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110000000110;
SIGNAL_B = 14'b1110010001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001010100;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001111011;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001111100;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001111100;
SIGNAL_B = 14'b1110010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b1110001111110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b1110010000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011001010;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100011000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011111110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001100;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100110;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101100110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101110100;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110001110;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110011011;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000010;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110100;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111101001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000110111;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000010001;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000110111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000011110;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000110111;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101100;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001111001;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101011;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001101011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010100000;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010010011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011100000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011111011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100011;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111101;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110001;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100110;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000001101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001001110;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001011011;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001101001;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000011;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000010;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b1110001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000011;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011011110;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101101101;
SIGNAL_B = 14'b1110001101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b1110001110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100001;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110010101;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b1110001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000001010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000010111;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111111101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001011;
SIGNAL_B = 14'b1110001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001011001;
SIGNAL_B = 14'b1110001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010001100;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010001101;
SIGNAL_B = 14'b1110001101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010110100;
SIGNAL_B = 14'b1110001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011100111;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110111;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b1110001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011111;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110000100;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110011111;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010011;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b1110001110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101101;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111001;
SIGNAL_B = 14'b1110001110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001001000;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b1110001111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110000;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010110001;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011001011;
SIGNAL_B = 14'b1110001110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011100101;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011011000;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100110011;
SIGNAL_B = 14'b1110001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011100101;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101001101;
SIGNAL_B = 14'b1110001111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011011;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011100;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111000011;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111010000;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110110101;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111110110;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000000011;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b1110010000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b1110001110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001010010;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010100000;
SIGNAL_B = 14'b1110001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011001000;
SIGNAL_B = 14'b1110001111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011100010;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b1110001111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100001001;
SIGNAL_B = 14'b1110001111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b1110010000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101010111;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110001;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b1110010000100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101111110;
SIGNAL_B = 14'b1110010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000000;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111101000;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001101;
SIGNAL_B = 14'b1110001111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111110100;
SIGNAL_B = 14'b1110010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010011101;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101010;
SIGNAL_B = 14'b1110010000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101010;
SIGNAL_B = 14'b1110010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010101011;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000101;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011111001;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100010011;
SIGNAL_B = 14'b1110010001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100101101;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101100001;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110001000;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110110000;
SIGNAL_B = 14'b1110010001001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010110;
SIGNAL_B = 14'b1110010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111001010;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111100100;
SIGNAL_B = 14'b1110010010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001011;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001010;
SIGNAL_B = 14'b1110010001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b1110010011011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b1110010011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b1110010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101001;
SIGNAL_B = 14'b1110010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b1110010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011011100;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b1110010100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100101010;
SIGNAL_B = 14'b1110010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011110;
SIGNAL_B = 14'b1110010011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101010001;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b1110010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110000110;
SIGNAL_B = 14'b1110010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110010010;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100000;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b1110010100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111101110;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111011;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000111100;
SIGNAL_B = 14'b1110010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000101111;
SIGNAL_B = 14'b1110010101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001010110;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b1110010101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b1110010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010010111;
SIGNAL_B = 14'b1110010101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011111111;
SIGNAL_B = 14'b1110010110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110001;
SIGNAL_B = 14'b1110010100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100001100;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011010;
SIGNAL_B = 14'b1110010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011010;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101011011;
SIGNAL_B = 14'b1110010111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101110101;
SIGNAL_B = 14'b1110010110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110110110;
SIGNAL_B = 14'b1110010111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110011100;
SIGNAL_B = 14'b1110011000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101010;
SIGNAL_B = 14'b1110010111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b1110010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b1110011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011111;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b1110010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011111;
SIGNAL_B = 14'b1110011000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001010011;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001101100;
SIGNAL_B = 14'b1110011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010100001;
SIGNAL_B = 14'b1110011001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010000111;
SIGNAL_B = 14'b1110011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b1110011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010010100;
SIGNAL_B = 14'b1110011001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011001001;
SIGNAL_B = 14'b1110011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101001100;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b1110011001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b1110011010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101100101;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b1110011010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b1110011011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b1110011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110011010;
SIGNAL_B = 14'b1110011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000010;
SIGNAL_B = 14'b1110011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b1110011011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000000001;
SIGNAL_B = 14'b1110011100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000101001;
SIGNAL_B = 14'b1110011011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001110;
SIGNAL_B = 14'b1110011100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b1110011100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000100;
SIGNAL_B = 14'b1110011100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001111000;
SIGNAL_B = 14'b1110011100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001110111;
SIGNAL_B = 14'b1110011101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011110;
SIGNAL_B = 14'b1110011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011000101;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011010010;
SIGNAL_B = 14'b1110011101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b1110011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111001;
SIGNAL_B = 14'b1110011110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111010;
SIGNAL_B = 14'b1110011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100000111;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100100001;
SIGNAL_B = 14'b1110011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b1110011111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111100;
SIGNAL_B = 14'b1110011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101111100;
SIGNAL_B = 14'b1110011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110010110;
SIGNAL_B = 14'b1110011111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110000;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110111101;
SIGNAL_B = 14'b1110011111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110111101;
SIGNAL_B = 14'b1110011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001011;
SIGNAL_B = 14'b1110100000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000001100;
SIGNAL_B = 14'b1110100001001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b1110100000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000111111;
SIGNAL_B = 14'b1110100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b1110100001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001011010;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b1110100010001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b1110100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010000001;
SIGNAL_B = 14'b1110100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110101;
SIGNAL_B = 14'b1110100010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011001111;
SIGNAL_B = 14'b1110100010111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b1110100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000011;
SIGNAL_B = 14'b1110100011001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011110111;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b1110100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b1110100100001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101101100;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101011111;
SIGNAL_B = 14'b1110100011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b1110100101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b1110100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110111011;
SIGNAL_B = 14'b1110100100111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010100;
SIGNAL_B = 14'b1110100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110101101;
SIGNAL_B = 14'b1110100110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b1110100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b1110100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111011;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000010110;
SIGNAL_B = 14'b1110100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b1110100111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100010;
SIGNAL_B = 14'b1110100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000110000;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b1110101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010011000;
SIGNAL_B = 14'b1110101000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110011;
SIGNAL_B = 14'b1110101001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010001011;
SIGNAL_B = 14'b1110101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100110;
SIGNAL_B = 14'b1110101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010100110;
SIGNAL_B = 14'b1110101001100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b1110101000010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000000;
SIGNAL_B = 14'b1110101000110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b1110101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b1110101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100101000;
SIGNAL_B = 14'b1110101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100110101;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b1110101010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b1110101011110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b1110101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110010000;
SIGNAL_B = 14'b1110101011100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110111000;
SIGNAL_B = 14'b1110101101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011110;
SIGNAL_B = 14'b1110101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111000101;
SIGNAL_B = 14'b1110101100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b1110101100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010010;
SIGNAL_B = 14'b1110101101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111010001;
SIGNAL_B = 14'b1110101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b1110101110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b1110101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000111010;
SIGNAL_B = 14'b1110101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110101111111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001100001;
SIGNAL_B = 14'b1110101111001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010001000;
SIGNAL_B = 14'b1110101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010110;
SIGNAL_B = 14'b1110110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010110000;
SIGNAL_B = 14'b1110110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010101111;
SIGNAL_B = 14'b1110110000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b1110110001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100011000;
SIGNAL_B = 14'b1110110001101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110001;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100100101;
SIGNAL_B = 14'b1110110010001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110010101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011000;
SIGNAL_B = 14'b1110110011101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100110001;
SIGNAL_B = 14'b1110110011111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b1110110011011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b1110110100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001011;
SIGNAL_B = 14'b1110110100001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b1110110100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011011;
SIGNAL_B = 14'b1110110100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101110011;
SIGNAL_B = 14'b1110110101110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110110100;
SIGNAL_B = 14'b1110110100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110101000;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001111;
SIGNAL_B = 14'b1110110101100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b1110110110010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b1110110111010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b1110110111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011100;
SIGNAL_B = 14'b1110110111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101000;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b1110111000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b1110111000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001011101;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b1110111001000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b1110111001110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010010010;
SIGNAL_B = 14'b1110111010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b1110111010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101101;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b1110111011110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010011111;
SIGNAL_B = 14'b1110111100100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b1110111101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011000110;
SIGNAL_B = 14'b1110111100111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111011;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010100;
SIGNAL_B = 14'b1110111100010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b1110111101101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100001;
SIGNAL_B = 14'b1110111101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100001;
SIGNAL_B = 14'b1110111101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100000111;
SIGNAL_B = 14'b1110111101001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111011;
SIGNAL_B = 14'b1110111101111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100101111;
SIGNAL_B = 14'b1110111110101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101010110;
SIGNAL_B = 14'b1110111110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1110111111001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1110111110011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101100011;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100101;
SIGNAL_B = 14'b1110111111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b1110111111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100101;
SIGNAL_B = 14'b1111000001101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b1111000010001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b1111000001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000010011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110001;
SIGNAL_B = 14'b1111000100000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b1111000010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b1111000011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b1111000011011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b1111000100010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110011;
SIGNAL_B = 14'b1111000100110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110011;
SIGNAL_B = 14'b1111000101010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b1111000111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b1111000111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001101000;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111000111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111000111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b1111001000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111001010000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b1111001001010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b1111001010000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b1111001001100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b1111001010010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b1111001100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b1111001100001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011010000;
SIGNAL_B = 14'b1111001100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b1111001101011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101011;
SIGNAL_B = 14'b1111001101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b1111001110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011111000;
SIGNAL_B = 14'b1111001110001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010001;
SIGNAL_B = 14'b1111001110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111001110001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b1111001110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b1111010000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b1111010000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010001011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010000011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100101100;
SIGNAL_B = 14'b1111010001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b1111010010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b1111010010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b1111010010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b1111010100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010101000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b1111010100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b1111010110010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b1111010110110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010111000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b1111010111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111010111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100010;
SIGNAL_B = 14'b1111011000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011001010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111100;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111100;
SIGNAL_B = 14'b1111011000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111110000;
SIGNAL_B = 14'b1111011010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101110;
SIGNAL_B = 14'b1111011010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b1111011011011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111101;
SIGNAL_B = 14'b1111011011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b1111011011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b1111011100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b1111011100001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b1111011110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010110;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b1111011111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b1111011111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111011111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b1111100000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111100011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100011010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111100100000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001100;
SIGNAL_B = 14'b1111100011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111100011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111100100010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111100100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111100101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111100110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111100111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111100111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111100111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111101000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001010;
SIGNAL_B = 14'b1111101000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111101010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101001111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111101010101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111101010101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010110100;
SIGNAL_B = 14'b1111101010011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111101011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101100111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111101011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101110001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111101111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111101111001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111101110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111101111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110001;
SIGNAL_B = 14'b1111110000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110001110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010100110;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111110100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111110101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111110101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110101010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111110111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111110111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111110110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001110010;
SIGNAL_B = 14'b1111111001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111001111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100101;
SIGNAL_B = 14'b1111111011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010011001;
SIGNAL_B = 14'b1111111100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110010001100;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001100100;
SIGNAL_B = 14'b1111111101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b1111111100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b1111111101101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001111111;
SIGNAL_B = 14'b1111111101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b1111111110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001010111;
SIGNAL_B = 14'b1111111101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b1111111110111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b1111111111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111101;
SIGNAL_B = 14'b1111111111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b1111111111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001001011;
SIGNAL_B = 14'b0000000001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b0000000001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111101;
SIGNAL_B = 14'b0000000001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100011;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110001011000;
SIGNAL_B = 14'b0000000010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000000010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000100100;
SIGNAL_B = 14'b0000000011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000111110;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111101111;
SIGNAL_B = 14'b0000000100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110000;
SIGNAL_B = 14'b0000000100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000000101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000001001;
SIGNAL_B = 14'b0000000101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010110;
SIGNAL_B = 14'b0000000110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000110001;
SIGNAL_B = 14'b0000000111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001110000010111;
SIGNAL_B = 14'b0000001000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100011;
SIGNAL_B = 14'b0000001000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000001001111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001001011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111010101;
SIGNAL_B = 14'b0000001001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001010101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111001001;
SIGNAL_B = 14'b0000001100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111111100;
SIGNAL_B = 14'b0000001011101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110101111;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110111011;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001100001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001100011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101111100010;
SIGNAL_B = 14'b0000001101001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110010100;
SIGNAL_B = 14'b0000001101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110100001;
SIGNAL_B = 14'b0000001111010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000001111000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000001110110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000001111000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101100;
SIGNAL_B = 14'b0000010000000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101110000111;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010001000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101111010;
SIGNAL_B = 14'b0000010001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101101101;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101100000;
SIGNAL_B = 14'b0000010001110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101000110;
SIGNAL_B = 14'b0000010010010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101101010011;
SIGNAL_B = 14'b0000010010110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111000;
SIGNAL_B = 14'b0000010011000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010100000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100010010;
SIGNAL_B = 14'b0000010101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000010101000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100011111;
SIGNAL_B = 14'b0000010101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100111001;
SIGNAL_B = 14'b0000010101010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011110111;
SIGNAL_B = 14'b0000010110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011101010;
SIGNAL_B = 14'b0000010110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000010110001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101100000100;
SIGNAL_B = 14'b0000010111011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011110;
SIGNAL_B = 14'b0000010111101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011000011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011011101;
SIGNAL_B = 14'b0000011000101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110111;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011000111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000011;
SIGNAL_B = 14'b0000011001011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000100;
SIGNAL_B = 14'b0000011001001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101011000100;
SIGNAL_B = 14'b0000011001101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010110110;
SIGNAL_B = 14'b0000011001111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101010;
SIGNAL_B = 14'b0000011010011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011011001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011010011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011011111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011100011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010001111;
SIGNAL_B = 14'b0000011100011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010101001;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011100111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101010000010;
SIGNAL_B = 14'b0000011101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001110101;
SIGNAL_B = 14'b0000011110000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b0000011110100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001001110;
SIGNAL_B = 14'b0000011110100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100111;
SIGNAL_B = 14'b0000011111010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101001011011;
SIGNAL_B = 14'b0000011111100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000011111110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000110100;
SIGNAL_B = 14'b0000100000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000100000010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000100110;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000001101;
SIGNAL_B = 14'b0000100000110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100000110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001101000011010;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111111111;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100010100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100010010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111110010;
SIGNAL_B = 14'b0000100011010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110111110;
SIGNAL_B = 14'b0000100011110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111011000;
SIGNAL_B = 14'b0000100100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100111100101;
SIGNAL_B = 14'b0000100100011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110001010;
SIGNAL_B = 14'b0000100100110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b0000100101011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111100;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110110010;
SIGNAL_B = 14'b0000100101101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100110100100;
SIGNAL_B = 14'b0000100110101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101111101;
SIGNAL_B = 14'b0000100110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000100111011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000100110111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101110000;
SIGNAL_B = 14'b0000100111111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b0000101000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100010;
SIGNAL_B = 14'b0000101001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100101001001;
SIGNAL_B = 14'b0000101000001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100111100;
SIGNAL_B = 14'b0000101001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b0000101001111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101000101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b0000101010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b0000101010101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100100001;
SIGNAL_B = 14'b0000101001001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011111010;
SIGNAL_B = 14'b0000101010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101110;
SIGNAL_B = 14'b0000101011011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100100001000;
SIGNAL_B = 14'b0000101011111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101011101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011100000;
SIGNAL_B = 14'b0000101100110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011101101;
SIGNAL_B = 14'b0000101100100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010101100;
SIGNAL_B = 14'b0000101100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100011010011;
SIGNAL_B = 14'b0000101101110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010000101;
SIGNAL_B = 14'b0000101110000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100010111001;
SIGNAL_B = 14'b0000101110000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000110111;
SIGNAL_B = 14'b0000101101110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b0000101101100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001101011;
SIGNAL_B = 14'b0000101111010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001111000;
SIGNAL_B = 14'b0000101111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b0000110000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000101111100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001000100;
SIGNAL_B = 14'b0000110000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100001010001;
SIGNAL_B = 14'b0000110000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111110101;
SIGNAL_B = 14'b0000110000110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111101001;
SIGNAL_B = 14'b0000110000000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011100;
SIGNAL_B = 14'b0000110001000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000010000;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001100000011101;
SIGNAL_B = 14'b0000110010010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111011011;
SIGNAL_B = 14'b0000110011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111001110;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b0000110010100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011111000010;
SIGNAL_B = 14'b0000110010110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110011101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110100111;
SIGNAL_B = 14'b0000110010110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110101000;
SIGNAL_B = 14'b0000110011000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110011010;
SIGNAL_B = 14'b0000110100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b0000110100101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101011001;
SIGNAL_B = 14'b0000110101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110000000;
SIGNAL_B = 14'b0000110101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011110001101;
SIGNAL_B = 14'b0000110100111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001100;
SIGNAL_B = 14'b0000110101001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100111111;
SIGNAL_B = 14'b0000110101111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b0000110110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101100110;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011101001011;
SIGNAL_B = 14'b0000110111111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011100010111;
SIGNAL_B = 14'b0000110111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000111000001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011110000;
SIGNAL_B = 14'b0000110111101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011100011;
SIGNAL_B = 14'b0000111000101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011111110;
SIGNAL_B = 14'b0000111000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011010110;
SIGNAL_B = 14'b0000110111111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011011001001;
SIGNAL_B = 14'b0000111010001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010101;
SIGNAL_B = 14'b0000111001101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010111101;
SIGNAL_B = 14'b0000111010101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010010110;
SIGNAL_B = 14'b0000111001011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001111011;
SIGNAL_B = 14'b0000111010011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011010100010;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b0000111010111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001101110;
SIGNAL_B = 14'b0000111011010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000111;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111100000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000101101;
SIGNAL_B = 14'b0000111011001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011001000110;
SIGNAL_B = 14'b0000111100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000100000;
SIGNAL_B = 14'b0000111101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000010011;
SIGNAL_B = 14'b0000111100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001011000000110;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110101010;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b0000111111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010111101011;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110111000;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110110111;
SIGNAL_B = 14'b0000111111000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b0000111111100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110011101;
SIGNAL_B = 14'b0000111111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101001111;
SIGNAL_B = 14'b0000111111110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101101001;
SIGNAL_B = 14'b0001000000110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010110000011;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101011100;
SIGNAL_B = 14'b0001000000010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010101000010;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100011011;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100000001;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010100001110;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011001100;
SIGNAL_B = 14'b0001000010011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011110100;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b0001000100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010011011001;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110011;
SIGNAL_B = 14'b0001000011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010010110010;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001111110;
SIGNAL_B = 14'b0001000100101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001010111;
SIGNAL_B = 14'b0001000101101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010001100100;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100010;
SIGNAL_B = 14'b0001000100111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000111101;
SIGNAL_B = 14'b0001000101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000001001;
SIGNAL_B = 14'b0001000101101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001010000100011;
SIGNAL_B = 14'b0001000101111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b0001000110011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111101111;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111111100;
SIGNAL_B = 14'b0001000110101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111010101;
SIGNAL_B = 14'b0001000111011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111100001;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001111000111;
SIGNAL_B = 14'b0001000111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010011;
SIGNAL_B = 14'b0001001000001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110100000;
SIGNAL_B = 14'b0001000111011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101111001;
SIGNAL_B = 14'b0001001001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110010011;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000111;
SIGNAL_B = 14'b0001001000011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101010010;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001101000101;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001110000110;
SIGNAL_B = 14'b0001001010010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b0001001001111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100101011;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100011110;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001100000100;
SIGNAL_B = 14'b0001001010100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011011100;
SIGNAL_B = 14'b0001001010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010110101;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b0001001011100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001011000010;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b0001001011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010101000;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001110100;
SIGNAL_B = 14'b0001001011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001010001111;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001001101;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b0001001101000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001001000000;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000110011;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001001000100101;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111111;
SIGNAL_B = 14'b0001001110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111110010;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110111101;
SIGNAL_B = 14'b0001010000000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111010111;
SIGNAL_B = 14'b0001010000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000111111111;
SIGNAL_B = 14'b0001010000010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000110110000;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101001000;
SIGNAL_B = 14'b0001001111100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b0001010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101010101;
SIGNAL_B = 14'b0001010000110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000101100010;
SIGNAL_B = 14'b0001010001000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b0001010001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100101110;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100000110;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111010;
SIGNAL_B = 14'b0001010001010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011100000;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011111010;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000100010100;
SIGNAL_B = 14'b0001010010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011101;
SIGNAL_B = 14'b0001010010111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000011101101;
SIGNAL_B = 14'b0001010011101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010111000;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010011110;
SIGNAL_B = 14'b0001010100001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010010001;
SIGNAL_B = 14'b0001010100011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000010101011;
SIGNAL_B = 14'b0001010011111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001101010;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b0001010100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001010000;
SIGNAL_B = 14'b0001010100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b0001010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110110;
SIGNAL_B = 14'b0001010101001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000110110;
SIGNAL_B = 14'b0001010101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000001000011;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0001000000001111;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111101000;
SIGNAL_B = 14'b0001010101111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111011011;
SIGNAL_B = 14'b0001010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111100111;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b0001010110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110100110;
SIGNAL_B = 14'b0001011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111111000001;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111110001101;
SIGNAL_B = 14'b0001010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101011000;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111101111111;
SIGNAL_B = 14'b0001011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100111110;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100110001;
SIGNAL_B = 14'b0001010111101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100001010;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011010110;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111011111101;
SIGNAL_B = 14'b0001011000011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111100001001;
SIGNAL_B = 14'b0001011000110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010111011;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010010100;
SIGNAL_B = 14'b0001011001110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111011;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111010010100;
SIGNAL_B = 14'b0001011011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111010;
SIGNAL_B = 14'b0001011010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001111011;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111001010011;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b0001011011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000011111;
SIGNAL_B = 14'b0001011010110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000101100;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000111001;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000111000000101;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111111000;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111010001;
SIGNAL_B = 14'b0001011011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110111000011;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110101001;
SIGNAL_B = 14'b0001011011100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101110101;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110011100;
SIGNAL_B = 14'b0001011101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110110010000;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101101001;
SIGNAL_B = 14'b0001011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110101000001;
SIGNAL_B = 14'b0001011101100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100011010;
SIGNAL_B = 14'b0001011110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100001101;
SIGNAL_B = 14'b0001011110000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110100000000;
SIGNAL_B = 14'b0001011110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011110011;
SIGNAL_B = 14'b0001011110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011011000;
SIGNAL_B = 14'b0001011110010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110011011001;
SIGNAL_B = 14'b0001011110110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010111111;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010110001;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110010001010;
SIGNAL_B = 14'b0001011111100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110000;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110001110001;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000100010;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000111100;
SIGNAL_B = 14'b0001100000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000111100;
SIGNAL_B = 14'b0001100000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000001000;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000110000000111;
SIGNAL_B = 14'b0001100000111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111111010;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111100001;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111010100;
SIGNAL_B = 14'b0001100000001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110111001;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101111000111;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101110011111;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011110;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101111000;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101011;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101101100;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101101011110;
SIGNAL_B = 14'b0001100010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100110111;
SIGNAL_B = 14'b0001100001101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110110;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101100010000;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011110101;
SIGNAL_B = 14'b0001100011011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011101000;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011001111;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101011000010;
SIGNAL_B = 14'b0001100010011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010100111;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101010001101;
SIGNAL_B = 14'b0001100011001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110011;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001110100;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001100111;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000111111;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000110010;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101001001100;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000101000001010;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111110001;
SIGNAL_B = 14'b0001100100111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111111110;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100111100100;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110010101;
SIGNAL_B = 14'b0001100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111011;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101110;
SIGNAL_B = 14'b0001100101011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100110100010;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101111100;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100111010;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101010100;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100101101111;
SIGNAL_B = 14'b0001100110001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100101101;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000101;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100100000110;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011011111;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011010010;
SIGNAL_B = 14'b0001100110011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100011000100;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010010000;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010111000;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010011110;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100010000011;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001101001;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100001011100;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000001110;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000110101;
SIGNAL_B = 14'b0001100111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111011010;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000001;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000100000000000;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111001101;
SIGNAL_B = 14'b0001101000110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011111100111;
SIGNAL_B = 14'b0001101000100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110100101;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101111111;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110011000;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011110100110;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101110010;
SIGNAL_B = 14'b0001101010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011101011000;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100110000;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100111101;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011111100;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100111101;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011000111;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011100010110;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010101110;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011001000;
SIGNAL_B = 14'b0001101010100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011100001;
SIGNAL_B = 14'b0001101011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011010111010;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011011101111;
SIGNAL_B = 14'b0001101010000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001011111;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001011111;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001000101;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011001101100;
SIGNAL_B = 14'b0001101010110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010001;
SIGNAL_B = 14'b0001101010010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000011110;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000011000010001;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111101010;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110101000;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110001110;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010111010000;
SIGNAL_B = 14'b0001101011010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110011011;
SIGNAL_B = 14'b0001101011010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101100111;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101110100;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010110000001;
SIGNAL_B = 14'b0001101100100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010101011010;
SIGNAL_B = 14'b0001101011110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100001100;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100100110;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010100011001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010111110;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011010111;
SIGNAL_B = 14'b0001101101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010011001010;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001001;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010100100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010010001001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001101111;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001111100;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010001010101;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111100000;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000010000100001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010100;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111101101;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111010011;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001111111010;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110010001;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101000011;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101101011;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001110010001;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001101011101;
SIGNAL_B = 14'b0001101101100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100011100;
SIGNAL_B = 14'b0001101110110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100101001;
SIGNAL_B = 14'b0001101101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100001111;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001100110110;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011110101;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011011011;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001011000001;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001111111;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001111111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001010000000;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110010;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001110010;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000111110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000100101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001001001011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111111101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000001000001010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111111101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110111011;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000111010110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110111100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110010101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110100010;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000110101110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101100000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000110;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101000111;
SIGNAL_B = 14'b0001110000011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000101010100;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101011;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100101100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100011111;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100111001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000100010010;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011011110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011000100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000011101011;
SIGNAL_B = 14'b0001101111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010101010;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000010;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010000010;
SIGNAL_B = 14'b0001110000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000010010000;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110101;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001110101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000001000001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000110100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000011001;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000100111;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111110010;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111100110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b0000000000000000;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111111001011;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110111111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110110010;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110001011;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111110100100;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110001;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101010111;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101100011;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111101110000;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100100010;
SIGNAL_B = 14'b0001110000001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100111100;
SIGNAL_B = 14'b0001110000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001110000101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111100001000;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011101110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011000111;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111011010100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010111010;
SIGNAL_B = 14'b0001110000101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111010100000;
SIGNAL_B = 14'b0001101111101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000110111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001000100;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010010;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111001010001;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000000011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111111000101011;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111001111;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110101000;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110111000001;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110110101;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110110001110;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110100110010;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110101001100;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110011110001;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010101111;
SIGNAL_B = 14'b0001110000011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010111101;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001001;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010001000;
SIGNAL_B = 14'b0001101111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010110000;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110010010110;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111110001101111;
SIGNAL_B = 14'b0001110000001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111111001;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111101100;
SIGNAL_B = 14'b0001101111111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111000101;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101111010010;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110111000;
SIGNAL_B = 14'b0001101110101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110010001;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110000100;
SIGNAL_B = 14'b0001101111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101110000100;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100101000;
SIGNAL_B = 14'b0001101111011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101100001110;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b0001101110000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010011001;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101011001100;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010110011;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101010100110;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001110001;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101001100101;
SIGNAL_B = 14'b0001101111011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000111101;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111101000010110;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100111101111;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110010100;
SIGNAL_B = 14'b0001101110011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b0001101110111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101101101;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b0001101111001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100101010011;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100110000111;
SIGNAL_B = 14'b0001101110010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100011110;
SIGNAL_B = 14'b0001101110000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100101011;
SIGNAL_B = 14'b0001101110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100100010001;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011010000;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100010011100;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011101010;
SIGNAL_B = 14'b0001101101010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100011000011;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001100111;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001101000;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b0001101101100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000100110;
SIGNAL_B = 14'b0001101101110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100001000000;
SIGNAL_B = 14'b0001101100010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111100000110011;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011111100101;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110110000;
SIGNAL_B = 14'b0001101100110110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110001001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011110010111;
SIGNAL_B = 14'b0001101101000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011101010110;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100100001;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100101110;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011100010100;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011111010;
SIGNAL_B = 14'b0001101100100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011011010011;
SIGNAL_B = 14'b0001101100000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b0001101100110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010111001;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010010010;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011010011110;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001010000;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011001000011;
SIGNAL_B = 14'b0001101100010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111110110;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111011000101001;
SIGNAL_B = 14'b0001101011000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111011010;
SIGNAL_B = 14'b0001101011100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111001110;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010111000001;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110011010;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b0001101100000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b0001101010100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010110001101;
SIGNAL_B = 14'b0001101010110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010101100110;
SIGNAL_B = 14'b0001101001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100110001;
SIGNAL_B = 14'b0001101010010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010100111110;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011110000;
SIGNAL_B = 14'b0001101011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010100010;
SIGNAL_B = 14'b0001101001010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010010010101;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010011001001;
SIGNAL_B = 14'b0001101001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001100001;
SIGNAL_B = 14'b0001101001100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010001000111;
SIGNAL_B = 14'b0001101000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000010010;
SIGNAL_B = 14'b0001101001110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000011111;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000000101;
SIGNAL_B = 14'b0001101001010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111010000011111;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111111000;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111010001;
SIGNAL_B = 14'b0001100111110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001111011110;
SIGNAL_B = 14'b0001101000100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110110111;
SIGNAL_B = 14'b0001101001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110011101;
SIGNAL_B = 14'b0001100111100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001101110110;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110000011;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001110011101;
SIGNAL_B = 14'b0001101000010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100110101;
SIGNAL_B = 14'b0001100110101111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100100111;
SIGNAL_B = 14'b0001101000000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001100000000;
SIGNAL_B = 14'b0001100110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011100110;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001011110011;
SIGNAL_B = 14'b0001100110011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010100101;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001010110010;
SIGNAL_B = 14'b0001100111001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001111110;
SIGNAL_B = 14'b0001100101101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001110001;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001001001;
SIGNAL_B = 14'b0001100110001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001100100;
SIGNAL_B = 14'b0001100101111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001001010110;
SIGNAL_B = 14'b0001100101111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000100010;
SIGNAL_B = 14'b0001100101001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000010101;
SIGNAL_B = 14'b0001100100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b0001100101011110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111001000001001;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000111100001;
SIGNAL_B = 14'b0001100100001100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101111001;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110100000;
SIGNAL_B = 14'b0001100011111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000101101100;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000110000101;
SIGNAL_B = 14'b0001100100111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b0001100100101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100111000;
SIGNAL_B = 14'b0001100100011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000100011110;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011010000;
SIGNAL_B = 14'b0001100011011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011101010;
SIGNAL_B = 14'b0001100011101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000011000010;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000010110101;
SIGNAL_B = 14'b0001100010111011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001110100;
SIGNAL_B = 14'b0001100001111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b0001100010101010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001100111;
SIGNAL_B = 14'b0001100010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001011010;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000100110;
SIGNAL_B = 14'b0001100010001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000001000000;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111010111;
SIGNAL_B = 14'b0001100001011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1111000000001011;
SIGNAL_B = 14'b0001100001101001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111111110;
SIGNAL_B = 14'b0001100000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111001010;
SIGNAL_B = 14'b0001100000011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110001001;
SIGNAL_B = 14'b0001100001001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111111011000;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b0001100000101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111110010110;
SIGNAL_B = 14'b0001011111111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111101101111;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100111011;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101101;
SIGNAL_B = 14'b0001011111101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100101101;
SIGNAL_B = 14'b0001011111110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011100000;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111100100000;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011101100;
SIGNAL_B = 14'b0001011110100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111011100000;
SIGNAL_B = 14'b0001011111000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010011110;
SIGNAL_B = 14'b0001011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111010101011;
SIGNAL_B = 14'b0001011111010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001110110;
SIGNAL_B = 14'b0001011110100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001101010;
SIGNAL_B = 14'b0001011101110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001000011;
SIGNAL_B = 14'b0001011110010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111001001111;
SIGNAL_B = 14'b0001011111000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b0001011101000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000101001;
SIGNAL_B = 14'b0001011100100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110111000011011;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110101;
SIGNAL_B = 14'b0001011100000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111100111;
SIGNAL_B = 14'b0001011101000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111011011;
SIGNAL_B = 14'b0001011101010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110111110100;
SIGNAL_B = 14'b0001011011010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110110011;
SIGNAL_B = 14'b0001011011110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110011001;
SIGNAL_B = 14'b0001011011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110110011001;
SIGNAL_B = 14'b0001011011000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101110001;
SIGNAL_B = 14'b0001011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101111111;
SIGNAL_B = 14'b0001011011000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110101001011;
SIGNAL_B = 14'b0001011010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100110001;
SIGNAL_B = 14'b0001011010000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100100100;
SIGNAL_B = 14'b0001011001100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100010110;
SIGNAL_B = 14'b0001011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011101111;
SIGNAL_B = 14'b0001011010010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011100010;
SIGNAL_B = 14'b0001011010000010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110100001001;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110011010110;
SIGNAL_B = 14'b0001011001010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010100001;
SIGNAL_B = 14'b0001010111011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010101110;
SIGNAL_B = 14'b0001011001000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110010010100;
SIGNAL_B = 14'b0001011001000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001111010;
SIGNAL_B = 14'b0001011000100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001101101;
SIGNAL_B = 14'b0001011000010000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001000110;
SIGNAL_B = 14'b0001011000001111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110001010011;
SIGNAL_B = 14'b0001010111111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000101011;
SIGNAL_B = 14'b0001010111101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000111000;
SIGNAL_B = 14'b0001010110101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110110000011111;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111111000;
SIGNAL_B = 14'b0001010101101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b0001010110001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101011;
SIGNAL_B = 14'b0001010101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101111101011;
SIGNAL_B = 14'b0001010101001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110110110;
SIGNAL_B = 14'b0001010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110101001;
SIGNAL_B = 14'b0001010110011101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101101000;
SIGNAL_B = 14'b0001010101011100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101110011100;
SIGNAL_B = 14'b0001010100101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101011011;
SIGNAL_B = 14'b0001010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b0001010011101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101011011;
SIGNAL_B = 14'b0001010100001011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101101001110;
SIGNAL_B = 14'b0001010011111010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100100110;
SIGNAL_B = 14'b0001010010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101100110100;
SIGNAL_B = 14'b0001010011001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110011;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b0001010011001010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011110010;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010111110;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101011011000;
SIGNAL_B = 14'b0001010001011000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010110010;
SIGNAL_B = 14'b0001010010001001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101010100100;
SIGNAL_B = 14'b0001010001101000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001111101;
SIGNAL_B = 14'b0001010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b0001010000010111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000111100;
SIGNAL_B = 14'b0001010000111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001010110;
SIGNAL_B = 14'b0001001111100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101000101111;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110101001001000;
SIGNAL_B = 14'b0001001110110101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101101;
SIGNAL_B = 14'b0001001111000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111101110;
SIGNAL_B = 14'b0001001111010110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111010011;
SIGNAL_B = 14'b0001001110000100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100111000110;
SIGNAL_B = 14'b0001001110100101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110111010;
SIGNAL_B = 14'b0001001101110100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110101100;
SIGNAL_B = 14'b0001001101100100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b0001001101010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b0001001100010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001100110011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001100100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b0001001011000001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100101101011;
SIGNAL_B = 14'b0001001011100010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100110000101;
SIGNAL_B = 14'b0001001011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b0001001011110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100110111;
SIGNAL_B = 14'b0001001010110001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b0001001011010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011100;
SIGNAL_B = 14'b0001001010110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b0001001001011111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100100010000;
SIGNAL_B = 14'b0001001010000000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011011100;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011101000;
SIGNAL_B = 14'b0001001000111110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b0001001010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110101;
SIGNAL_B = 14'b0001001000111111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100011000001;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010011010;
SIGNAL_B = 14'b0001001000101110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100010110100;
SIGNAL_B = 14'b0001001000001110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b0001000110111101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001100110;
SIGNAL_B = 14'b0001000111001101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001001011;
SIGNAL_B = 14'b0001000110111100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b0001000111101101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001110011;
SIGNAL_B = 14'b0001000101011010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b0001000110101100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000110010;
SIGNAL_B = 14'b0001000101011011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100000001011;
SIGNAL_B = 14'b0001000100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110100001000000;
SIGNAL_B = 14'b0001000100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111010110;
SIGNAL_B = 14'b0001000100101011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111110000;
SIGNAL_B = 14'b0001000011111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b0001000010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b0001000100011001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011111001001;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110101111;
SIGNAL_B = 14'b0001000010111001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b0001000010000111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011110010101;
SIGNAL_B = 14'b0001000010111000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101111011;
SIGNAL_B = 14'b0001000011001000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101010100;
SIGNAL_B = 14'b0001000001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b0001000001000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101101110;
SIGNAL_B = 14'b0001000001100111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011101000111;
SIGNAL_B = 14'b0001000001110111;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0001000001100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100111010;
SIGNAL_B = 14'b0001000000100110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010010;
SIGNAL_B = 14'b0001000000000101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011111000;
SIGNAL_B = 14'b0001000000000110;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100101100;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100100000;
SIGNAL_B = 14'b0000111111010100;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100011111;
SIGNAL_B = 14'b0000111111010101;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011100010010;
SIGNAL_B = 14'b0000111110010011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010001;
SIGNAL_B = 14'b0000111110100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011010010;
SIGNAL_B = 14'b0000111101100011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011000100;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010010001;
SIGNAL_B = 14'b0000111110000011;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111101010010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010101010;
SIGNAL_B = 14'b0000111100100001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010110111;
SIGNAL_B = 14'b0000111100110010;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011011011110;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010011101;
SIGNAL_B = 14'b0000111011110000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011010000011;
SIGNAL_B = 14'b0000111100010001;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001110110;
SIGNAL_B = 14'b0000111011100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001000010;
SIGNAL_B = 14'b0000111010100000;
#5;
CLK_ADC = 1'b0;
#5;
CLK_ADC = 1'b1;
SIGNAL_A = 14'b1110011001011100;
SIGNAL_B = 14'b0000111011000000;
#5;
CLK_ADC = 1'b0;
#5;


$monitor("Simulation_ended");

end


endmodule : TOP_ResonantConverter_control_loop_tb


