-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DOqa28vq/O9Gu6mChwJudQrf+LpZgRwqPzyRfW0C77p+RfN6isagRWY9+XoHJ1zyIfU+cntrrHuw
M43zCQ7e56tsq7GvBlWCbAExdlB0/HsT1nz6iMaalO6BzQciBleTZsRnWRQdiDEzwdo7/j8uybBY
G4J4bjt3uOM4YyD6bUwNOXMkFREY/ylxxLAvFDgpNtN6+wxWNLuoEcQJZ3vtApmvMXH58TkgTtK2
SXsRLu/1W7D/9gPiWQZYHYdPYPG4IP9baKmKwjZBgozMJa3Ls8mHoFWBTn8KGwO+iH7k625VnhOc
ejzdfR2JfNiim5RudZJPUfu2DhPxkiG+wrQtZA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2640)
`protect data_block
Rxw31XyY/a26Tta8DCkfVkWz5j7k7rtF76wVsb2KSKwjOlA7iPs23Y7jR1FRhUn/Ixk6D7z/tbwF
xPbNGkPmIn4PXHmVMp0c1u8SDU2QQH5t7Ow1AxdoexIBgaqrMAskaXINqexYjAIPpUupY60EtF3a
I9tbEVtx3l6D99V44J4OAtZn5mbpsyF5ZE/8BUAsHs4bPgdsIJK+T/JKSzD7Tu1B4wyjWPNdxNPE
iX7qPTK13iW8VGlW13IlyQsuXw3YSeaCY+C3yNMdZQAd6J+wek4v31uvoRX/7mG/DnV+0zY2Be0a
qslk4sfD6jE8p9Vpo4F62XYLcoh6+/bvT8s1kD4I/Ul9TxTXdNa2snT7KHgk/0QP9fPN4Evu+QHi
yfcR+gdvw4Skm3Lo4HabW0XXVTps3oCuZKPyqMR/GzDQnCLv+PxpuylgGOQtmEj5TD95RU8Na+Df
T/ecY1yCa1EN3QyKflwcqSBjQu5SgpMJ+Q95kBiXdL0NrQMnpNOxThk6XnoKTyN9UmuotrqWkWdO
XDPgHLZAbBmCRs18n2ZgFtm44LqqHuq138/5w/53BfRVgOI3R5r7m0Coz+JKAmVA9+AQBvDZPPF6
Nld+Xv/8m8CUBIVNxj3sCLA26fxmjc+xg2LHgkNk3J0jEsvqxlVsnS//DOHDNoV/ajTq/JVoXd8o
rsBA9xXWk9UvNcdLiYm+AvYmHw7JdTho9EW5v/tsfpybgz8Ajx7nMkMSURTrXvpMo7fT3ARH9dRy
17Tq38it5/r2BC/1SMoPQ4pC+FKUKCjQR3+BC74cIUJDREusKsj0VOATjBXottIuR3/ZIT4hdHVF
4ZEhJefL63nqbIbmsaSYLIPUXiuVJuZPuPRMMY+ncaKI2XZkFGzVpsZXAS8UFmRH3FHteo5hDpX0
f1I2VHrOOuAxjV0mUFhJpdXgaBuzNIT/0tc92C9wW0Mrx0we4PJNSmjK85XAiXJw7gR7bXCLhndF
nl4Rkn9rk5jOmSh+ouwLoSU82qKUF1a0t0/9l4oeNDiTsU6MwuQPb4jhIdF7OYTgI+f1IUu9EnmD
lzXvl2K0NAZEZGk5ArHFuNWW9F9lW7fAo5NTr6AsBDuZKvqneE52Qbx8Tn/e8iATRVB1TbPu6jiO
Ar8+CbkaLG6Z/8hB7a1CJ7priewkMhrRSh2i+SHrQQdPMlCcBbvd0fwOxlenCP0oIxMkaoXR7Oyb
RDbBpNG+/uAV6OPcvPn8HN6uwKa6CY47kEv5XTfY7ZUGdZwtFYS1WODnbn+wusUr/MdpXzGnWm1a
3ej8BJHEMDzz0XkWL0/pHAU6h//S/ixxO47X9pYp7tsxyLT3smsWfkT+azFboXseD8x4UnoJf0Xi
QQenT7ZeA+CVdyNcXQGb3jIV1G6XyXwcrFusqiNuitWEVIfmEbih8Nm3yv96x4dJBN6uGGaXYiHA
K6QFf8OLaJwRzbGtRBWCAaG/+HHxWPOg/0HUKwvkJU0Xhv5nbKaqTCltQqZa28J3pHFYfH+01n2M
mxB5kJbo2kJ3pWn4wXmxo5Tjb7FBtbhTUIf64BXf3TiynnyZFaN1XX1USCsGurzcox613E0Kgywq
mQh1Q81Vk2wDmEmE7RMgip8EKQuCHmHUum6E8oTQQLNWHbX5bAxiT6tInPX8HeC0ubK4xvK2g2rp
U+OA09eN202cbjyqQ8FwfViD0kJUG2Jd6/gz9EW6a9mxaARNuaZSk9S8DVxr5fhmY8W0h1/XE7w9
pl6tYf8L+8k88EEUfieMRr+QIzpIKTB2a7tDMBjjKltY7QPHSZugRiLxI59r6PpVPxsjuvBrpfn/
rrB534rgpa2weiLUs679/iZf12+8IBeGwsoZ1db3ENCc67ULJDcUXVj7GSdlFbYS96rrYhDDshMd
rWBiWft0W2lw9urh4iOLEQCibI5AJMFGnjAeEqZifDydv9dVm0JKXYh8jUOOAfJ24GVvwMXxj9lb
Ohjs17gb95mPZCCF3AATgOrcHEF88HbXku7wAfI1JJpPkm/WGaSWFR2n067nMeHc2++dWWrJLYDa
8QSp2ZJU3+96KnddpwoE7LadhZ3Og4K81fyMlQF6OJqgUQzGgxOEreo09kkLpEhLIWZKaKhJWl9T
RqdKjnS1/TM7PMsLO2P1+8aUQzo4Wyuv7do+jpDZFgDLcXEjGtf5q8RUHMtlAEF+DyGj35dhkslI
CLccjtghK/1GdZ4MXkfrqk0ShANOLDwvh43eTltIIQnkdDo6eG7tfpa8QOx0vH4hrcqr6tj/GeFy
NDGvPPqf2cbzvKgtc5MzbPv4iPhPQM5rRZ47u+W22hafNiO7IT90rpSBY64jt/mVhZsBpUING3V/
AxnTPW785mWfpxtazOnAUaTpDjjj0i8dbvfwom7/ryCf2fnYxVeEHyWHV1wvZJ3fJ7H8blghesBl
naqA6F3dhPvgfqd5wF3/i/mKh5t2lu5qKdcnF4sRJvikbY4oQIr+nAQ1pBfyUcPdpFGzQOE1cjl0
1x4cz1ibqZ/VqRNV9ZdUlz8K3Lr0t7u5a3Fxi9U9grgLSGHZyc3C3G35pfJENwBaTru1yXyqk8xU
Hko+5XmNfB1/QUkClm/7kaE0GghCpMPi5WNE8i7K4ikCwPr92fycsRSGbEQI3QaXmtjr6YoqxpyN
twucuzg5/NAXD9hO2Xw+g9nPZMnIdv3o7CwjAK3UkkYcnHgVd3zzyVea1eRPokhBEtBvohmlyzlS
PC/+fdcjRtUwuLnNri7vUnVI5F+gOsnkkUDQhffqXLOueChjxV+1XKzjeH8/sdEkwkNlv7rJ7Laf
3YH7ykAQVUr6/aHIjOkZr1UZvxPzKFU9ASUbBwjP+2cNskaULMzEwJ0ZugjhiMVF9qMPP8JrA613
CIY5XFsPIkVpcFmm5vyDFcSf6hJzetvKhuEo/gy2cab5Qm3gc9c4g2D+IkDYt9r6PrTOx1ppEjJb
/S6mYPOMB8fxJbVlB8bUn9bkabYTratPldb/b+chGhvJLexJLzo82yQOpUgSsdanxveCOOGd/6d/
SH5V/R31193j9s0irxK1u0rZLwZT9z7nVdwjlgOc4alDH43QuSisGcxBrkYfT1hA83QyJSjVUtjR
K9VyegXwth8KJflcDvRaKyJGepOD2CRPSd2L+GCFkN37PhdfJDEy7S8oIWzrrfUF+KtoJ2pB48Nf
t4WfJy6YwMvZ3p8izDS6dmvFENxolIQeX2MdJIkaigkKixRV38CiXQMWa5R2efkZynuvyh4c3SKb
jGDThSSkAVa1JOz3qrOdAOG93fV2Cn0ZgEYiyHJ/EKrYP4c7qjfSEW063LuXu0oD4y6e0BGlikD6
sO2ci6xwWFE6frvv65TpHU/ZlUnixrss6ExWRv5X9MsVZGjvuYqyI2a8zTyRqe+QIElH/tLRoLMD
BA8WRbkwmEDzBvQkgSv8rdGK1szwALGxhiHIzCq+iCo0sCabYRuDp/3XHBSF5M3KEM98h2h7wYkJ
oj+X3sZKgsQ7bOdmtd/N+hnD
`protect end_protected
