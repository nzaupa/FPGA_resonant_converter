// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
0VrQ/RXSOTK/s6k2QtE7phijKVMTAiFufo2jB54qhqsUQyTtkMubaaF5NP4D7lZUt/5/ickB2Fx3
op6mUsTGh+2PPqEPCtLw7m6MiRnway2e1xVoR46OJQXebW5n484fAe3CiJ2zikG+fWGoIFDxyWpH
cxTWVEaouuWgHogJTk4dlPRtUeVMEv+AOo7hCfBqz6X/KBFgo+/E8IWlJV+TD0/k8xhE+rFWfrvG
iDXoYJE2RyDdQO+m6b6qhXFK9yfj7GEX9AD79LYSKKVvXWDBn2+mildyV6zIcp+MrBwvw566Rqm3
zjkY8sv70UaT3hQgD0qbOB9bh04UG35/w5xjLw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 1984)
HnbKykyBOCow39AQLSFNeiiDXvuzvkPrOrUyxnuf0NKWJ9OG8Fq8nyrAGMx5BWcWD2889aEZ5nDI
xyJz39sKD5xXWuircbvY+H684J4itELBpq9QaIWAMs8bhCPMpg5PDB7UswjTBaqgHBzJJ/skS1rw
2c2eKOSOVcvZ53UgTQwNHd1JdQ1dKq0T7PC2ijcoZlP6qIYy55safEInmhxkfOgsrTsgpTx/EU66
gL8wwXgEGXhBrK7XUSytJ+qspS6H9e1PRB4ECMieDzdL773IcVYD6pVRiqsyWgnIWhwMKYs4bdBg
aKU5vlsshZ7OJlhgUq8rsU3IJEN0+rOqbenxEH5uFmMKMo4zPlhoHvpc7IWWIRyNIqYn6pUexkdd
hyoCpli2vO0/Xpl7CCSpJE4ncQUs8n6WA9QMgYsI5HlJtqckKCsCBty8g4s5GFQh324fai32vBNU
uJBj5nQ6ZjpeOdkA/qHcQOEpXmAT22LuUgAY7/nMpUEkoZNyK6pv5puKt02pAHO8G1Pq4vVBjebv
+6/kVghMhgHrjOb9O4dp7J030xDY7lWXIPfo3AEN1VU3AIgsT4gzFDKKQSTh8jdW43xCFMyYzpmF
DYQR8riPD6xP1vHnDQg84moIbvHCAxqSh8XP4F6WNbN6Bkur7ChQUFsXHz99h/KVIBYYcCOjUmcf
mBkNZ+oT6tP2hfGVx+hpAhKl8vYv4PLRGyo/GN3MNc9xu0Uea114KKgYRPAMDowTOeYqyqg7L8DR
jfT2X2zlr16OEb/boClXxGa9wLdT/gZwVc4UPMq5sodcqFlnyXgBOXzzzyGy7Gcf+S1Z86wdUWLJ
pmp64pdU/YNWSRByBtsWKtoJa5O7wOjX6mPCZqPL9wBRoo6MhDM6c/OgssL0Gq9qXhKKMPtvCmdJ
ycl9tL7BPhhCqzPWtxRO/BtL1W5TreeOlLsWggpRw8+OAIXzNH5ovL5G37SMovHNPka0b8MwtdZN
JVhcuobvcupy0kiAPNOWFguZlInq03RCbpw+pAawHT44hTUW/t9bSEHUEcQYBSjvGDf8LYUWJccH
Z1l79erjIhA5oj9dFcKgeazeCYvExMSldRUAlHF+C1BSPRusxbVDN14dPdhA40ysug3MJTi1oi4O
7+EzJUFsO/N3p4CyRn63xKyxH+FjNs84F+PLnZbJrAQmVVvK8hhH6jJGF0BKKBCBBMiy5c0FgrEe
TOyLxTB2Sz6bs6s8jQaE4zeZhmR98gjnvkVB7iYQ5OHYAqBF1RzeEj1lQpgWvLxPw3TweRNVrySm
17XGotw8pDCT6nbPVS++3+rcWYUEJfaDyWwI/UZHYLS6h99F6+dPZAcEsVKHUt30iKglMnt0OUqq
BGogx8zSvKOKzRMqw2kRANo8vNU+GFn2ozCR682TO+8vaLwSCBf/mMS+csDu1mo8ZOl7sY9adZXK
ODjgynwjDDy/90Mhniu7HABS8ljpo/it6evp7Dj7HweY9jNAVZ1MpQWF98NaA6Yqq4xGu5wtB+RI
aM+0VvKjfk60CjWfIUD2fqzsGc/aGsTiBmH2C0sukD9qRnJX3NTE6ZHCV8awbt/xbe8DOrlDnIhr
4YupBKcT6H4e7lF4dbqM8DbipKc8j7wEK2Ok2sM1VGEKH5d0PcH6ZPSZZkqOey7Oxx7hL5aofM5+
SlNvopcJXUfRN9Dq81+fXfl6GWBgZ2aKn0uPvQmvxUkIFdcMLFg/XcHrpUeWIanZd5FTtOZRXMET
+tTsFv9kEwcvUyzOw8Ue/qrbC0/rcxIWzJsfj2UNpUl6QCRbIKBmNwfiG4l7PTy039CWQuhpxkGy
wvzmkN3EE4JZKP8/CFMMuyV0QJ3LeQcwSJGJdQdD5KtRoQThWZgXPJxVF2qR+wDdYnalfAyzpDPH
CeyCcW9hp93HBh6iL4b9M1stKXfU7ZlEUHmUHuoNCFSHxit6F2qqMaymETmOFu/lJI8rFGXHX8O6
hDvwL3aQTQaEAJ5zqnv0ys/eYmIg2ZNPUqWpiR27QL2x8pEELEfKLQIxqfU6msbT7eucXEfreAAB
DsdnGcmRGii/MGeiFm4q8VhJX6sOn+yLviXxpS1SyVmxR2uhg0bFnGrbWCtbkXuhFozn4C47sQLF
NV4ZMqv3myb1MY5VasqEEbhTdA/NFLS6c1LcYzuHLQSMZZMli1oyA+y8scq9SvShDz81TZCKVKTS
hFmUtpZuyhdUnN7oe6rL74sDEEgPR1Zm7/CFeMOJhsH6DWqVhoEieIuRy2eASO4FQkKoMSzrDApQ
cGeT2ouN+37GGXMv8b8v6VcvrdjkFy+3sCCwVgAF7J/SY5jF/LHz3D8mNRe4E9wpWP2VqUvqt4sU
aZBObx2KWYOGjv1w2NHaanhnqPRuJGyQndUnDMwx+IIfH1WR4EDjRtQ6PoaQYolOn5ZlIP2xunjn
blaZHs8dgXPYHMQP+DrhbtYaAtWxQ35/8I8Ynqm7qveg75ZcmmYwrAckBK7mivQYw81HcweqHKqm
xETU0BOP49mGOpISMRzHt7B5BZET8xqCXYM8JEJaM19cCwYxfG+dF90osxeZ2Slph+dKYKyDgEld
bDKv8U8n4Ihmq/BusrBoPwJ1jx22XCAEdbNc2E5P0m2nfpEpNyoUsefhD5UaTw==
`pragma protect end_protected
