-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Gd1/KiIR7DzxRR6v+QYWQtEGKLpxvoHlrq5fVcb+SY9UjkKML+OR5zMIiyNDQHAQv2+HrIGw/Vwa
iIHcPpvgo1mIZifUEgIjI60FCOVS3Y3FOGkPQedE1ypK8WP9NNurb4Ul3s85lrcpcsoHAHhYkGrl
QiS7t9JSAeq/UQZfqkz78DrZaiksffgK+k+59Tibyz+BrJmc2EExL38olluWI93ggB2SajxaOhBe
u0lLlsf8p03hBsLKCmTo/SddffD+6lh3OPQGSdRed9I3uZBvaX69cl5nQ3f1cG41LOqGX/aiZJpP
nwPDwThqHmllV7jjxsLybYyHqyBIXJH9gHgRNw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5264)
`protect data_block
CeIQbaOQHQ2fH9V9nSUCCYg/b0JgmcTD4dCQq0GprHwBI8caPZX3fdWU1CEUxTIrjczpvfPz/yBl
wMn3o0jOSivcSUj40lylr9bLvSlGCJ0DY8q0ydOaWRFvcXHMnO3biN75bQDJWkZt5E2o1M2KWCnP
ekeBtGtMWCOZNEWHHo+P4hvUpqZsUh/vz+v/4h3sCmBefL77Jx5fjqB1iElfe39uHwqoA9cS8LOG
dICZGGdFvc0/25Lpmgp8JzfejFiQheTqRSoerN7YxiwORygNNUxEE/rCZu4Q3Ab905QL18mcMSkM
UHn9Ri/jSAfSPIo4xi8bYLP/KBdtchYNnHzTWg1o0G7qVeMCqlkf6BvXnVDzYnR7XIvFaE9+c7zh
CHYQPHJh/GFdeBuclxgkjQI+vE1EuL5jcZoNXYMFjNIALFBADwHSxnnSUUZOxraty9aZsPclKjoV
TDnIXCknzUC0veJW3OKl85cPe9BlPAiIAbcWYmP6AXEhMIw2cRogYk5He/Z35xVNAfR0xMSTvLL6
ynm5CTfMmEOa7av7aSCljraiG4mpj3l4R21G20djbjQ/0H6DK5rbO1H4AWwCyo7Ww/eEXFKKmjgn
X0UTc4ZRgwXHKkvmhQncDsp6getSxQfxvhs6LAbk4OfEiZL6IOCcik2Xt4vkyBomZBnaqg+lE8EI
uOffHAhnceb47YBgpshZwvsYwADLkY97nERMUwiIU1vSPtDw52OR5LWhsmgBtaQkWgEtJcOfcEeu
TdvT8i5VK+gEbnH6aD46omom9opfWvNBAou759qfojKWNuy8A8hdyzrJB9U38U215ApbYSU9TUd+
xdHAGqY2+l4nsp9olhEuWyVniNLXpCSNDdlfbLSNJ+NCYIK7zu7Uimti3oSkfl4HD3V1R2oEQSVa
gla3EFV/4jtqd0+NuG3QUw/XYYpy4wj3YlNTsnLJt789HN/LOXOKZZuwtTGfGCJg7KIBI8e5K/dL
M/FZfqbbghhV4atUtlgw3pRGdTa97KQOBj2DVdtk6G3MeIWI0Owo0ioaudy2jEKdisFqmQacwKGO
U0QhLSEwaDL9mD7chUkN9u19Bb6cTVrCXJMnpg5uek2LMtcla9kD7/Sa1gToV8w+RNHiQJABf6Ob
jLy2bigjiJg/ckJm6CVqvS24mIjTZkmqugVkRDdExltnX7DJgRctcGqzuS0TFRjvIK4X5CVYDWyY
s8KgsNs0zP8s2132SNBCdE/4hmSDQqDFhz2d7P0zcBdRWgZxvcV9llstqcQFgGAokGanKyWX9CE/
noqu7aAGw/05jSVGWsXgzgpTyx8ZQvbL/qT/uVsqSYjvhLkv/BcB4FU1Da2rA0N219E/zdkHKBmb
xPeQPESgWUDnWn7XoDsC1g78GS8F6EpqaUX+I+pF3guoBIgYoIfaoxhdwA2y2qlhChGl7ZSFGuhb
mhb/c3XjM8BY8u8VHDr6+vYzXzDyNgeJNOqYeWFdQoXhbubUuaMBZe6oJAObJBLiMOawzTHaKcL1
DXqFh21rTPEfeV1OCQjgz0Hqv77BTU7B1fIr/TiJIY7Nw6tB3GNExtJSd6pGk365bBZH2q0UKzyD
R9AvMnl1ICdFBEXSwogJNNCDlyKu6sau09GLPpiV/hy5wWQFVhWb3rqaOW1bVAuWKMeZTuurdLCE
EE8O1UcTOAG5ZZykM/aH7v/Ve7zz3YmToa/pvgz2hQoyJMp2pqyo/vruNE11Qcx8MF5be//U8/Ae
tv2Yxau3mUaMiaj0tQ4QPT2iwNglkmnHo7ZSU3m4p5hAWF4PdfjnGwgtV4bvppA04GlBJkI7PPu8
j8Vf2lIwRzsn6/EaUY0C3LjhS9asX/bodf4wsmns2y7O11iu15VWdu4eQDEZmh2SCAXKzZJD552a
4kex0bDPdiEBWL6FcWZj4qvk3OlZ2R7PBmfi38Du1/vReNbJ11xmCrDcOFSDvTD+GYRvY1Eswz6T
/pFeCsvottjcbToqpJrQ/HZdPK3MjlBWvZQ+fy+Lrfp20uAgj3XeZXrQB054T9hnJRF9ECbPFX4G
4Lz7IBa6zRgVYuugFCyZazh8LLhbRILwM+zTYrLLKDv9XStqZlAps4BQ7fZ+MXeQW5J/2EEnf/FI
Sv84YtHEPfb2mks5QmA3UgiPJRlQAanXfFfPYxxjG6MxPdzvAOAXwFgdv18/e9Z1vQ3X6DUUYIr4
FM4C9OnQFrb29A1uhYnrPP9kIRUEkS3w9GhsJQrts3PESIfIRv+eR83cseqvUixqEIyaCyELlv2r
lZ5l7M4GY+GsAEWqGEHP6Dkf2v8v5AobElhKddTd/R6h/wNfRTTv3Dk8SM+XVvEw+epu3XwSN5Tt
cj3QqtNVe9Mq0PGz8bbnYn0uo5ShquNi9tT3r2LKQdfp61fEFU7DYYZApvCNKs2JshS7uulQx++c
7ZvFGi+9ssqRrZXm3gTwAR4TMPe7gx1YoBSM8+nqqDgJ2cdn9GMPoLfoNlb6G74luGCfO3OhJnZK
eYWatnBhK3lTtmlanID35CUGCbN9CLWukihLJCoIskhc28Ax6nJ6CXOIugb/u/ulgQ/l2xiFHGAW
igeBVzqwZCUD8u9bTbVMiq15oQ8JILii0MC5j4rM6b7suMcL6BcrbFj/O7DZlVi3oX39bd9RcnQJ
odr+PVzJDRpa2s81M77WhrMXqYzBhxr8/6wsCdQlyZV7gdH2LSRqyZzREW0cBFwsGuJ0N5aNdVH6
kj3dj3V74ko5nEAc3tjSE2fNBw8GrZK652pvtfM9pHiZ6UUVUDj4McWn1ssdnEmix+G3NNrUOQ3G
lIIXyy2vMVIB0oF7j+j0wujT9M0pTbHO5vfRaNeCjrR0ZPNZkONf/KeTw+SwkJ/rDd/gmLbxjrlh
f32P5+0hVN5+QfiI8w6L4czdM1IyjC35HZMJbCJ/V12AzM54a6SnlSq2HU4P6D8YQiZqjcljhiAK
jyjcim9IM3FvNnKOMiyoan56ioY/n42dXD12OjI+iMhVkPZAUqLnseGhi3Gtafu8n7Wa10GMUn+C
2miY5FehIuXixETGiR9yQjj0dPZrGtCXlwDIJ4wg/lJ+Mj2JwMQmIqq6HsQuheGn2w2d3TZWcp+e
ZavdS/Xw3aPDqsxU7k6+wxVp1sCYPB0L8s47favKhSRoGCp3HRuAgvL1vy70LqKu1IBoLDvudED8
LghtmX+pUvPCAVlB6f2k/XRxJR2cTaFnC7f+8BIzZipbFwXdv9kZ2J4FDcxqSRfEUSd5KS5ddNO4
d612SDKZcf62+2cZCL2LRc5ypqqFas9OLO8RFe5Ke18jwNqFNN2lYX6xTjmBe8ySjl6zC+B7IHKC
yTVJKdSQWrCWKazXXV9liXncP2PgHumK/2xiujJVRNQQn25BOhskjDYAgtDWvxWq2IjHsS8qqGnC
ZZ7WLrB4j0pW2ZipKlyYbmpky2TIm1x/wM6Ok5uD/LG/4Xglf9jAsWkbkp8LOe3GrtxpJWWLPxbe
qv/pwNrZ5gJT/o/5YEX/kz7TqVTmnAzswWTT0KLFY2vBWc2Du+SvMb6d9+lkZWkmjanHgSVq38Sc
rJGHRcztcJA6RBeZh9QI2jJEsw9QUkwDHlU7pHj1XQ5gId3bJK3EvpmsluuhCy53v+q38VJtm1Az
UuEhRvxqROx94Lcdw6BNvG2pokQ64RN0SVlmwSjrmmiPn6qO+1TdQDBJe+CNI9QpiStuF88irbJp
sZhO6nA5AazLwi8RnqNBkLAgE68nk516WL+mz12WCjDA+Ij5sQmu+HOti3qD2So7GZlCboSwwqvw
yxb42mkU73y6j8WNGJ1q8Anqz9m2dZqXL4ZkIrrwquqjuaHz7WrAzZLCX1iNJya5hDXAlNVsxmOH
LSFgak0qjeaNdTKlUnG+5359mi3nA8DXpcEoFEgeIey5Hvoz6XDk9u1WG4lkVccuv9rdpEmKfX0v
ytqqA/IRKIxCfCd+HlAiAEs8SycvHqadbm0vQ1TviPkj9u2kplfI7zxCa9EaYEmWt/3kkOGuhJHq
qiTR+S691KANkvrFFUCAkAS8LUInZHyuFYFR8LARrfV8Ey2/bN2LkgQppjEBOOSf6MTd3Fi29S9u
IN2lKoh8cT+447jCtAO0Sg9qjvKx9e8recmBPdJOE9fQJOk4l3A983xavTRU7h5GK63sTgmS6fBi
dtNFGtwhrjlwGl9lPCmbasXAMWhR9uwQ+Cj8Fz0vzYYepMRkcK9+NCxwljR9tzIkHy7F2ot29jy4
PTUl/wvkTO40I5Hej5h0LkJYz6a055WZBWqYIZIxv3eq8ciokND2C9mpvNJUJy+y/LwfM7uj9ekK
i/IVjJENMgi9f8URcHJzT/csQYIMTI4TPZC7SZAp0CKCV5c8fUb1RZ9xqmgP8ovgtLujElpSgua1
XtpH1MWumtozQXT3sReyC93a3xWQrLRonS0lESGDBRi5AdGEK3AP6gYyitpCEALCEBjw++S/n3fc
3hbonNShX5QHjFnrEGFQU8lcSYu17sE4mwDpKt3T7g26j5WeotTiwP31z+9TIwX+fVlTmd9DTFnI
6AWajZxCsiwxyIosdaRNHfY5dZFttsvF7lsjOZ2pkW2Gf6UmJWHpzBox/d9qZzHRXM8qfp1tM8Ma
gGsKaH+ygYy1uBPHZizN4MJ9yKZ81wNNYuQa+IYS37VFf4zQOQ5nIyfQ8tSNLHoqtEDI5Li5K5nA
Fm2SkBjKSAP7nV5e6+z2MyUINWKpXw0FKjK85Fh5TRyJOlCdXOWrw7f+X8HEcBOCTAT8tmPaOfwx
Pz9QmxDDJdwdrh6mp+e9JXyZ60Mye/IAjgC6xaToXxQbFHa7JwegVvEaP/Of4HX5d9gFqzpuEgBK
AlamvR5qPX8Bc5gB0gYZPq6XPu65/M9IFf3IoimNuUyA08QcRdTeMPnGLkN6MUFRFFnZe4QmUWLn
W/XLy9arrM4g1Gfzry0p2kDMxg86inx1PWSXpP8d9da/WrJp4Cd67ZbUSXgYbBaK2Fe+Wm9puTBU
AVM+ItTEov0WsQj8pS+ZhS4drJ1RXkvl46IOX2UykttctJyoosEBxdjndGfBZupFlbxHpikeSn85
o0/HvENDipkAqin/GMAtcHnh3uyVL4ApRKlslHz7LvbQDtE4ZMoLpL/fQNfWLV4Qh3DT8o5i/e8U
Th2xXju0e9X1NCikTp99W9Vd8G8MlWhIIhiPHbK1U0MgCRkFC4eUpbL4w+A94wxzXfjMst1K5WdJ
2bZwyZjPVMGS2FmeSrftqKwK8fgDgK9+W/ZBL2lLpfxqs+GvstkgYGFN0RklegVW0SVX1zhmT7nb
frTJWg5Y/jZUAKTNG2IcAHe2B8fngtPIUsugsoQ10t2xW/o+uZk0FpOnfp617yeg1qce8T2S7jFl
PZuq0LLlGlOUq9Zpj8Ff0Bu4KF9zC+93Mj7yfzPZJC5PgNdboYND7I9VRwYQ4OygdI2mgTzgLzAI
Fl/e5+Ds7KRQAjj6e85RLEMae4kEbI1bYKrCgSv8pRY0QHS2q9txuBXK9xlSxltdAmouOBfZn6OT
r4IdOKTVOCPauqdBzFqGvEtMikjwQIIX4AQ+8Vp/LZEm3UgH3qcZ7KmZ7QrO/VOHQUkhEeEVbV5b
C24ANizrJmJk2OngDVze0L6gR8IptRT2NsGDG0sQ0qvxva+sglOX+dja8fJ46Q/93/ylWtnB6iya
eu7pbwdd8gnWt08ltsBLvq8aklcEc/EdGKA3C4nF9uN2z2AomLCqBiFtm1S6Veb/erGubV0ktFnO
hKmkhrJFjzwdq1bPSoeajsTyr8S+cLaJiodWXwN28tEcdgm0qTYUiC1uFiXwhbJ03uUj4U8iCAHI
h3H0ctEvpfIzsojIfg5VDDEExl3nSVOz4GSttTgJ4rVApTtHhoarbkZ6GHK1Lh/hlxx8oJpQU6j+
LTRDb9sz+xrMgfeO4yfyOdK/41xxD9zb701x1Q3iqINTPccigcqDhistHs9iXxJCSX5EF8ytRcvd
F4ygspV4EGpiEphyNE9lzDecs+GWXkafrJb0GUeFSK2gqrrN8zCgpFMi/qkKKPswamTVuAErYJUk
uC+zUVqyzZwJq+XHP7bRHVT8ZhiALC97GiJFKfZRFLn2NAY8ellOW+qUB0Ge8GQQgkAknN1lJQpz
solb2m9zb7T1U5IOAhIlrw71Lpt1TBk8dgd7hOxv38me/m9KR8/NTJAJ2fRqGMai6CQ0GE7VqPMN
H7Ek+kqVWp+LNJlZZspvO/V5NwjXX2Mx5VTAu7tk/oJ2BM8kRxOkftQvt0hfzzbZNsFSHeXFWEkP
3PFPGlVGzn2vLz53747RgXCEe5jQDidb7LFF7epWrNAFa2ljdUeljJnrZo5aE/0SKmlmegi5VLp2
8FPIgQYMxJzDlflcSGrLI6PPFK6T0zRuO++dinHYOPxj1gml54poWN6MfMGOnRokj7bLmv9at8qO
nEgiRfBK9JrIp1QBYoiP0m3vlb/r4MHfy+R8EhZNV4TpCwTkw20vbNIjxSyavnLsDWd6PrDicT0j
oZ0CA2exPzN5f864DVsPjbkYUbO/DFSdyFR1MxFyk4s6ZQQBVUR1uM5fWpN0y/REAJ2v9R6rP3Vo
LKLH/s/Vrcwmq7G9p+Ab/eSEpxm5/DjknH1REGmx5zVCjSEo46H3kXhapxQnCsKaf+Bx3fESz+6Q
DIVCkQ0Rwg3mezIlypLCVBXrq3Pxk0k0rhTNPW5hor1pOLeWKaawoPpcEvyM9r+hqAe/S+vSi/jL
6nhQzWwtTgmJ0GOVuJD+Xf+ocG6R33wzgcc+ZNuliLl1YG2IExEdEGyX6vAIXsCUcY3xMzSogXXP
hy8qPkZKjvNoaeIU4qpyf9IAVri/FtNQQ9gO1LOtUQVQOm1oVHI3EK3GxIHugkOmf8vc74LihN+V
1vGQWnNyYVBcLEB3S7Z5CC+0Z0xuIYE1R9pepxGOdyEOd+XzgX43p98NwCvls+LkIMsBl1o/SM7C
jGA9wDFEgkSR/45HwbJoRJBKL1s=
`protect end_protected
